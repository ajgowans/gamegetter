D��������������������������������Ė����                _]}]_]U�      � � \ W �e�h�� �0�0�0�0�0�0k0�pVpVpVpFppFpppp<�7���p����]���_�T]]]]uu��������7@��UVE  @DUUf����:??:jf��UU�DD    P � ��V��������tu��_W����W3�303�4�L�L3��>D�  PDDUUofԙK�t���������t�[f�UkUDD P U���������5O3S��� 7�>�>f:�� ������9r9qNqN\N�S�      4 � � &)��<�<�����<�<f�%�%I��{���[}��k��=PCU��=�C���  ����ff��d&��c�S�S�S�S�C�p��   � |�W | � <���h�� �0�0�<�<�>�>i-�}T�T�U�F�W���~�����U�����UU�� �*���f�� ���U�����������������w�� � � p � �f��UU�DD Z �Z�����_��W��Z��jڑڨ6�6f6�6f6�6U6U6U�T�Qj�� � w�v�� \ L � < U������������UU��  ���� �� ff�� �� UUUU  �� � ��u��0u0�pW��&)��̿|��������fl%�%oIo�[���_���_U���������U��� �j��� �����&������ �U�U� ����_ \ � \ p p p p�h��#�>�>�7�5�;�>k>�V}VyV~F~Fuvv6�6���jU�j�ڪ6�M��jcj��dژ�TZT6D66D� j� �                 P � �rVq��U������*��cɓ�N�PUUDD�O\5��U}w�u7��75u5�� U�����V��������������q�r�©ɩ&����D��D� ����^k��wM]��7�=�&3)֪X�\�ܿܪ|�|�|f|%n%�I��[��������j�VU��U����j��6(6�6�6�6f6�6f66666��j�|w_]]��WwW����h��'�7�9�9�;�>�:i:�vT�T�U�F�W��o~��z��M�7��V]�v����_��
���ff��`���Wէڧکj��l^s�py�y\ww��}W{Z �Z��j�媤�Sw�]�Z�(l��|��f��f,T,D\D\_�]�y��|�p�ܗ��L�L� U���>��?��w�_uU��|U��uu_]�W����oW\]\_\]|=�0�0�0��� 3 3  &)�������f%%I� � 5       �?0U�]u�=��W�]qWq�_��w]���u�q�w��5        ��_�� � � � � p � p��  U��UT���������j�j����o��f��?T@�Uo�� ��9m6�9g��f���� PU���
��U�� �        5 7 � ������������U��W �         � � �         ���P�PUP������  ���������������Z���]\[�[[VlV�Z�[�k��U�V�j����u�ϫ�^�s�ӬS�T�t��0005���0 3 �jjj���������ڪj�ڪڪڪڪv�]�]�]�jjj�j�jǪ��j�j��ݪ]�v�v�v��Z��g-�m�k�lű����V\V�[ݯ~�7]?�9~y_�חwW7��=���|7���        {�{�{=�u�u�}�u��ww�W�^�~�ޱ^�]l\l�����w�u����������ww��������1����]�u�u�w�׷^}zu���u�}�w���u3ww0�       �����q\qq�q��1�qp�q���3����������]q{qrq�}�s����5�5��q�s�q�q�]���_�w�uw�]����u�u�u����]�W\�\w�]1W3�1p1�3 <    ����������������� � = 5 � � � �  9 9 � }�� ]� < 7 � � � � � 7 5    1 1 1 � � � 1 1    3�OO�L��6�N�N�SӔ��3�3�3�O�LnLnOnMn7n5n7:�8�83�<�4��s�s�]��;��^�]�]ow{�{uv}�u��]7u7�����u\�p�p� �         S���ĩũq���������������������������u�u�u�q�q�q�ũĩĩħĞĞs��M,M,=-<��S�T�뤧��>�:�M�O�M�3����\�0�0��uWu�SuSu��L�L�LWpW�u������ 7  ���������ꩤ�����S�T�>�C�T9U:UN�O�L��^�W�^u�}u�uusuq}\w\��wwW� � 0       ���������������j��g?� ? 8 � � ���� �<��U��_��5_7�7 � < ��p��lf���g �W�W�W��U�? ��  �����������V��g�W�~�_��U� ������j�� ? 9 6 9 ? �� U��UU��UUUUUUUUUUUUUUUU��WUWUW�WWW�WU�UU5W5\5\5W5U5WUW�W�W�W�WW�UUUUU5W5|5���\UWUWUW�WWW�UU5U5W5\5\5\5WWWW�WUWU\U��\5\5\5W5U5U5U��WWWWWWW�\5\5\5\5\5\5\5WWW�WUWUWU\U��\5\5_5U5U5U5U��WWWW5W�WUWU�\5\5\5\5\5_5]5W]W}W�WWWW�U5U5U5W5\5\5\5���WUWUWUWUW�WW�UUUU5W5\5\5WWW�WUWUWUWU��\5\5W5U5UUU� ����?                   ? ��������            �_� � � � � � � � � � � � � � � � � � � � ����            ������_U�_�__U���W�_}__}_}��_}_}�_�W�W�W�W�W���W�W�W�W�W�W_}_}_}��_}_}_}�U�U�U�U�U�U�U�U_}}}�}�___}�_�__U_U_U_U�_�_�_�_}_}_}_}��__}���}�}�}�}�_�_}��__U_U_UUUUUUUUUUU�W�WUU                U�U�������U�U�UU��������������UUUUU�_�z�_UUUUUUUu��u�]���^w^w{��]�u��U�UUWUWU]U]UuU�U�U�U�U�UuU�U�U�U�U�UuU}UsU�UU}U�ժ��UUUUUUU�UUU}��u�u_�uu�U��Z�U�V[l�o�l?��[UdU�uUUUUUWU}U�����[���ֿտտ�o���j�j�������������z���������^��U�UUUUUUWU]U]U]UWUWUU�W�^UyUyU�U���_�UU�ZUcU]U]UWUW������|�_�_�_�_�_�������}UW�w��ꪪ������  ��  ��������UUUUUUUUUUUUUUUUWUWU^UyU�U�U��y}^W�Uu�u�_�{y�y������U�U�U�U�Uޕו�����w�y{yz^�W�Up�_�p���������UUUUUUUUUU�U�W�W�U^UWUUUUUUUUUUUUUD�D�1DOD�W�}��_7p�s6s�_DDMDuD�UGDwWD\�DD��_qUUUU}U]���W�U�U�U?���1sqs~LzzLt]���?1�?����1�����۪l�m}�U�U�UG�qDMDMDD�DG�DOD�W�|��_7p�s6s�_DDMDuD�UODwWD\�D��WtUqWUUUu�_}�W�U�U���U3�s�1sq^zLzzL��O�?1�?��?�����תW�\�qutUqU��G�uDMDODD���=DGD�W�|�]UWUwUvU�WDDMDuD�UODwWD\�D��WtUq_UUUu�_}�W�U�U���U7�w�5su^zMzzM��O�?1�?��?�����תW�\�qutUqU��^^G�uDMDOD��LDGDGDGDGDGDGD����DDDDDDDDDDDDDD����DDDDDDDDDDDDDD����DDDDDDDDDDDDDD��DDMDMD]D�M�4MMDGDDD�O|=�O�OODD�O|=O|=�ODD=O|=O|=�ODD=|�=�?O|DD�O=O|?�ODDDD�?�DDDD=|D=|D=�DD��D��D��DDD�?OD�OODDD�?OD?�D�DDD|�D��D|DDODGDODDD��G��G��GDD�O|�G��DD�O|�D|=�ODD�xO-OO�?DODD�?OD�D|=�ODD�OD�O|=�ODD�?O|�G��DDD�O|�O|=�ODD�O|�?D|=�ODD_�G�����D�DD����������DOD����������D������������GD�W������������WUWU�������������������������������\TG�����oN]N����TUEF�U��iN���Uq�����}��O������������������gf��gf��gf��gf��gf��gf��gf��gf��gf��gf����������ff��ff��ff��ff��ff��ff��ff��ff��ff��ff���������f>��fޙ�fޙ�fޙ�fޙ�fޙ�fޙ�fޙ�fޙ�fޙ��ߪ��?��gf��gf����������ff��ff���������f>��fޙ��ߪ��?�g>��g��g��g��g��g��g��g��g��g��������W=W�W�W��߬��?��ff��ff��f���fޙ�fޙ�fޙ�fޙ�fޙ�ff��ff����������ff��ff��f���fޙ�ff��ff��gf��gf      ��      ? ���V��f۪��?   ��UU  ff����   ��וۀ˖۪��� �����[��?�:l4�4l4�4l4�4l4�4l4�4l4�4l4�4l4�?��[����W�W�W�W������  ��  ��  ��  ��� +�WU� \�W����   ��UU  ������   ?��U� 6�5���� ?<<��[�kլ6l4�4l4�4l4�4l4�4l4�4l4�4l4�4l6k�[���<<�\0g�gŧ՗�\5�  ��  ��  ��  ���?[�k�����k�[��?l4�l4�l4�l4�l4�l4�l4�l4�  ��ww33ww����    ��ww33ww����  DDDDDDDD��ff��ff��g���gޛ�gޛ�gޛ�gޛ�gޛ�gf��gf��g���gޛ�gf��gf����������gf��gf��g���g���ff��ff��ff��gf��ff��ff��f���f��f>��f��f��g��f��f��f��g���=��|=�׻ݼ=�UUUUUUUUUUUUUUUU����?                   ? ��������            �_� � � � � � � � � � � � � � � � � � � � ����            ������_U�_�__U���W�_}__}_}��_}_}�_�W�W�W�W�W���W�W�W�W�W�W_}_}_}��_}_}_}�U�U�U�U�U�U�U�U_}}}�}�___}�_�__U_U_U_U�_�_�_�_}_}_}_}��_�?� ��? <�?��?�?    �?�?_}���}�}�}�}�_�_}��__U_U_UUUUUUUUUUU�W�WUU<<<�?�?<<<��������      �?�?      ��?<<<<�?���?<�?���?�?�? �� �?�?�?�?������<??�?�?�<�<�<�<                U�U�������U�U�UU��������������UUUUU�_�z�_UUUUUUU]U�U[Wm}����U[U[U[UmUmUmUmU[U[U[U[�V�V�V�V�V�V�VU[U�U�U�U�UUUUU�UUU�UUUUU�U�UUUUU�U�U�U;�6�6�5�յUmU[U[U[U�U�VWk]}��u�]�]�W�W�W]WUWU]U]U�������^U������������  �  ���V����UUUUUU�u]���w�w�wW�W�~��� 7 7����yUYU�U�U�W�~���W��]��usu[uU�UW�W�W�W�U��������������������Zl�𯯪������UUUUUUUUUUWU}U�U�UUUUUUUWU\U\UsUsU�_UuU�u�U�UuUuU]�W}UWUU�U_W_]�uUuW�]�}u�_�_�_�W�]�]�Yj[jW�^�_5p�_ \�W�U�WZ]�UUUUUUUUUUUUUUUUUU�?�?    �?�?<<<�?�?<<<����������?<<<<�?��?�? �� �?�?�?�?������<??�?�?�<�<�<�<                <?<�<�<�?�??<��?<�?�   ��<<<�?�?<<??������          � �   UUUUUUUUUUUU��������UUUUUUUUUUUU   � p \ W ����5�55u5u5u5u�u����U�U�U�Uu�u�]U]U]U]UuUuU�UU_U�U�   �  � 3 3 ��_|UWUUU�V^ p p   ������  ��k�UWUU]UuUUUUUUUUUUU�U]UWWU? �   � �U=U�UU���    � ��0�p��  �/p�kU�U�uU]UUUUUUU�~UUUUUUUU�    5 � � W\\�\�\]\]\]Z]W]WWUWUWUWUWV][]UuUuUuUuU]U]UW�U_U_UU_��u�uu����}U�U@��_@]����U}U�p��Wq�����U W W \\ \����*�)�͞q�J�"�9�9�;����٦٦���©ª������ܭƮ��:�:���ų��#�-�-���=���= � �		*0	>D	R �
!+1
?E!S �"&,26:@FJNT �#'-37;AGKOU^ � $(.48<BHLPV� �%9��	��hqyW �)=��	��irz� �/C��	��js{ �5I��	��kt|� �M������_clu}� �Q������`dmv~� ��������XZ\aenw �������Y[]bfox ��� �gp+ �* �� �)	
) �)) �)� �)� �)� �)� �� �29 �3:@ �-4;AF �.5<BG �/6=C �07>D �*+, �18?E+�, � !"# $!# $%&'#(( ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	ZH�KZEHI�LZFIJ�MZGJZ
H�KZEH
I�LZFI
J�MZGJZH�KZE
HI�LZFI�LZFI�LZF
IJ�MZG
JZH��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	ZH�KZEH�KZEHI�LZFI�LZFI�UJ�MZGJ�MZGJ�YVZ�FXO�PZNO�PZNO�PZNO�YVZ�FWO�PZNO�qPZNO�J
Z�rZH�KZsOPZNOI�LZrZJ�MZtOZO�PZN
OZH��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	ZO�PZNOPZNOZO�PZNO�PZNOZH�KZEH�KZEHI�LZFI�LZFIJ�MZGJ�MZGJZO�PZNO�PZNOZO�PZNOZ�EKZEKZEKZQZEKZEKZEH�GMZGMZGMZSZGMZGMZGJH��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	ZH�wO�PZNO�vHI�LZ�FI�LZuO�qO�KZFI�LZRZ�RZ�rZFI�LZRZTZQZSZNPZrZFI�LZRZ�RZ�rZFI�LZtO�MZNO�MZFI�LZ�FIJ�WO�PZNO�PZNOJZH�KZEwO�vHKZEHI�LZFLZ�FILZFIJ�MZGMZEH�KZGJMZGJZ�GJ�MZH��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	ZO�PZQZQZuO�qO�vZ�RZRZRZ�RZ�FKZNxZNO�yZRZSZNMZNOJLZ�SZ�RZRZ�WOPZNOPZRZtOZ�R
ZO�PZNW
OZO�PZuO�qO�v	Z�RZ�RZ�FHwO�PZQZNOMZQZSZNxZFILZ�rZ�RZ�RZFJMZNO�WO�MZNO�WOJZH��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z
\�]Z[\Z�^a^a^a^Z^a^a^a^a^a^�_Z_Z_Z_Z_Z_Z_Z_Z_Z_�`Z`Z`Z`Z`Z`Z`Z`Z`Z`Z\�]Z[\Z\�]Z[\�]Z\�]Z^[
\�]Z^\�]Z_Z�^Z�_\�]Z`[\�]Z`Z[\�]`ZH��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z\�]Z^�Z[\�^Z`Z�^_ZaZ[	\�]ZaZ_`Z�`\�]Z^Z^Z^Z^Z[\Z�_Z_Z_Z_Z�aZaZaZ_Z`Z`Z_ZaZaZ[]Z�`Z�`Z�^[\�]Z[\�]^�_Z�^Z^Z_Z�[\]^Z_Z_[\�]Z_Z�_Z_Z_Z_�`[\�]`Z`Z`Z[\�]`ZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z\�]Z^[	\^Z�_Z^_�Z[\�]`Z^[\�]Z_`Z�_Z_\�]^Z^_Z[\�]_Z�_Z_Z_�\]Z[\�]`Z`�ZaZaZaZ_Z_\�]Z[\�]ZaZ_Z�^Z_\�]Z�_ZaZaZ[]Z_Z�_Z`\�]`Z[\ZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z\�]Z[
\�^Z�_aZ[\�]Z[\�`
Z�^Z\�]Z�_[\�]Z[\Z�_Z�[\]Z[\�]_Z�[\Z�^Z�_Z�aZaZ_Z[\�]Z�`\Z�_Z�[\]Z`ZaZaZaZaZaZaZ[\Z�a\�]Z[\ZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z\�]^Z[\]Z[\�]^[\�^Z�_Z�a`Z�^_Z^Z`[\�]Z[\]Z�^Z_�Z_Z�^Z�`Z_�Z_[\�]Z_Z^[\�]_�Z_Z�_Z_Z�^Z_�Z`Z[\�]^Z_Z`aZ`ZaZ`_Z�_Z_Z�_Z[\]^Z�_Z`[\�_Z�_Za_
Z�_[\]Z_Z�_Z^ZaZaZaZ[]_Z�`Z�_Z_Z�`Z[\�]`Z`[\ZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�zZzZz�ZzZz�ZzZ�zZ�zZz�Zz�Zz�Zz�ZzZz�ZzZz�Zz�Zz�ZzZ�z
Z�zZz�ZzZ
zZ�z
Z�zZzZz�Zz�ZzZ�zZ�zZz�Z
z�ZzZ�zZ�zZz�ZzZzZzZzZzZz�ZzZzZz�ZzZzZzZ�zZ�zZ�zJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Zz�Zz�ZzZ�z	Z�zZz�Z	zZ�zZzZ�zZzZzZz�ZzZzZzZzZ�zZ�zZzZz�Zz�ZzZzZzZzZ�zZzZz�ZzZ�zZz�ZzZzZz�ZzZ�zZz	Zz�Zz�ZzZz�ZzZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Zz�ZzZz�ZzZ�zZzZ�zZ�zZz�ZzZzZzZzZz�ZzZ�zZ�zZzZ�zZz�Z
z�Zz�ZzZ�zZ�zZz�Zz�ZzZz�Zz�ZzZ�zZ�zZzZz�Zz�ZzZz�Zz�ZzZzZ�zZ�zZz�Zz�Zz
Z�zZ
z�ZzZzZzZzZzZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Zz�Z	zZ�zZ�zZ�zZzZ�zZzZzZzZzZz�ZzZ�zZ�zZ�zZz�ZzZ	zZ�zZz�Zz�Z	zZ�zZ�zZzZ�zZz�ZzZzZ�zZzZ�zZz�ZzZz�Zz�ZzZ�zZzZz�ZzZzZz�ZzZ�zZzZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Zz�Zz�ZzZ�zZ�zZz�Zz�Zz�ZzZz�ZzZz�ZzZ�zZzZzZ�zZ�zZz�ZzZzZz�Zz�ZzZ�zZ�zZz�Zz�ZzZzZz�ZzZ�zZzZz�Zz�Zz�Zz�ZzZzZ�zZ�zZ�zZz�Zz�Zz�Zz�ZzZzZ�zZ�zZ�zZz�ZzZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�cd�eZfZfcd�ef
Z�gZgZg�cdeZfcd�ehZgZfZigZ�gZ�gZgZg�ceZigZcd�ehZgceghZ�h	Z�gZ�gcd�eZcd�eZfhZigZ�fZgZ�gcd�eZfZhZhiZig
Z�gZ�gfZfZ�fZfiZhcd�eg�ZhZiZhZhZ�fZ�ghiZiZiZiZ�fZifZhZfZg	Z�hZ�hZ�hZhJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�cd�eZcd�efZ�fgZfc
d�eZfZg�ZgZ�gZg�ZhZc
d�ehZgZg�cd�eZcd�eZgZ�iZ�ighcd�eZceZcd�egZ�fZ�gceZiZhZc	d�eg	Z�fZ�gcd�eZfZhZfZ�fZfZgZ�hZ�hcehihihJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�cd�eZcd�eZcd�eZ�fZ�iZf�Zfcd�eZgZcd�eZcefg�ZgZ�gZ�iZgh�Zhcd�eZhifZcdeZgZ�iZ�gZ�fZig�fcd�eZhfiZgZ�hg
Z�gZ�gZfZg�ZiZfcd�eZihZ�hZgZg�fZ�gZ�fZ�fZ�gZgh�cehZfceZgZcehZ�hZgZ�hZ�hZ�fZ�gceZcd�eZcehZihZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�fcd�eZceZ�fZcd�egZ�iZ�hZ�fhZcd�eZcdeZ�cegZ�fZ�iZ�iZ�gf�ceZgZcd�eZ�fd�eZgZ�hZ�iZ�gZ�gh�ZceZifZceZ�hiZcdegZ�gZ�iZ�fZ�gfcd�eZihZfZcdeZhZcegZ�fZ�hZ�iZ�ghiZfZhZcd�eZcdeZcegZ�hZ�iZ�iZ�iZ�gcd�eZ�iZ�ceZcd�ehZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�cd�eZfZcefZfZfZ�fZ�gZ�gZhigcd�eZfihZcegceZgZ�gZ�gZ�hZ�hZ�gceZcehZfceZ�iZiZiZigZ�gZ�iZ�iZ�gfZceZcegZiZiZ�cd�hgfZ�hZ�iZh�ZfZfZi�ZiZiZfcdefZ�hZgiZ�iZ�hZ�gcd�eZhZfZi�ZiZ�iZgZ�giZ�iZiZi�Zgcd�eZhZiZ�iZ�iZ�g	Z�iZi�ZiZhJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�konkZkn�kZko�ko�kZ�mZ�mZmZ�mZ�mk�ZknkZkmZmkZkZkokZmZ�mZ�mZmZ�kZ�mk�ZmZkZkmZmkZ�kZko�kZ�kZ�mZmZ�kZ�mkZ�kZkmZmkZkZmZkZmZ�mZmZ�mZmZ�mk�ZkZkZkmZmkZmZkZkokZ�mZ�mZmZ�mZ�mknokZkZk�Zk�ZmZk�ZmlZ�mZ�mZ�mkZk�Zkok�Zko�kZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�ko�kZkokZkZk�ZkZkZ�mZ�mZkZkZkZko�kZkokZkokZ�kZ�mZmZkZkZkZk�ZkZ�kokZmZmkZkZkmZ�mZ�kZ�mZmZ�mko�kZkZ�kZkmZkokZkZmZ�kZk�ZmZ�mZmk�Zko�kZ�mZkZkokZ�mZ�kZmZmZ�mko�kZkZko�kZkZmkZkmZ�mZ�kZ�mko�kZko�kZk�ZkZ�k	ZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�kZkZkZkZkZkZkZkZkZkZ�ko�kZkokZkZko�kZ�kZ�kZ�kZkZkZkZkZkZkZkZkZk�mZ�k
Z�mkZkZkokZko�kZkZko�kmZ�mZk	Z�kZ�mkZkZ�kZko�kZ�kZ�kmZ�kZ�kmZ�kZ�kZmkZkZkZ�kZkZ�kokZkZmZ�kZ�kZ�kZ�mkZkZkZk�ZkZkZkZkZkZkZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Zk�Zko�kZkokZkZkZkZkmZ�mZ�mZ�mkmkmkm�kZmZkZko�kZkZkZkZkmZ�mZmZ�ko�kZko�kZ�koko�kokZko�kZkokZ�mZ�kZ�kokZk�ZkZk�ZkokZkZkZk�ZkZkZkZkZkZkZkZkZkmkZ	k�mkZkZkZkZkZkZkZkZkZkZJ��p%&'()*p�!# p�+,-./0&3p� "$p&�@?>=<;:pB�CDABZ�}	Z�ko�kZkZkZkZkZkZko�kZ�mkZ�kZ�kZ�mZ�mkZkZkZ�kZkZ�kZkZkmZ�kZ�kZ�kZ�kZ�km�kZkZ�kZ�kZ�kZ�kZm�kZ�kZkZ�kZkZ�kZmZ�kmZkZkZkZmkZ�kZm�kZ�kZ�kZ�kZmkZkZk�ZkZkZkZ�mZ�kZ�kZ�kZ�kZ�kmkokZkZ�kZkZ�ko�kZkmZ�kZ�kZ�mZ�mkZkZkZkZkZkZkZkZkZkZJ� �� �� �� �� �� �� �� �� �
� �� �.5 �(/6 �#)07 �$*18 �%+29 �&,3: �'-4; � !" � 	 
 �d��� �  �! �"#$%�		
	�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`>�>�>�>�>�>�>�>�>�>�>�>�>�.�>�>�>�>�>�~�>�>�>�>�>�>�>�>�>�>�>�UUUUUUUUUUUUUUUU��WUWUWUWUWUWUW�W�W���W*�
gJ�Jg
�)W���W�W�WfW�W�W�W�W�WUWUWUWUWUWUWUWUWUWUWUWUWUWUWUWUWIWWeW�WUWUWUSUSUCUU+T/T�P�B�
+��           ��c�W���@   � W*W�WUWUWU����UUUUUUUU�U�T
TPUTUTUUUUUUUUUUUTUPURUBUJUJUBURURUBU
U*T� ����UUUUUUUUD@ *�*��U�U�U�UUUUUUUUUUUUUUUU@U
T�P� � �        �
�*���������*�
�
�
�
�
������U� � @     �
X�VUZUe����UUUUUUUUUUUUUUUUUUUUUIU	U)U)U�U�U�������UZUUUUUUUUUUUU�U�U�U�U�U�UmUmU�U�T�T�P�ԪVjUUUUUUUUEUU����.����< *���������������� * * *�(�"�"�"�����������jU  ��ZUUUUUUUUU��UUUUUUUU�_���ZUkU�U�U�U�UUUUTUPURUBUJU
P�B�j�jU�U�U[U[�V�V�V�V�V�[�[[n[YVUVUV��U]U����������U�U]j���տU�UUUUUUUUTUPUTUPUTU@U
T��� ��
 
 
 
   ��*�*������������������UU      �U�UUUUUU����UUUUUUUUU�U�UmUmU[U[U��6�6�6���[^mzm굻���횭��^�w�������u�Wj�U5U5U5U�U�U�U�U�U֕W�W�_�{������}�p5z����u����@_S]�z-�?�UUUUUUUUUUUIUJU
�*������ >       @ P  U           � � ��*�*U @      * ��UUUU����UUU��k�VZ�U��U�UuUuUU��� � � �����0�3��5��wV�[�m�m�m�m�}���p��� � � \ \ � � p ����߿�k5VVV�U�UUVUYUfU�Yjf�����3p3�0���������U�UU�UUTUTU ��0                              � ������� � � ��
U�UUUU����UUU�_U�U]Ws_s}]}�u�W}\]p�p=pp�s3�����zU�U�_�������]_]W]�]?_�]�]�]W�U����5�\�ܷ��l}l�[�V�� u]��UV�       ���������wkݩg���VUUUUUVU[Uk�����      � 0 �:�5�U�V�j � �              BU    � UU�����UUUUUUUUWU]Uu�u�w����v�v�v�]�]�]�]�]�]UWUWU]U]W]WWWW�U�_��3�0 00090�0��[��;�:V�U�U�U�UUU�W?� �����������������������ff��PUBU
U)U)@�
�:��         0 � � U�              TT UU          ����UUUW�UuUUUUUUU�_UUUUUUuU�UUWUUUUUUUUUUUUUUUUU��5�_�UpU\�\�W�WUWUW�Ww\w\wpw�U_0�� ��5�5���?�0�0000?������������������wf��fUUUUUUUUUUUUT��Z�o?�     � p p � � p �        � \�5W5|� U T   UTUPU    ��UUUUJU* ��U�UUUUUUUUUUUUUUUUUU�W |��UU5U��U�UU_UUU�_wU�WwU��U5U�� |�_WuWu��WuWu�_WuWu�_����U�}�U�����w( ��Z�VUUU�U�:��>   1 3�3\1�     5 � \p��W \ p � � � l l �  �T�  U��jhUVU��UTR�T�T�T�T�R�
U�U�UUUUUUUUUUUUUUUW�\�p�sh�h�U�U�U�U�U�UsUpU\UWUUUUUUUUT�
�*��`�R�R�JUI_IIU�U�W�WXUZUVU�V��   �p=\����5  5 5        0 ���\U��[U�q�q��quq���p���:  * ��U�UU����� ���UU:U9U9U9U9U:����� � � � ���U:U9 8�0�2�ʥ�U�U)U%U�U�U�U�U�U�UUUUUUU�U5 5*0�2�ʙ
e*�)U*�)U*��U�U�U�U�U�U9�:�� >                     � p l � l � � �3 � �<Q�_���U�W�]UUUWU]U�Z�o � ê�U}U�U�����                                             �                        @@T @ PU           ���p�p��Ӭ���\������<�>������U�U�u�UUUUZU��� � \ p � |��5�_���5����UVU[UZU_�����  ���
�
�� ��*                      U                 > �_��_W��Z��UU���s���� � � �p�_UU�W�^ZuVu�_U��>ϖpU_U_UU�U���?�7�u�  �����             � 0 � s�\0W�U0� 3                       @  T             �            � fÞz��ÿ��U3U�U�U3�0�|��U�U�U]U_��� �   M
@  ��ZpUpUpU_U_U����     �  �����  ?<������UUUUUUUUUU��33      U@         0000�    ����  ��C�<���0 _?��3;   ���j�UUUU��������[��U�j ��@  T	 �*U�UUUUUU����    �   0�� �<��<�0<�
����UUUUUUU�U5��3      � 0    ? � �    �<��C?<��Pp���������V�UoUZUUUUUU�W�\�\�WU�U�?�  PP� ` X�VYU�UUV���� � � � � � � � � � ��������5���3��� � � � � � � � � � � � � � � � ��<���=���P�O�u�_�z���ϕ�U�UΕÕÕ�����9��� �T�� ���U�U�U�U�U�U���UUUUUUUUUUUUUUUU����������������������:�ꫪ��+��+��������������������������������������������*��k��������j�������������������꫺���n�k�[�>�ꫪ�������VWVWVWVWUWV���������������������������������꫺����������������������������������䪓�N�:��:�ꔪ��@��:������������������������������������V��j���������꿺��ź����[Vko��������ꪺ���������������������i�V�֪�������������������ª*�*�����������������������������������������������ꪩ����P�S��>��T�@��:��������������j��j��������������꿺Ʈ�k�����\U �� �����ƪª������������ƪƪƪƪƪƪƪƪ�Zƥƪƪƪƪƪƪƪƪƪ��ƺ��ƪƪƪ�����������ꪺ����������������������������ꪩ��P�C�����Ϫ������ꪹj�j�Z�Z�V�V�V������U��������������\�:���ê����j���f�Y�V�j�U���j�j�j�Yjf���櫺����������ꪪ�������������������������������������������������ꪪ��j�VUUUUUUUUUUUUA <��O ; ����WU? ���:�꿪��ݪݚk[�Us�V       � 00�0̌̌00P0`0��U0P�C�� ��� �W����������������������������������������������������������������������������ꪫ�������n����T�W�W�^�y�u��U����UU  �� � @ ����V�UU@� 00000��0��TUeeiijZViYf�j���jUU�?�����ѹ���������}���������������������������*��������������������������������������ꪪ��~�ꪪ��������� ������j��ꦾ�����ׯת�Z�U����U���� ���W@��@�f���T�P�@e � T P @     ��0032322@1%�%i�F�0�P��� ��W�������������������������ê�>�ꫪ�����������������W��_�����_?�    ��j�j����g����u�u�0�0��������������3�<���UT� ������������������e���d���P���PVP�P���\���P���e���f���������������������������������*������������������������������������:����<��#�":�鿧��V�U�UnUnkkj V�U�U�W�W�����^U� ����� �TT:P�P�C��������������������j�j�j���jU�j���������������������������������:�:����������:�:��������ꪪ����3��ë���j�Z�֫�ڶ����U[UmU� �������������������UU  ��������������媵��������������������������Zj���>���:��ΪΪ���?�:?�CCW�\���ЪC�>�������*�������������������������������뾾��뺮�j�֫����������k0�üά�l�;�ꫪ�����������������C�C^C:O�y�:������:�:�:�:�:�:�:��N�N�N�N�N�N�M^N���P���:�:�:�:�:�?C�T�������������꫻��U� �������������������*����������������������������*��������������jj������������S������������������꫺��*���������������������� � ��>�Z=���ꪯ���꺪������������������������������������������������������j������j��j�j���������������������s�s�CUNUU;P���������������_���㵯������.������������`:X:�V���Uc�cUc��U��V�����������������������������������������������������������������j������j����Z���}�������������U�W:]:u:t*��  �U�����������m;Tꐪ����N��î?��MzCzSzS�SUSUUjU������e���f�������������������f������������ꪪ������������������������������������������jj������������T� �?�ꐪC�N��:U:U:V�Z�Z�V�U:V:�:��������:�������@�?�萩C�N�N�N��;�;�:�:��N�N�N���������N�N�N��:�:�:������������������������������������^�z�ꪪ��������:����>�:��z�z�������z�z�z�_�U�����j����j�������ꫪ��殚�����j�j�j�j�j�誸������ڮګڪڪv�ݿ��몾��k����������j�j�����������j�j�j�j�j�j�j�j�j�j������䚤�����������������������������������U�U�WUWU^U^U�W\p?p�p�\�WUuU������|�WUUUUUU�U�ի����������j��������j���������ꪪ�����������������������꫺��꯫�����������ꪪ����[������j�j�j�j�j�j�j�j�������������������������������������������������������������������������������֩�f�����������j�Z�Z�Z�Z�Z�V�i�j�j�����������������������������UUUUUUUUUUUUUUUU��           CA  WU       ��<3�3��3<��_��� C�    ' � WWW	W�WeWUWUWUWUWUWUWUWUWUW�W�W�W�W�W5WWC�P7T7T����]�}�7�7\7p���p�\WWWW�U�U�uw�wUwUwU�uWWuW]W]Wu[�gf��gf����������                        @ U              �s��U�U�U�UpU_UUUuUUpU������?� <       (��`UZUUUUUU�U�ի�ꝺ]^W�W��u�uյյ����PUS��U]?�<�<� W�U�u��UW�]�W��j���j�}k��]�uk�k�mݭ]�u�v��U���5T?UUMUNYCYSZSZ�� ��3��0�0�70�\�W��    �      M@5 5@��T� � � � � � <        � h�ViUUUUUUU�����[꫾�W�U�U���������k��V髥��wu~�^�^�S�S��������Z��Z���Wv_�|�|��W�U�UUWUWUU�]W]�W}�ת~�֫j���֭ڭj������ ��s�p�p�p�\�ת��U�U��� � ?�      P @     UU @                   ) � ��UbUbUYUUWU^U^UWU^Uz�z�_�\�\�uu��~�WuU�_�U3�554���S�L�MC<���N�N�N�C� 55���3�3��W�WU_U��UUUUWUUUUU��   @NU   0���� 0       T T      UU D               ��bfYUUUUUUU�՗5T��Us��WsU]��0��� _�]���U�U�����_�_���M�O����溵鯤*��>�:�QG�E�Q�����u�w�~�uj]�W]U�U�UuU�U�U�����           @ P       UU                               @@     �`�`eXUVUVUUUUUUUUUUUUU_U�U�W�^�^_^�~�w�w����<�7z5_5W=�7z?{�^]zu{u^u^�W�\��?�?�������z�z�^������������}�w�w�{�v�y�v�y�������          TP          U @  @                   @ @� p    \ p p�) �U	U�UUUUUUU�UW�U�U�]�UUWUWU]�=�@�P��Z�V�U]U]U]U�UT_C�?��?\]u3��uu]�6�6�ڥj�����������������z�z�z�z�z�z�z�^�^�������              P @ P@     UU                     @ =�<_��� ��}uU_U\U\UWUWU_����W�U�ZUkUUWUUUU�US���x�x�y�׾שWU�U�U�U����k�Z�UZUTUUUUUU����_|UT�P�@� |×}������������֪֪֪֪V�Z�Z�Z�Z�Z�Z�Z�j�j�j��       P              �<0S���� ��}u�_UUUUUUUUU]W_�W�UUUUUUUUUUW_�_�_}_��w�}�յU�����V�U�U�U�U�U�U������UW����������������������������ڪZ�Z�Z�Z�j�j�j�j�j������������         @  T              @@    : 9 � � � ����W���� @@PP��55C�@��TCUC�P�P���4���S�C}>U�T�T������������������ꪪ��������Z�Z�j�j��������������������������     T@   UU                 D@      �  � ?��\�W�\�]�]�]�W�W9W9V:Z:�:�:�:��~����ߟ��:����V�U�իu�]��U�UsU]�_^]�]�W�W�UWUyU]z瞻����Z�j�j�j֪֪Z�Z�Z�Z�j�j�j�j�j���                   � \ � w w � \�D�pp�� ���<�ܮ_�z��`�XUTUUUUoպոToTUTU�[�n4n�[CUOUU: ��� �{�ꪥ���U�U�U��n�k�[��������������k�[�^�^�z�z�z���ꥪ����������V�V���         �0�ܬ\�\�G
G��������{U���<� ����S�T����U_U�W��� �����U�W�~��U�U�U��[�n5n�[UU�W5}=���_�w�}@���|�������]UqUqU�U�U���������~VzUyU�U�U�U�U�U�U�UyUyW�WyW�^n^��n��ë����    7 � \ \ p p � \ � ; ;�Έ���������{�]UU�j����� � � ��p���{��U~�^������ZzUzU^UWU�ժ��^�W�U��z�zUyuy���6��yZ9U=U7T�@U���W�UUuU�U�U]W}Wu]�]�u�w]�u�u]�}�uU�U�U]U�U�U�U�U��eթթ٩�������i�e�g������0 ���p�\W�u��5u5��U��?     @��C�� � ������ � :     M77@5           �(i�UUUUUUU�U�W�W�\�\ps��Ϊ������\�W�U��W�U5�4p0\�WU_UuU�UUUUUUU�U_Օ}�חU}ի�w�]��W}]]u�VU]U_ծ���WV����������j�Z�ګ֭�����                 P@   @U                          TP P@    @D        ��`	`	XeY�VUUUUUUUUWU^U^UzUzUzUzUzU{U]�{�꽥k�V�UUUUUWU]�u}�W�UZ����[��A�z\��]]t����N�N�O��:y:y�T�T�T�S�S�����     T   P                  @@       ( ��UiUUUUUUUUUUUUU�UUMU�U�UCUMUUUM�C5 @ P�u5u�]�WuU]UWUUUU����W�Uzx�_��uW_�]]WU��W�U�U��W~qWqUq�q�q�qqqq\q\q\�ťT���� � � � � � � � � � � � � � � � � � � � � � � � � �@���� � ���Z�U�U�U�U�U�U�U�U�U�W���]���w�]�����w�u���U���U�U�U�U�U�U�U�U�U�_��թץא޿��ޥו���w�U��ު����מ�^������^�n�n�n�ŷ����UUUUUUUUUUUUUUUU������j������������������������������������������j�j�����������������������������i�i�i�i�i�ij�j�j����������Z����Z������i�ij�j������������U{U~U��ꕪU�UUUUUUUUUUUUUUUUZU�U�����W�����������������������������j�j�j�j�j������������������������������j�j�jjjjjjj������������������������Z��������������������������f�j�j�Z�e�j�����������������������j��^�W�W�������Z�VUUUUUUUUUUUUUUUUUUUUZU�������U������������������������j�j������������jjjjjjj�����������������������j�j������������������������������i����������������������������j�jZe�Zj�������������z�z�^�^�޵�կ�j�VjUVUUUUUUUUUUUU�U�U�U�U�UUUUU�����U�WWUW]��ꪪ�������������������������������������������j�������������������j�j�jf�f�f�f�f�f�f�f�f�f�f�f�f�f�f�f�������������y�^�^�^�ު����z�zmzkz[�Z�V�V�V�U�UkUVU�W�W�U�U�UyUyUyUyUyU�U�啧����������꪿��]�]�u�����������������������j�j�j����������������������������j�j�j�j������������������z�^�W�W�W�ת��z�^^^U[U[UkUkU�U�Z������[�VUVUVUUUUUUUUUUUUU�U�U[U[U[UVUVUVUVUVUVUVUVUUUUUUUUUUUUUV�V5j-�.�����������j�j�j��������j�j�j�j�j�j�j����j������������������yZ^�޿��k�VmU[U[UVUUU_����Z�V�Z�[�Z�V�V�Z�[�Z�Z�Z����U�UUUUUUUUU�U��ZU�U�U�UUUUUUUUUUUUUUUUU�U����ەVUUUUUU_�p���
����������������j����������������j�j����j�j���������������U�U�_�UUUUUU�U�������VmU�U�U��k�nU�U�U��k��U�U�������U�UuUuU�U]Z][]k�׻W�W�WUU�UuU�UUUUUUUUUUU�U�U�~�W~U�UUU��ݿ������������������������������������������j�j�j������������^mWmW�պ����j�U�UUUU�_�p�� � � � ������UU�_=�333333=��VU���     U@U��AU@ �U� T   �U�WU@] u����U�U��y�zU^@� WU�T�U� U �Ͽ������������������������j�j�j����ꚺ�n�[�[�V�ZZjUUUUUUUUUUVUZU[UVUZUUiU�U���� p p p�����UW� 3 � � 5         � � �P��W ? ��PU   �T� T    � U�@U     �U� U    � U�@U  ? ��P�ë�Z�V�UjUj��-��������������������꫾Z�UVUUUU��� 9 5�5��pU3U�UUUUUUUUUUUUUUU�U�U�V�ZU[U[UkU�U�Zǫ�              UPW���T���_�� � ���_�� � ����� � � o�m_k[ [�Z�V�V�U�UkUZUVUU�����U�UU�߰���������f�f�f���������龕�UmU]_ukulլճ5�5��oU�Z���UzUz�z��ե_�zUUW�� � �ÕÕ�U�������������������pUpU�Z�[�[�[�[������Z���������������������ժժUkUkU�U�U�U�U�U�U�U�U�U�ժ��������������������WU�U���������������j�j�j����������Z�V�U�U�U����� �<�?�7���U�U�_��ZV�[�o�o}YUU�W5�7;�:��V�����������������j�j�j�jۛ۝۶[�[�k��ھ��ֻ���������������f�f�f��������������j�j�������������������U�U�]�]�ת������WWUUUUU_U���������������������������j�j�j�j�j����j�j��������j�j�j������ߪժժu�]�U�W�׬?�:����������i�i�i�i�����������������������Zi�����j�j�j����Z�����������������z�z���_�UU�W�W�^����W�U��U������0:�� ����������i�i�i����������������������������������矚�V�k�����ڪ���������������������j�j�j�j�j�������������������������������������������z�꽪��������W�_���UWWW�WUWUU�U�U�U[U��U�=�=��p��_�W��UU��  ��    ��  �����������j�j��������������������������^����K�
��j&� %�V꛾f�몾������������������������������j�j�j�������������UU��������=j�h�ڪ��]�u�u�w_��wUUUUUUU_U�խ�����կ?��7p�_UU���U}�_ �� 0 0� �������������������j�j�jj�i�i��毐� 夺�����������������������������j�j�j�j�j������������j�j�jj��U������𪯪��������:�:�:�z�:�N�^�^����W��_z�޵޵ߵ��u�_�^�����������������������������������������������f�i�i�i�j�j����������������������������������j��������������������������������j�jjjjjj�i����Z�������������Z��������������������������������������j��������������j�j��������������������j�j�j��������������������������������j�j�j�j�j�������������������������������������������j�j�j�j������U��������������������������������������������������j�j�������������������L�L�L�L�L�L�L�L�L�L�L�L�L�f�L�L�L�L�L�x�L�L�L�L�L���L�L�L�L�L�( ��.;HUb������� � "/<IVco{������� �#0=JWdp|������� �$1>KXeq}������� � �%2?LYfr~������ � &3@MZgs������� �'4AN[ht������� �(5BO\iu�������� �)6CP]jv�������� �	*7DQ^kw�������� �	+8ER_lx�������� �
 ,9FS`my�������� �!-:GTanz��������d �( �'2I������ ��=Jax����� �3>KVbmy������ �(?LWcnz����� �)4@MXdo{������� �*5ANYep|������� � +6BOZfq}������� �!,7CP[gr~������� �"-8DQ\hs������� �	#.9ER]it�������� �
$/:FS^ju�������� �%0;GT_kv�������� �&1<HU`lw��������d �( ��?LY����� �'3@MZfA������� �(4AN[q|�����A� �)5BO\gr}������� �*6CP]hs~������� �+7DQ^it������� � ,8ER_ju�������� �!-9FS`kv�������� �	".:GTalw�������� �
#/;HUbmx�������� �$0<IVcny�������� �%1=JWdoz�������� �&2>KXep{��������d �( �(5@KWco{����'�� �)6ALXdp|������� �*7BMYeq}������� �+8CNZfr~������� �,9DO[gs����'�� � -:EP\ht�������' �!.;FQ]iu����'��� �"/ GR^jv�������� �	#0 �S_kw�������� �
$1< �`lx��'����' �%2=HTamy�������� �&3>IUbnz�������� �'4?JV'���������d ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`րx����^�p���������ʋ܋� ��$�6�H�Z�l�~�������ƌ،���� �2�D�V�h�z�������ԍ���
��^����$�f����,�n���Ԑ���
��.�@�R�d�v���������Бb�������j���������Ԗ��"�<�V�p�����6�ȘZ��~���
���@�қd��������>�Пb�r�0�����������������������������������꫾�������������ꪪ�����������ꪪ����������몪����������������������������V�����������j�U�_����������WUU���������j}UUUU}��������WUUUUէ������v�UU�W�������]}�WUU}u�����jWWU]UU�թ������  pUUUW������5 �pUUU]�����v5 ��]UU]�����v ?�WUUu�����] ��WUUuu����] �WUUuu����] �WUUuu���jW5 �{}UU]թ��jW5 ��UU]թ��jW� �W�WUWթ��jWU|UU}�Uթ���UU�WUU�_UU����UU�U_�WkUU����UUzU]�U�UU���vUUUUUUUUUU���]UUUUUUUUUUu��]UUUUUUUUUUu��]UU�UUUU]UUu��]UU��UU�_UUu��vUU�U��W]UU���vUU�  @]UU����UUU  @WUU���j_UU=P�UU�Y�jU�UU�O�_UU_����W_U�U��gg? ���_UUտn� �  ������j�9 ?  p�V�o�k��� 8  ���W�Z׿j��  gg�~�j��jg�  ��իj�je����Z�jկm0�����������������������������������꫾�������������ꪪ�����������ꪪ����������몪����������������������������V�����������j�U�_����������WUU���������j}UUUU}��������WUUUUէ������v�UU�W�������]=�W�|u�����jW \5 �թ������  p  W������5 �p \�����v5 ���? \�����v ?��� p�����] ���� pu����] ��� pu����] ��� pu���jW5 �{�� \թ��jW5 ���? \թ��jW� �W� Wթ��jWU|UU=�Uթ���UU�WUU�_UU����UU�U_�WkUU����UUzU]�U�UU���vUUUUUUUUUU���]UUUUUUUUUUu��]U�UUUUUUWUu��]U�_UUUU�WUu��]U��UU��^Uu��vUU�����jUU���vUUU���ZUUU����UUUUUUUUUU���j_UUUUUUUU�Y�jU�UUUUUUUU_����W_UUUU��gg? ���_UUտn� �  ������j�9 ?  p�V�o�k��� 8  ���W�Z׿j��  gg�~�j��jg�  ��իj�je����Z�jկm0�����������������������������������꫾�������������ꪪ�����������ꪪ����������몪����������������������������V�����������j�U�_����������WUU���������j}UUUU}��������WUUUUէ������v�UU�W�������]}�WUU}u�����jWWU]UU�թ������UUUUUUW������uUUUUUU]�����vuUUu]UU]�����v]UU�WUUu�����]]UU�WUUuu����]]UU�WUUuu����]]UU�WUUuu���jWuUUu]UU]թ��jWuU���VU]թ��jW�U�W�kUWթ��jWUW~UU��Uթ���UU�WUU�~UU����UU�U_�WkUU����UUzU]�U�UU���vUUUUUUUUUU���]UUUUUUUUUUu��]UUUUUUUUUUu��]UU�UUUU]UUu��]UU��UU�_UUu��vUU�U��W]UU���vUU�  @]UU����UUU  @WUU���j_UU=P�UU�Y�jU�UU�O�_UU_����W_U�U��gg? ���_UUտn� �  ������j�9 ?  p�V�o�k��� 8  ���W�Z׿j��  gg�~�j��jg�  ��իj�je����Z�jկm0�����������������������������������꫾�������������ꪪ�����������ꪪ����������몪����������������������������V�����������j�U�_����������WUU���������j}UUUU}��������WUUUUէ������v�UU�W�������]=�W�|u�����jW \5 �թ������  p  W������5 �p \�����v5 ���? \�����v ���� p�����] ���� pu����] ��� pu����] ��� pu���jW5 �{�� \թ��jW5 ���? \թ��jW� �W� Wթ��jWU~UU��Uթ���UU�WUU�_UU����UU�U_�WkUU����UUzU]�U�UU���vUUUUUUUUUU���]UUUUUUUUUUu��]UUUUUUUUUUu��]UU�UUUU]UUu��]UU��UU�_UUu��vUU�U��W]UU���vUU�  @]UU����UUU  @WUU���j_UU=P�UU�Y�jU�UU�O�_UU_����W_U�U��gg? ���_UUտn� �  ������j�9 ?  p�V�o�k��� 8  ���W�Z׿j��  gg�~�j��jg�  ��իj�je����Z�jկm��??�?�<?<�?�����������??��� �?�?��?<��<�?���<�?�? �� ��? <�?���? ��?<�?���?< <  ����?<��<�?���?<�?�? <�?���<<<�?�?<����?<�?���?<  <�?���?<<?���?�? �� �?�?�?�? ��   �?�? �?�?<�?�<<<�?�?<<<���������?�?������ <<<?<��<<?<<< < < < < < �?�?<??�?�<�<�<�<�<<?<�<�<�?�??<��?<<<<�?���?<�?�   ��?<<?�?�?��?<�?�����? ��? <�?��?�?������<<<<<<�?�<<<<<<���<�<�<�<�<�???<0<??���??<0<??��� � � �?�? ?��� �?�?      ��      �/�����������/                ���\UUWUU5WUU5W�W5W\5W\5W\5W\5W\5W\5W�W5WUU5WUU5\UU��� �?  |�  W�  W�  W�  W�  |�  p�  p�  p�  p�  p�  p�  p�  p�  �? ���\UUWUU5WUU5W�W5WW5��U pU \�  W5 �U |U�WUU5WUU5WUU5������\UUWUU5WUU5W�_5� \5 �_5�UU�UU �_5� \5W�_5WUU5WUU5\UU���  � �U \U WU�UUpUUpuU\�U\�U\uUWUU5WUU5WUU5��U �U  � ���WUU5WUU5WUU5W��W  W��WUUWUU5��W5  \5��W5WUU5WUU5WUU������\UUWUUWUUW��W  W��WUUWUU5W�W5W\5W�W5WUU5WUU5\UU������\UU5WUU5WUU5W�_5W\5�\5  W  W  W �U �U p�  p�  p�  �? ���\UUWUU5WUU5W�W5W\5W�W5\UU\UUW�W5W\5W�W5WUU5WUU5\UU������\UUWUU5WUU5W�W5W\5W�W5WUU5\UU5��W5  \5��W5\UU5\UU5\UU����_�_}��_�W___}��_U�_�__U���W�_}__}_}��_}�W�___}_}_�_�W_}�_�W�W�W�W�WU_�_�[�W�UUU�U�UDD�O|=O|=�ODD��G��G��GDD�O|�G��DD�O|�D|=�ODD�xO-OO�?DODD�?OD�D|=�ODD�OD�O|=�ODD�?O|�G��DDD�O|�O|=�ODD�O|�?D|=�OD��DDD�}�1�_MDDO7p�suDD�6s�W�_UGDwUUU?WU}��D\U]�1���sqDD�s�W�~L�_U�zqUU�zLt]������G�?۪�1�l�qD?�m}��UMD�ձU1լUMDD��DDDG|���_MDDO7p�suDD�6s�W�_UODwUUU3WUu�sD\�_�1�}�sqD�W�^�WU�zLtUU�zqW��zL����OתG�?W��1�\�uD?�qu�tUMD?�qU����ODD��DD��|�=]UMDDGWUwUuDD�vU�W�WUODwUUU7WUu�wD\�_�5�}�suD�W�^�WU�zMtUU�zq_��zM����^Oת^G�?W��1�\�uD?�qu�tUMD?�qU����ODODDDDDDDD�D��?������D�ODDD���������������������O������������������?�?�������GDODOD�CD��GDDDDDDDDDDDD����GODD|DD��G�����?��������������D�������O��������������DD�����D�GDDD}D
��<<��?�?<<�<<<<?<<<?<<<<<?<<<<<�<<�?<<�<<�<<�?<�<<�?<�<<?<�<<?<�<<<?�?�?<�>��<�
� �?���? �?��?<  <<<  <<   <<   <<  �?<�?  �?<�   <�   �?�<  �?�<  <��?�?�?<��?�?<>��<��<<�?  ��?�?<��<<�?  �<<<� �<<   ??<<?<� �?<<   < <?<� �?<<   > <�<� ��<<   / <�<� ��<<�?    <�?� ��?<�?  � <�?� ��?<   � <?� �?<   �<<?� �?<     <<<� �<<   ��?�?<� �<�?�?  ���<� �<��?  ���?<<<<<<<<�?���������������?<< /��� >  �?�?��?<< <�� <<<�?����<<<�?�?  ��   ��? < <<�?���?<  ��?<<<�?���?<? ���� � � � ��?<<<��<<<�?���?<<<�?�? < < <�?�        ??   ���    �    _�   �UU  p}}  p��  �<<7  �07  �<<7  \��5  W}}�  WW�� �uu]]��UUW�U��U W�z�  |�_=  �W�   �?    p    _�   �UU                           ??   ���    �    _�   �UU  pUU  p}}  \��5  �<<7  �07  �<<7  W���  W}}� �UW�U�Uu]U��UUW W_��  |�_=  �W�  ��         ??   ���    �    _�   �UU  p}}  p��  �<<7  �07  �<<7  \��5  W}}�  WW�� �Uu]U�UUUU�U�U W���  |�W=  �W�   �?    p    _�   �UU         <?    ��    �    _�   �UU  pUU  pUU  \WU5  �UU5  ��U5 �o_U5 p�UU� \UUUU�UUUU\UUUUpUUU� pUUU5 ��UU  W�   ��        _�   �UU         ??   ���    �    _�   �UU  pUU  pUU  \U�5  \UU7  \U_7  WU�� WUU]�UUUU5�UUU�5�UUUU5 WUUU WUUU \UU_ �U��   _U   ��    _�   �UU  < � ���?�����?��� <            ��  �����? �� �������w?��������3���?0 ���?  ��������?����  ��?�����03��  p��  p�_  ��x�-�x�C-�p�B��@�����������������?�����? �� �������w?��������3���?0 ���? ���������? ��� ���?0����00��  p��  p�_  ��x -�x�@-�p@��@�����������������?�����?�W����w����������������<���������?����?�����������������������������?����00���������?���  <�������?��3� ������?�����?�W����w����������������<���������?����?��������������������������00����?������� ����������0�0���?������3��?������?�����?�?�����?�������_�_�����}��������������??�����?���������� 3� ���3���<<���3���0����� 0��0�<  <��?��+�3��?0������?�����?�?�����?�������_�_�����}��������������??�����?���������� 0 ���3���<<���3���0�������0��0�<�<�<�?<���3��?0������?�����?���/����������������?<��?��?  ��?  ��<���3��0�3 2����:�#�� �,�8�� � ����*�� �� 0��� �� ?�� �������?�����?���/����������������?<��?��?  ��?���<����3 2�3<�0����:�#�
#�,��� � ����*�� ������?� �� ?�� �������?�����?������_?������������?���������<���� 0��Ï
����/���L?0���<�1���<�1��� ��,  ��0����� ���@��������_���S�������?�����?������_?������������?���������<���� 0��Ï
����/  ���  0���?�0��<0�  �� ��,���0���������L��������W���S�������?  ��    �������   � � |�l�����,�<�`�����̣��8�\�����Ȥ��4�X�|���ĥ��0�T�x�������,�P�t�������(�L�p����4�d���ĩ��4�l���ܪl���������$�  ���������  ���������?  UUUUUUUU�  _UUUUUUUU�  _UUUUUUUU�  _UUUUUUUU�  _���W�W��  ����_�_��  �UUW}}W]u�  ��UW]u�_u�  _�WW]u�Wu� �_UWW��Uu� ���WW�WWu� U�UW]uW]u��[UUUUUUUUU��UUUUUUUUUU�p�WUUUUUUUU�\�UUUUUUUU�����������?< ���������  �/   �W�  |UU=  WUU� ��_�Wpuu]]p]�Wu\]��u5\]��u5V]��u�W]��u�Wuu]]���_�W��UUUU�VW�_Օ\���5\�Z�^5p�V�WpU_�U�U�_U WUU�  |UU=  �W�   �/  �?���� ���?���?����?������������?�<?0����������/�����?lU:��?�jlU5�U��������}��}߬V5��   ����9ly9lU5lU5lU9�U-�e�� � ��������pw�U5|w7��=�U5���kV���?  �� �Yp�5pU���\������ � �     �  O�9pDt8�LD���D44��3�    | � ����U�����:�:��*����������?��{��{}�{U��U�_��{U�����꫾���?��?��꫷�������_��������꫾���?��?ת�����U�{]�{]�{��{U��U���������?��?WU�WU�ww�w�ww�ww�ww�w�WU�WU���? � 0 <0��pyl�5��6��6��6�5�k���? x�\UwW5wW5wW�WU������\U�pU���?�� �U�]�]5�]5WU5��W��WU�WU�\U5�����W�u5l}5p]5pU5\U5\U{U��;<�: � � �U�]k]-|]5pU5pU5pU5|U�����??<  �� ��?���ܽ=����6��6�z7��6��ګ������� ��?���|�:���������6��6����pUpUpw=w�ww�U5pU\U\_�p ��� \U\U�U���]WU\�\U\W\_��<��u=w����ի�5�W��U�\U�pU���?\5����pu\w5|w5�u����{U�\U�\U�p�5�W �  � �U\U5�U�W��WU���?�<7��77��7��<0 � �U\U5W���U�WU���?p}\�5��7�<70  <  � �U�Up�\�5WU��U��U7|U=\}5��? <  � �U��U�W��W��\U5pUpUpUp}��   <�<�U7pU��7\U5\�5\�5p}�U7<�<    �7 �� 7p��U���U�Up�� 77 � ��� ��l�ܝܝl���:��:��:��:����             � �l�:۝�۝�k�ꬪ:���� pU�_�]5�]5w]5�W5WU5\U��p� ��  ? ���_w]5�]5�]5�W5WU5|UWU7\��  � �UpUpU\�5\�5\U5\}5p}p}�U �  � W�U5�U5p]�p]�pU�p��p�7p�5�U �    ���p�:|];{W��W�kU�|U5pU5�U �    ���p�:|�:�����k��|�7p�5�U �?���<\�7p�lt�P�pJ\�1�<� 0     00��-�,��<����0                 � �6� �  <             ����������������W���__UWU�����__��_���������_�_�__�WU����W��_�_�_��������WU�_�_���������__�W�WU�����������������   l  [�[��6[m��[m��[m��[m��lo���l�� ��6 � �  � �l5lo�6[m��[m��[m��[m��[���[ͳ�l�6�       �6����l���[m��[m��[m��[m��[m�6[m5l� ��         ��l��6[m��[m��[m��[m��[m��[m��l��6��                 �  \7  79  �8  �  �                          �   _ �Z9 �V9 �>� �C� �W� ��� ��:            �  ��? �V� lU�lU�l����:�9�oil�Ul�������<  <   �  ��? �V� lD�  L�0!#2���8 #)L�U,�������<  <           0   L  1 �  0  � � 0  ���  22            ��       � �    �U   �U5   W�   ;W� �;W��5��UUs\�UU}�U]U}\UWUsp�U�p�_�\ ��\ p�?W �W�U �W�  �_��  ��7  �� �UUU \U�W �� �  ��       � �    �U   �U5   W�   ;W�  �;W� <\�UU�\�UU�5�UUU�5\UWUsp�U�p�_�\ ��\ p�?W �W�U �W�  �W��  ��5  ��_  \U�   �U=    �   ��       � �    �U   �U5 ? W��� W�p5�;W�p��UUs\�UU}�U_U}\UWUsp�U�\�_�\ ��W p�?W �W��  �W��  ��7  ��=  ��_ �}UU p���  �� ?    ??   ���    ��  _=p5 �}�\ p�p_ p�W p�}�  \�s�  W]]5  �V�5  W_}5  |�W  �W�  �_�= ����� p�[�_p�W�_p���_p�W�_�_}_�  \�U  W5W5  ��?   ??   ����   �p  _=p �}�\ p�p_ p�W p�}�  \�s�  W]]5  WVe5 <W�_5 ��W W��� \�_�= �����  �[�_ �W�_ ���_ �W�_ \}_�  \�U  W5W5  ��?  � �W� pUU\UU\}_W}_5W}_5W}_5UU?�_�5\�W\UUpUU�W�  �  � �W� pUU\UU\UUW_}5�u�5WUU5UU?�_�5\�{\�^p�W�W�  �  � �W� pUU\U}\U}WU}5WU}5WuU5W�_5WU�?\UU\UUpUU�W�  � ����ˮ�F���ï
�[��� �`���3��������x��������4���]�������������Ʈ>^�>���� >!>�^�� �^��>>� ��׮ޮ������ >�^^�N~��^^� �N~�~!N^�^~�  �^��#��%�.�5�:�A�.'>�^'^�n#n�~� >n�~'.�^^�.>� �^�^~~�T�Y�`�i�p�y���n�n^>�^� � %>��.>�^.�^%n�n �>N�N'N�n'������������>�^^��� �.%NN� >>�^n�~#~��.�>�NN�n�ѯد߯����� .�n'N�^~�Nn�~�� �..�n�^!~�~#�!N�^��� �N%~���!�*�5�>�G�P�.>�^��>!n�n'~� �.N�~��.�>>�n�N'N�^!~�  �.#^�>�n~���k�r�{�����������.#>�n �N!^�^n���>N�Nn�.�^#n��%�� � '~%.�>�N�n�N^n���ưϰڰ����.�.���>�N!n�~� % �^���.�N�^'n� �^n~���N^�~�~ �N'~!����"�-�6�A�J�U� �>^�n #N�^'~�NN�n�~!~�.�^�n�� �>^�~�~!.#N�n��.�N^�^��N'N�^!~��p�{�������������>�N^�^%��.#^�nn�>N�N%~�� �^~���� ^#n�nN�N~��#.'>#N!^n �N�^��!ұݱ�������(� � N^���.�>�n�n~N~����>�>#N#n�n#..�N�^!^� �.N�n�~>�Nn���%.'>!^�^~ �.^!n���E�P�[�f�q�z�������.�N^�^#�� �^�n~�~.N�N^���N^nn�~'.n�~�~ N�^�n���.#.�N#~��^�n��� � #^%^������Ųвݲ������ �.N�nn���.�NN�~#~�>'N�^�n!~�.^~��� �.^�n��>�>N�n��# � '.�Nn��.^�n!n�~�.�^'~'��/�:�E�P�[�f�o�z�  �^�nn�.N�^!~�~%N'^�~���.�>�>N�N.^�n#���'N�n�~�� �.^�~�� N�>#~�~%��������ǳԳ߳� � .�N�^%n�>>�N^�^#��.�Nn�~~�.#.�N�n!~� �>^^�n�~�>N�^�~��.�N'N�n�~~�N�^n�~������#�0�;�F�S�`�m�.�>N�n~��� '.�^'^�~! �>�N!N�~��..�^n�n!>�>'^�~'��N!N�^'n���� �.>N�N~�>N^�nn�~.�^~��!������������ǴԴߴ�.�>>�n�~ %N�N'^����.�.^n�~~�>�N!n!n���.%.�^#~~�� �N^�nn���.�>^�^#~�>�>�^�n~�! � >�^�~!����'�2�?�L�Y�b�q��� �N^�~�~% ^�n~�~���#N�^#~����.�>>�^^��!.NN�n�~!~�.�>�^�nn�� �>~�~ N�N^�^n�n#.�>#^�~%~����.>�NN�^�nn�������ȵ׵����� �N%^�^!n�>N�^�nn�~�� .�^�~���!..�>�N�^%n�~!.�N�nn�~�NN�^�^%~���.�>>���n~� �N'N�^�^#~'��>�N�^#n!n�~��.�=�J�W�b�q������� � !N�^~����.#>�>N�^�~.�N�Nn�n��.!>#^�n%~�.�Nn�~!~���� >>�N�^~��>�N#N�^�n%n�N�^~�~���.^�n����¶Ѷ������'� #>�^'^�~��� �>N�nn�~�~.�>�N!N�^�~��.>^�n�~��� �N�^'^�~��� ..�N^�n~�>�>N�n�n#~'.�.%^�~'~����.n�~~����F�U�d�s�~��������� �..�>�Nn�~� >N�^#^�~%��.�N^�n�n'���.^�^~�~>�NN�n�~����.�>�^�n�~��� .N^#n!~!�%N�N'^�n�~���>�^n����շ�����'�6�E�T� �.#>�>^�n�� .�N�^'n�n�>�>^�^n���.�^n�~�~#�'.%N�^�n%n� �N^�^���>�>#N�n�n~�~.�.N^�^���! � .�>NN#^%^�n'n���q�����������ɸظ�� � ^�n~�~��..�>�N%N�^'n�>�N%^�n#n�~�� ..�>^�n�~N�N^n�~~���>>�N�^�n#��.�.!nn�~����>�^n~~� #^^�n����.�>�>N�N~�~;�3�;�3�3�;�3�3�B�3�B�B�K�K�K�B�B�K�K�U�K�K�K�K�U�U� � � � � 	�����Թ�T���Ժ�T���Ի�T���Լ�T���Խ�T���Ծ�T��� � �>� �^�>  ^  �> ��� � � � � �  �> ^�^  � �>�  �� � � � � �>� � � N�^~� �� �� � �>^� � �~  �^� �  � �>� �~  � � �N  � �  �.� �> >�n .� � �^� �. .� � � �^ � �n�>� �> �^� � �n  � � �.� �> ^�N �� �n  �n�  �N� � �>  �n�. � � � ��  �^� �>�^ n� � �.�> n� �~ N�.  �^� �n~�N N� � � �^ ��N� .�  �^� �n N� �n� � � � �. .�^� n�~� ��� � ��N� �N� � �^n�n~� � �� ���n  � �^  �.�.^�n  � � � � � �>�.~��  � � �^ �n���~  � �^�^    � � �  � �.  �>�  ^�n  � �~�^N�>� � � �.� �� �~�n  � � �~n�~�   � � �.  � �>  �~��n�L^�>� � �.�   �^�n�~  � � � � ��� �~� �. ^�~  �.  �~� �^^� ��N  �>>�^�~  �.� � .  �^�N� � �^  � � � �N� � ����  �N ^� � � �~ � �.  �>�^ ~�n  �^�n �� � �~~�n n� �.  � � �.�   �^�n~� �>  �^� �~n�� N�>� �.�> � �^ .� � �^N� � �.   � �. N� �n^� � � �N�^>�  �^� ~� �~  � � �N �^� �N>� �N  � � �~�� �^N� �>  �^� �nn�^�N>� � �.^  �n�N  �~��  �.  � �^  �.� �^  �n�n�� � �. >�^�>n�~� �� ^�^  N�N�� �n�^  � .� �. �~ ^�>>�n N� � �   �^� �� � ��~�n �^ n�~�> >�.  � �^N� � � �n n�~�> �^� �>�.  � � �^�n ���n� �^ N�>�~ �^�>�. �~�� n�   �  �>� n�^�. N� � �^n�^�>  �. �.�.N ��. �>� �^�.�  N.�N� � �.�>>�  .� �> .�  ^� �n ~�~  �^� �  N>�.  �^�~n�n��..�n  �. �^ > N� �^�N  �.�>��n ~ n� �> . �^�n ��~ n�^ �N�^�N  �N� �>�^ �^ .� ��n�� �   �.�  n�~ ��� �n ~�>� �..� � �^ ~�^�� � . .�^�N �^�N  � � �   �N�^  ���� ~� �n ^�NN� �>�.  >�N�  .�.�>  �.N�.  � �^�n �~�>N� � �. >�� � .�   �N�^^�>�n ~�n�^  � �> .� �N�^~�^ ���^�n ^�~ .N� �n�~N >�. � �.^�>� � �N� � � � �.>�N  �^   �.�  >�n�~�N��  �.�>^ ��~  � ��n�^  �~�n  ��������������������������������������������`��
�������l �m��� -� =���! ]�� ���h�`� � ������`��V i�!�W��"��# I��`�xph`X�0�"�H�# I�` ��` t� ��`�	)�悥���� �������! ]�`  ��`����	`� � '�`�h���P���@� � �@� !� ��`� �P�Q�R�S�T�U�f�g��e��8�4��\ ���5``�`��
�������l �W�� �%�8�&�&�
��
�&�%�� �% i+�!�U��"�0�# I����� ���l�� ���`@P a� �� ��`�	)�)��U� �8�!�X�"�g�#�_�$ �`�� �`������(� � '�@� ��@��������m��� !� ��惥�)��`���  
        ������8��������4�5` 	
���4�5`� � � �!�x�"���#�$ �!� �`��
��?�@l C�d� `� |� �� �� é ���t���8�`��` i�!�z"�8�# I��`�x�Pe`�P�Qea�Q� �P�
�	�
�P��P������P i�!��"�H�# I���P �V �����`��P �V ��`��V i�!��"�(�# I��`�xph`X� ��!���"�Å# I�����`(8H�J�!��"��# I�K�!�`�"��# I� �%�8�&�&�
��
�&�%�� �% iM�!�bÅ"��# I�����`HP �� k�`��`� �8���ݥ������]�8ݪÐ�!���4�5`�5��Å4`3������(� � '�@� ��@�x�������m��� !� ��惥�)��`��
���Å��Ål ��� $ĩ�� �ĩ ������ >� _� ���` ~� 4� U� ��`�L�!�(�"��# I�`����	)���I��iW�!��"�8�# I�`��� �	)����zą!�p�"�8�# I�慥�)��`YZY[�0A)�:����ą!i�#�@�"i�$� �  ॆI����\�!��i�A��ą"�@�# I�``� �P�Q�R�S�T�U�f�g��e �¥��� �4�5`��\���	)�P� � '�0���������Fō@�@�  !� ��� '�`���������FōA�A� !� ��懥�)��`000-./00��
��_Ņ�`Ņl gřŠŧũ ����@������ 婠�������6�M�@��� ���` �� �` b� �` �� � ��`�	)�M� ��@�:�JƝ��VƝ��@� ���Ɲ@ ��戥��� � ���i� ����@`������`123455�	)�8� ��@�'I�@)� �JƝ��VƝ��@� �
ie �@ �������`8`�8`�8`�0000PPPP�	)�H���H�B� � ���!i�#���"i�$ �΍΍΍΍悥���� �����ƍM�� ��`� ���9�M�� �� � ��`6787876�	)���I��i9�M�� ��`��4�5`�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
��ȅ�ȅl #�?�������Lԩ���� K� � �� � �� IɩE�! C��` =� �� s��`� �%�8�&�&�
��
�&�%�� �% i;�!�}ȅ"� �# I�����`8@� �%�\�&�&�
��
�&�%�� �% i;�!�}ȅ"��# I�����`��P i;�!�Ʌ"��# I���P �b �1�����? B��\ ȥei�e�e�
��
�e�f�f�
��
�f�g`��P �b ��������80( �8���
��3Յ�4Յ� �� ��K��`� ��@����`�8�����XɅ�` Z�������������������������� �����i���������������	�_�`�a���������� ������`�@� ��@�H��� ��� � ��`�8���
��`���a��� ��`��@��`  � O� 2� �� � n� n� �� �� �� �� �� �� `� {ҥ��� �� ��`�	)����=ʅ! C�恥���� ��`EFEGEF���"� �# I�`�	)����I��iH�!�H�"��# I�`�	)�B�_�	�_慥����a���A� ���`	�	�`�a`��_ i;�!��ʅ"��# I��`ph`�i�8�	)��0�)�+�)� �L�ʥ)� �̥)� *�L�ʥ)� ��`���������)�L��`��)�`��)��L�˭�)��L̭��!�q������������)�]��)�V 7ͥ#��M���!��i�" L� ������������)��#��ƈ �� ��扦�� �P���� ���B�  �`��ɐ�si	������������)�\��)�U 7ͥ#��L���!���" L� ������������)��#��ƈ �� ��扦���P��������@�  �`���v8�������������)�_��)�X 7ͥ#��O��i�!���" L� ��΀΀΀΀��)��#��ƈ �� ��扦���P��������A�  �`��ɘ�ri	������������)�\��)�U 7ͥ#��L���!���" L� ��������)��#��ƈ �� ��扦���P��������@�  �`�	)���I�����3�e��@� � ��`���!���"�"8� JJJ�0� ��!� �� �!���!� �0�!��" ��#e�#��� JJJ���ͅ$�#� j�$��)�#`	��/�8�>�0�� ����/���� :� =����`��/�8�>�0�� ����/ =� :����`���!�����"�� L�� � ����� =����`� �A��)JJJ��΅!��� !� `�0����)JJJ��.�9 � `?���� �i�)0�`��)����)�����%��i�A �� 7� Φ��P��
��w΅�x΅l `ΑεΣέ�i�� �� ��Ɖ`��8��� �� �Ɖ`��8��� �� �Ɖ`��i�� �� ��Ɖ` ���P�P� �P�
�	�
�P��P����� ��`���!���" L�8�>� ��`����ɠ�ɴ�`�!���" L��/�8�>�0�� �/����� =� :����`�/i0�/��0`���!���" L�8�>��� � ����� =����`���=�_�`�,�a�(��������H����A�@��� �������`�
�? B���`�	)�/���+� ����@�0��ɠ� ��L�Ͻ�ɴ� ��搦����`�Ə��� �@`��Y�Œ�S�]���e����8���
��`��/�a��0�8���
������ ������ ��
��/��ȱ/��� ����ő��`� �Ц���������ȱ��@� )?�A�@�� 0�I�Ȅ��i� ���Ƒ�Ɣм�`
� ���@�����`����Ѕ �	% ������ ���@�  � ��搦����`?����Ѕ �	% ���������@�  � ��搦����`���@0��i���� ��L0ѽ�8�����������@)?���@I@�@�@)?� �@
� � �A��i� ��`� �����!i�#���"i�$�@�9���/i���i�0i� ;� ����@)?���Q�Q ��  � � ��搦����`8�
���х��хl ���������D�9�&��k��Q�Q�Q�Q�QL���Q�Q�QL���R�RL���Q�Q�QL���RL���RL���\��? B� �L���a�a�
��	�a�`�_L�ѩ �^���L�ѩ� � �@�)�e �@� � ���� ����L�ѩ �B� �� ����`����Ѕ �	% ����@� ��� � �@�+)?��%�@0�� ��ɠ�e ����i�� 7ͥ#��	搦����` `�	�? B� �� �������`� �_�����L��`�	)�
�n���j�)���Ӆ ���r�)�JJJJ�!�r�)�"�!�a�F�"�`�@ �Ф���
��`�*�������@��`� ɀ��@)?�AȘ� ���Ƒ斥�)��`e �ߖ����vtrpfeYTRGC@741'%$#		
	
	���
�^�
�� ��`�, `��? B���0���@���@��,�Y !� ����`� �i� �`��
���Ӆ� ԅl �ԭ�)�
��)��`L�ʥ���� =�`� ���@�  �搦�����\0 ȩ��`� �i� �4�5`� �i���'�	)� ����ԍ@�@� � � ��暥��	�� ��`���!���" � �� �� `�	�? B���`+*)))**++� `��? B�� '� ͩ��`�	)�H���P�#Ɯ��� '��\��? B��� �ƛ�# ��`�� '����������@� !� ��`L�ϭ �]�8�1Ր�!���4�5`2g�gղ���H֓���)�t׿�
�Uؠ���6ف����bڭ���Cێ���$�o�UUeUU���������������UUUUU���j����j����j�UUUUU�������������������������UUUUUUUeUU����������������UUUV�j����UUUV�����UUVUU��������UU�����UUUUU�����UUUUUUUeUU�����UUUUU���j�UUUUU���������������UUUUU�j���UUUUU�����UUUUU��f�j��f�jUUeUU������UUUj����j��YVj����j���Vj����j�UUUj�����UUUUU�������U�������UV�UUUUeUU�����UU��V�j��j�U�UU�����UU�UU�����UUUUU�����UUYYV������YU�f�����UUUUUUUeUU���j�UUUUU���������������UUUUU�����UUUUU������UUUU�������VUV���j�UUUUUUUeUU������U�UV����f�UUUV�����UY��U�����UYU�U������U�UZ����Z�Y�UZ�����UUUUUUUeUU������U�UZ������UYUZ��i��UViUZ��i��UUUUZ�����UUeUZ��ff�UUeUZ�����UUUUUUUeUU������UUUU������UU�U�����UUU�U�����U�U�U�����U�UUU�����UUUUV�j���UUUUUUUeUU�������UZV����f�UYUf������UY�V����f�U�UU������f�UU�e����e�UU�����UUUUUUUeUU���j��UVUU���j��UUUV���j��U�UU������U�UU������UYUU������U��Z����f��YVVUUeUU��i���UeUU������UfUU��ff���VeV���ffUUUfV�����UYUUU������Y�UV������UUUUUUeUU�����UU�Yf������U��f������U�YV������UYU���������YV�����UUVUV���ffUUUUUUUeUU�����U���V����jUYYYV��Z��U�UUV�����UUU�f����fUU�VV��Zj�UU�UZ�����UU�UUUUeUU������UVYV�jf���feYf�fj���eUYV�f�Z��YUiV������YUYV��j���YUU������UUUUUUUeUU������UU�V�j����eUY�������eUU������UUUfV���f�UUVUV�Y������VV�fY�fUUYefUUeUU������UUUV����f�UUUf������UUUV������UUeZ�����UeUUV�f���UUYUV����fUU���UUeUU�����UUeYV��f���UeeZ��jjZUVVVj����Z�UU�f����f��YYf����fUYYU������UUUUUUUeUU��if��UeeV����jUeVVV�f�j��eeeV��ii�UVVVV��f�j�eeeV�f�jjVVVVV��e��UUUUUUUeUU���jfUVVVj�jj�VUeVVV�����UVYeV�jfZ��VU�U�e�f�VieVV�fZifUV�e���e�VUUYZfUUeUU�j���Ue�VV���f�VU�eV�f�Y�VU�VV�f�ffUU�fV�f�fjVU�eV�f�f��UUe��j���UUUUUUUeUU���i�UVVff�jjUUUefff���i�VYVeV�e�jfUVZef���fjVUVfV�f�f�UVUVV��j��UUeUUUUeUU�����UUUUU���j�UYYUU������U�UU�jj���eUU��Y��ZU��Yf���jfUYe�V��fffUUUUUUUeUU��jff�VUj��f�ff�eUUU�j���UUUUj����jU�UUU��i��UUUUU�ffff��j�������UUUUUUUeUU�fff�Uie�V���fj��VYZ�Ye�V�fVe���fif�eUef�Zf��U�VVZ���j�UYU�������UUUUU��
��!�+�3�;�C�K�S�[�c�k�s�{݃݋ݕݞݪݷ����������� �	���+�=�J�\�( ��)** 8X56789:$0$"X$�$D&0D!XD&�D  d!&0d&Xd##�d&8! P !H(!	H8&^HP	H`]^]^`x!
H�]^]^"
H(
H8&]^]^HP" H`&^"Hx "	H�&^8!&^%!^ !	Pij t&"^^ !^j�!&^%!^"��������������������
���ޅ��ޅl �޶�?�E�K�`����ߩ� ������ ���`��� ��`�`�	)�)�&` ߠ ��ޅ!� �"��ޅ# I�����`_ac`bd(Px ߠ ��ޅ!� �"��ޅ# I�����`� � � �!�(�"�7�#���$ �`� � �H�!�(�"���#���$ �` ��` '��`�� ������ ���`��� z�`�]�� �4�5`�]�`�	)�)�` ߠ ��߅!� �"��ޅ# I�����` ߠ ��߅!� �"��ޅ# I�����`eg_fh`  �� �� ��`��
��4��8�5`����������������������������� � �!�"���#�$ �` L�!JJ

�!�#JJ

�#�#8�!JJ�%�%�$8�"�&�&� � ���%�� =��&��`�"�}���")��q���!�����JJe���` 0`��� P���@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^_____`````aaaaaabbbbbccccc�i0���`��!� �"� �#� �` L� ��7
�� ��/���0� �/�!�# ��/�" ��/�% ���#�� =� ��!�#�"��`��%��&`�/��0`�%��&`���`�������<�� ���^`� ��`�  I����I�%��`� �#�!��"��#e"�#�!��`� �#�$�!��"��"�!�#���$`� � ��� )@�� � �� �`��@����
�'� �(����!���" L��%��& �� � ��/�%Lx�%�/ �� ���'� =��%��&�
�'�(��`�
����/���0` �����������������������������!)
� �$���" L� ���%��&��@����
�!� ��"�@
�� ��/�-���0�.� )�� �1���$�_ �� �'�(� �/�# m�#
&(�$��'�# ��#�%�1�(�'� �(� �$ �� ���!�˥'�# ��#�%�1 =��%��&�
�!�"Т` �� �/�# m� ��#�% �� ���1�!�� =��1��%��&�
�!�"��`�� ��`�/�/����0`�� )
�� ���+���,l+ '���(�?�-�/�.�0�8�"�)��
��L� U�*��e
��0e/�/��0`�-�/�.�0�"8��) U�*L�-�/�.�0�"�) U�*��L� �*�)��*e
�*��0�)��`�� )�,� ��#jjj)���#

)0��#JJ)��#***)�#� `�4�!�8�H�
����2���3� �1�2=��)����� �#=����#)�#���� h�`�0?����4��H��D��@��<����6���/��0��%�8�>�&��(� � �%�/ �������%i0�%��&�(��`� � �/�#��`��!����"��0�$��`� `� � � �* �C�D��� ���A�B`�
���܅��܅� ��(�)ȱ�*ȱ�+� ȱ�,ȱ�!�+�"�,�# I�+i�+�)��(�)� �+�,i�,�*��`�	���0�� �`����������������������������xآ��� � ���&  t橠�  � � � � � �V�W�[�Z�]��Y��X� ��5�� ��ťm���ejj����5� ��Lo� �� �� F� �� ��L@��� ��� ��������������`�5� � �5 `�4���0�? B�  � �� ?� ��`� �� ��0��` �������������������������� �%�F�&��/��0� �%�/ �� ��%ɰ��&�\��` ��%� �6�6� �7� �!� �"�6 `������`�4���& �4
�������� � �/�*���@�0�0�) ���# �� ���)�0����)�) ���# ���)� ��Lc� ��ɍ& `������������������������������������/H�0H�4
��������#�!�!��i����!�� � �� ��/ �����
� �� :�L��h�0h�/�/i�/��0�*�*��� �*�0�/iX�/��0� `�/i.�/��0`�4
��W��X�l  � � � � � � �� � � � � �� � � � � �� � � � � �� � � � � �.���Nŀ�D��������>������.������~������>������Ė������*�)�͞q�J�"�9�L�;����٦f����©ª��x���ܭƮ��:�����ų��#�-���=�����H�H�H��� V� ���h�h�h@ ���9�=�>ȱ9�O� �@����0���@�OJ��?� �@�@��� �* ���`��� ��� �  �ޥ?
��C�9�D�:`� �@�@� �@�@����>�
�=�>��`
��C�9�D�:�
��9�;ȱ9�<��� ��C�� U�L�� ��L�� �� 0]��;�OJJJ���� ��C�Bȱ;�3�

��3� �O)�6� �� �!JJJJ�$�)pJJJJ	�0 �� �O ��`�@�-�>�����k�L��*��$8�'�$���)�* �� �`� �-�$ �� �`�*���'}$�$����)�* �� �`�-�O�O �� �� �`�*�Ž$8�'�$��!)�$L��!)�$���ǽ)�* �� �`�*� �� �`�@���)��O�0��)pJJJJ	�0�

��)�%�38�O�3��6� �3�6�3� �6� `�3eO�3���6�6��ީ�6���3��~i�@�

���� `�O���@�-`
eOe@����O��@)�*�JJJJ�'�O�-`��;���e`���ȱ;������.�@���*��� ��� �  `��ý	��	��L����ȱ;��	�L����ȱ;�L��
q;e@�O����Oȱ;��@�L��i���A�A05

����A�+� � �L�,�N)� � �M�-� � �.� � �C�C�c�N�S)x�OJJ�O�L��M�C��?�N0&�L8�O�L�
�M� �L�M�L� � �M� � L��OeL�L���M�M��ܩ �L�C�� � � �B0

����B�?�( �@�) �D�A�* �D�	�D�� �* `xy� ..< �l ���=���)���7�w���a�����e�������k�A�d2�	}T� T� T� P �	}T� T� T� P �	�}� }� }� 0  .	@T� T� T� P ��� � � P ��� � �q P ���q �q �q 0  �xq_ q_ ke  @   �  #�#("�#(#�#("�!�#�#("�#("�"!�"#�"�"\!�#�"�"\"�#�#("�#(#�#("�  !�!�!T!�!�!�!T �!�!�!T!�!T! �!!�!}!. �!�!}!.!}!T!    #("�#�  ���d0�0��0��1T�1.0�.T( @   �0�0��0��1T�1.0�.�( @ 0��0��0��0��0��0���( @ 0��0��0��0�T1.0�.�( �  T 0�0��0��0�0��0��( @   �(C(B�C�C(B�B\BB�C(B�C�C(B�B\B�BC�B�C�B�C�B�C�C(C�B�C�B�B�B\B@ C(B�C�C(B�B\BB�C(B�C�C(B�B�C(C�  ��������@� ����@���� ��� �� �@����� ������@����!����� ������� �����d2����� ��� �� @������ ������( }T@� ������� �x���x��x�h   �@"�!�!�!�"�!�"�!�"�!�!�!�"�!�"�!�#X"<"�"<"�!�!�"�"<!}!�"<"�"�"<#X"�!�!�!�"�!�"�!�!�"�!�"�#X"�"�!�#�"�"�#�#�"�#X#�"�#X"�#X!�!�B�  g���.	@h	.@	h�	�A�   �@ �  \ B�   �����}	���A� ��I���@� ���A ��@� ���  6@� ��� @� ��� ������� ������� �������  � ����� @ �����  �@<�}�B<�<�<B��X�XC��\�\B�  }����F ���@� ������� � � �� � �	.�1   ���@� ������� � � �� � �0�    d< � X � < � \ � < � � � � � � �   =�=��@	� 	� 	� 	� !T!�	} 	} 	} 	} @0 	� 	� 	� 	� !}�<	� 	� 	� 	� T  �0 	T 	T 	T 	T !!T@  � �}	T 	T 	T 	� 	} 	} 	} 	� ��d 0 	� 	� 	� 	� � � 
< 
< 
< 	� T  	} 	} 	} 	T . }   �@T}  C�C��@�!��� � �!�h} � �!}�h  @}�}!�  �!��� � �!�h} � �	} }�h@ @}��!�  �!h}@ @ �!@ h h!h � �h!@  �!h}@ @ �!@ h h	 h�� �@}!h    /�/��@	� 	� 	� 	� 	� 
< � 	� 	� 	� 	� 	� 
< � 	� 	� 	� 	� 	� 	� T 	} 	� 	� 
< � � 	� 	� 	� 	� �<� 	� 	� 	� 	� }} 	T 	T 	. 	. }!�	� 	� �\� <   ���@	T 	� 	T 	� 	} 0 	} 	� 	} 	� 	� 0 	T 	� 	T 	� 	}  	}  	} 	� 	} 	� 	� 0 	@ 	� 	@ 	� � 0 	@ 	� 	@ 	� 	 0 	@ 	� 	@ 	� �  �  � 	@ � 	@ 	 0   �����F	} 	} 	T 	@ 	} 	} � 	} 	} 	T 	@ 	} 	} � 	} 	} 	T 	@ � 	 	@ 	} 	T 	@ 	} 	� !}  	 	 � � 	 	 } 	 	 � � 	 	 } 	 	 � � � � � 	 � � 	 	} !    �����.. �.}.� � �ThT.T��A}@  �@� � \ � � � < � � ( � � b\   %���  ��� � � � ���@	} 	} }@� ��� � � � ���@� ���  � @T	} 	} 	} 	} }T@�� ��!@  	} 	} 	} 	} �}��A  }T	@ 	@ 	@ @� � ��� ��!@  � � ��� � 	 	 1@   �@ ���������������<��������X�X�X�  ��X�����X�������X�X<�<�<�<�X�#X �<���������X������<�<�X�X��X"�  �����	.	 � ������@T@��`� ���& ��� ���A�B� � � �* �C�D� � �< ����E�[�F� �G�H��I��& ��I���I y� "��G����H����i<���`�E��E`�E�G�>�]�:��8�G ��i0�J�i �K�G�����J����J�i0�J�K�i �K���G���  ���G�a�.�]�*�D �����ȑ���� ��i0��i �����E� �G�_��a�Ș J��G�a����G`�G`�F��F`�H�K�]�G��8�H ��i��i ��i0�J�i �K�H�����J����J�i0�J�K�i �K���H��� ���H�a�0�]�,�D ���ȱ����'��� ��i0��i ���ߩ�F�H�a����H`�H`



}g��J�h�i �K�J��� ��k�e��i ���J���`� � ��@�� ��������`H)��*��hJJJJ�
ei@}:��` 0`��� P���@p��      

�� �_�� � �����`� �/ �m�m� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������)� � �