                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��������������������������������������������ꫪ��ꫪ��ꫪ��ꫪ��ꫪ��ꫪ��ꫪ���*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �������������������������������������������                                  �����                                  ���*             �          ��      ��«*            �_          _�      ��«*      ��?   �U?          WU?      ��«*     ����  �U?         �WU?      ��«*    �UU��?  pU?         �WU?      ���    �WUUU�� pU?         �WU�      � �    |UUUUU�? �U?          _U�      � ���   _UUUUU���U?          \U�     �����  �WUUUUU���U?          pU�     �����  �UUUUUUU� W?          �U� �  ���*  �UUUUUUU�? W?          �U� |�  ��«*  �UUUUUUU�? W?           W� WU ��«*  �UUU��_U�? W?           \U?�UU ��«*   WUU? �U�? W?           \U?�UU ��«*   \UU �WU� W?           \U�pUU ���    �� �WU��U?           pU�_UU � �     p�  WU��U?           pU�_U� � ���    p�  WU��U?           pU�_U� �����    p�  WU��U?           �U�WU�  �����    p� �WU��U?            WUUU=  ���*    p� �U���U?        �?  WUUU=  ��«*    p� �U�?�U?       ��� WUUU  ��«*    p� pU�?�U?       U�? _UU�  ��«*    p��_U�pU?  �  �_UU� \UU�  ��«*    \���WU�pU? �U�  �UUUU\UU�   ���     \U�_UU� pU? |UU |UUUU\UU�   � �     \UUUUU? pU? _UU? _UUUU\UU�   � ���    \UUUU�? pU?�WUU= WU�_U\UU�   �����    \UUUU�� pU?�UUU��UU�_U\UU�   �����    \UUUU��pU?|UUU��U�?U\UU�  ���*    \UUUUU�pU?_UUU��U��� \UU�  ��«*    \UUUUU�pU?_UU��U��5 \UU�  ��«*    \UUUUU�pU?_��W��U�  \UU�?  ��«*    \U�UU�pU?W� _��U�    \UU�?  ��«*    WU��_U�?pU?W= _��U=    pUUU�  ���     WU |U�?pU?W= _��U=    pUUU� � �     WU �U�?pU?W= _�W=    pUUU� � ���    W� �W�?\U?W=�_�W�    pU�U�? �����    W� �W�?\U?W��W�W�    pU�UU� �����    W� �W�?WU?W��U�W� � pUUWU����*    W� �U�?WU?W�U�W���pUU_U���«*   �U� pU�?WU?\UUU�_U���?pUU_U�?��«*   �U� _U�WU?\UUU�\U���?\UUsU����«*  ��U���UU�WU\UUU�pU�U�\UU�UU���«*  �UU��UUU�WUpUUU�pUUUU�\UU�UU����   �UUUUUUU�WU�UUU� �UUUU�\UUWU�� �   �UUUUUUU�WU�UU�� �UUUU�\UU\Uճ ���  �UUUUUU��W�  WU�? �UUUU�\UUpU������  �UUUUU��� W5  \��  UU�?\UU�U������  �UUUU���? |  ���  �W��_UU�Wհ��*  �UU�����  �  ��    ��  WU� W5��«*  �����?                   _U�  �?��«*                           |U?    ��«*                           ��     ��«*                                  ���                                   � �                                   � ���                                  �����                                  ����� ���?              �              ���*�����            ��             ��«*_UUU�            �U       � ��  ��«*�UUUUU?            pU�     ����� ��«*�UUUUU�           ?p��    ���W�? ��«*�UU�U�          ��p���    |�_U�� ��� �UU��_�   �?    |�s��W    _UUUU�� � WU= |�   |�    _���_U    \UUUU�� ���WU= ���� |�   WU��_U    |UUUU�?�����\U= ����\���\UUUU� � pUUUUU?�����\U= ����\���?pUUUU��U��UUUUU����*�= ��W�|� _U��UUUU= _UU=�UU�WU���«* p= p�W�p��UU��UUU��UUU��UU_U���«* p= \�T�p=pUU��W�? pUUU��U� \U���«* p= \�W� p=|UUU W�  \U�WU�W� \U���«* p��W�W� p=\UUU= W�  W�\UW�|U����  p��U�\� p=\U}U= W�  W�|UW�p��� �  pUUU� p� p=\U�W= W=  W� \UW���?� ��� \UUU� �� p=\U\? W=  W? W�W��� ����� \UUU= ��p=\U� W=  W��U� W�   ����� \UUU ��p=pU�  W= �U�U? W�   ���* \UU� ��p=�UU  W= �UUU� W�   ��«* \UUU� ��p=�_U�  W= �UUU�  _�   ��«* \UUU�?��p= pU� W= �UU�  \�   ��«* \UUU�� �p= �WU W=��UU=   \�   ��«* \UUUU� �p=  \U= W=��UU �\�   ���  _U�_U��p=  pU��W���W� \�   � �  _�AU��p=  �U��W�WW��_5\�   � ��� W} �U�W\=  �U��U�WWU��W5\U   ����� W �U�W\=��U��UUU=WU�U�pU   ����� � �U�W�\=��_U��UUU=\UUUU�pU?   ���* � �U�W�W=\}UU��UUU=\UUUU�pU?   ��«* � �U�W�W=\UUU��UUU�UUUU�pU?   ��«* � pU�W�U=|UUU��UUU _UUU5pU?   ��«* �? |U�WUU=�UU���UU� �WU�p�   ��«* W�?U�_UU=�_U� _U=   ��? ��    ���  W��UU�\UU� ��?  �U             � � �W�_UU���W���    �              � ���WUUUUU���U                     �����WUUUUU� �U                     �����WUUUUU�  �W                     ���*WUUUU��   �                     ��«*WUUU��?    <                      ��«*WU����               ��     ��«*������                






(    ��«*                      




 
(    ���                       




 
(    � �                       �

��*    � ���                      
 

 

(    �����                      
 

 

(    �����                      
 




(    ���*                       ��    ��«*                                  ��«*                                  ��«*                                  ��«*                                  ���                                   � �                      �
��� �
��
 � ���                     
(�� ((��� �����                     
  
 
(� (  �����                     
  
 
(� (  ���*                     �
 
�((� (  ��«*                      ( 
��(�
 (  ��«*                      ( 
�(( (  ��«*                     
( 
�((( (  ��«*                     �
 �(    ���                             �    � �                              �    � ���                                  �����                                  �����                                  ���*                                  ��«*                                  ��«*                                  ��«*                                  ��«*                                  ���                                   � �                                   � ���                                  �����������������������������������������������ꫪ��ꫪ��ꫪ��ꫪ��ꫪ��ꫪ��ꫪ���*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��«*��� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����������������������������������������                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �    UUUUUUUUUU         @UUUUUUUUU    �   @                           @    �   @                           @    �   @��*(��         
����
(�J    �   @�� (
�         
��� (�@    �   @�� (
�         
��� (�@    �   @��
(��         ��*�� �
�@    �   @�� (
�         
���((�@    �   @��  
�         
���((�@    �   @���*� ���         
����"(�@    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �   @                           @    �    UUUUUUUUUU         @UUUUUUUUU    �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �    UUUUUUUUUUUUUUUUUUUUUUUUUUUUU    �   @                             @    �   @                             @    �   @                             @    �   @�� *�* �*�* *�����* *   �� @    �   @ 
���� �������� ���� � 

@    �   @ 
���� � � ���� ����

@    �   @ 
���* �*� �����* �*����
@    �   @ 
���  �� ���"� ������
� 
@    �   @ 
���  �������� �����

@    �   @ 
 *� �*�* *�����* *�

� @    �   @                             @    �   @                             @    �    UUUUUUUUUUUUUUUUUUUUUUUUUUUUU    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �   @                             @    �    UUUUUUUUUUUUUUUUUUUUUUUUUUUUU    �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �    �        ��*��
�                �            "          �*       �    "
��
�   "    *�
  
�  ( 
    �    �� "   � �
      � "  �     �      ��
�   �"        ��*       �           "   "             �      ��
�  � "    ��
 �
��
�      �                                      �                                      �                                      �                                      �                                      �����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����������������������������������������                                      �                            �  @QEQEQEQEQEQEQ  @DDDDDDDDDD �  PUUUUUUUUUUUUUUUUUUUU    �  T                      @D�OO�O��tD �                         �1�1� �  �
���*�* �����  @D�tO�tO�GD �  � (
���  <<<<<<<<<<   ��1� �  � ( 
���  <?<?<?<?<?  @D�tO�tO�GD �  �
( 
�*�
 �<�<�<�<�<   �1�1� �    ( 
�"�  <<<<<<<<<<  @D�O��O��pD �  � (
���  <<<<<<<<<<    �  �
�����* �����  @DDDDDDDDDD �                         ����?� �  T                      @�tO�tt�DOG �  PUUUUUUUUUUUUUUUUUUUU   �1�1� �  @EQEQEQEQEQEQE  @�OO�Ot�O�D �                           �1=1� ��������������������������@�tOw|t�DOG ��������������������������
 ���1�? ��                        
@DDDDDDDDDD ��                        
  ��                        
@DDDDDDDDDD ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@          ��                        
@          ��                        
@  �
��  ��                        
@  � ((  ��                        
@  � 
(((  ��                        
@  � 
(�  ��                        
@  � (   ��                        
@  � �(   ��                        
@          ��                        
@          ��                        
@�������                        
@<<<<<<<<<<��                        
@<?<?<?<?<?��                        
@�<�<�<�<�<��                        
@<<<<<<<<<<��                        
@<<<<<<<<<<��                        
@�������                        
@          ��                        
@          ��                        
 UUUUUUUUUU ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@          ��                        
@          ��                        
@��*(�� ��                        
@�� (
� ��                        
@�� (
� ��                        
@��
(�� ��                        
@�� (
� ��                        
@��  
� ��                        
@���*� ��� ��                        
@          ��                        
@          ��                        
@   ��   ��                        
@   <<<<   ��                        
@   <?<?   ��                        
@   �<�<   ��                        
@   <<<<   ��                        
@   <<<<   ��                        
@   ��   ��                        
@          ��                        
@          ��                        
 UUUUUUUUUU ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@          ��                        
@          ��                        
@��
�* ��                        
@��(
�� ��                        
@���
� ��                        
@��(
� * ��                        
@��(
 � ��                        
@��(
�� ��                        
@���
(�* ��                        
@          ��                        
@          ��                        
@  ���  ��                        
@  <<<<<<  ��                        
@  <?<?<?  ��                        
@  �<�<�<  ��                        
@  <<<<<<  ��                        
@  <<<<<<  ��                        
@  ���  ��                        
@          ��                        
@          ��                        
 UUUUUUUUUU ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@��                        
@DDDDDDDDDD��                        
@��                        
@        D��                        
@�
**�*��                        
@

 (
�D��                        
@*
  ���                        
@�
  �D��                        
@

� � ���                        
@

  �D��                        
@

  ���                        
@

 (
�D��                        
@
�
**���                        
@        D��                        
@QUUUUUUUU��                        
@        D��                        
@�?�?�?�?��                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@������                        
@�?�?�?�?D��                        
@�?�?�?�?��                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@������                        
@�?�?�?�?D��                        
@        ��                        
@DDDDDDDDDD��                        
@��                        
@DDDDDDDDDD��                        
 UUUUUUUUUU ��                        
            ��������������������������
            ��������������������������            �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���*      �?�?      �
    �
    �
    �
 
�  � �  � �  � � 
 � �  � �  � � � 
  �
    �
    �
    
                   
     PP            
   PUpp  P       �  
 P �ppPUp          
 p p pp�p         
 p ppqp p         
 p ��]pp         
 p p ��p         
 p pU p pU         
 pU�  pU�      �  
 �    �          
                   
                    �
    �
    �
    ��  �  � �  � �  � �   � �  � �  � �      �
    �
    �
     �
    �
    �
    � � �  � �  � �  �� 
  � �  � �  � �  
   �
    �
    �
  
                   
     PP          �  
 P   ppPU           
 p PUpp�P         
 p �ppp p         
 p p pqpp         
 p p�]�p         
 p ��p p          
 pUp  pUp       �  
 �pU  �pU        
   �    �        
                    
                  � 
�
    �
    �
    � � �  � �  � �  �    � �  � �  � �      �
    �
    �
     �
    �
    �
      � �  � �  � �  � �  � �  � �  � �� 
    �
    �
    �
  
 P                 
 p     PU          
 p   PP�P       �  
 p PUppp p          
 p �pppp         
 p p pp�p         
 pUppqp p         
 ���]pUp         
   p ��pU         
   pU   �      �  
   �              
                   
                    
 �
    �
    �
   � 
� �  � �  � �  � �  � �  � �  � � 
    �
    �
    �
     �
    �
    �
      � �  � �  � �    �  � �  � �  � � �
    �
    �
    �� 
                    
 P     PU          
 p PU  �P         
 p �  p p       �  
 p p PPpp          
 p ppp�p         
 p �ppp p         
 pUp pppUp         
 �pUpq�pU        
   ��]  �         
     �          �  
                  
                   
  �
    �
    �
    
 � �  � �  � � � 
�  � �  � �  � � �
    �
    �
    �
     �
    �
    �
     � �  � �  � �  � �  � �  � �  �  
�
    �
    �
    � 
         P        � 
   PU    p          
 P �  PUp         
 p p PP�p         
 p pppp p       �  
 p �pppp          
 p p pp�pU        
 p pUpqp �        
 pU��]pU          
 �  ��          
                   
                 �  
                   
   �
    �
    �
  
  � �  � �  � �  � �  � �  � �  ��  �
    �
    �
    � 
    �
    �
    �
  �  � �  � �  � � 
� �  � �  � �  � 
 �
    �
    �
   � 
                    
   PU    P         
   �PP  p         
 P p ppPUp       �  
 p ppp�p          
 p �ppp p         
 p p pqpp         
 p pU�]�pU        
 p ��p �        
 pU   pU           
 �    �        �  
                   
                   
    �
    �
    �
  �  � �  � �  � ��  � �  � �  � �  �   �
    �
    �
     ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WuU5 �_U pU�  �_� <�{5 ��k� W��� \WU� �WU? W�� �� ���? �_�      ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WuU5 �_U pU�  �_�  ܫ7  ��7  _��  W��  W��  ���  ��� �W�� ���      ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WUU5 �_U pU�  �_?   �?   ��   �_  �U  �U  ��  W�  �� �� ��� ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WUU5 �_U pU�  �_?   �?   ��  �W <�U� <�U� ���� ���� ����  ���    �  � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \U]� �U�?  WU ��� \�7< W��� W��� �U�5 �U� W�� ��� �WW? ��       � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \U]� �U�?  WU ��� ��7  ܪ�  �W�  �_�  ?�  ?��  ?�?  _� ��       � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \UU� �U�?  WU  ��  �7   ��  ���  �U�  �U�  ���  ���  �W�  ��� ���  � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \UU� �U�?  WU  ��  �7   ��  ���0 �U�< �U�< ��?? ��?? ��?? ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���ة�� ���  ��� � � � � � � �ߍ& ��"  �آ t ���� �� �� � ����� ��� ��XL �H�Z� � �P0� � � � ��  ��z�(h@H�' )�	� � �# �$ �% hX@                                                                                                                                                                                                                                                                                                                                                                          �ȩ��  �� 6� 	ة 3�:���  ٩�� �
��  v����� ����� �� Bɩ � [� q� {� �� � �� 5� V� y� � �ϭj �k � �n  3� V� y� �ũ �s  p����� ��  b� i� |� ��L� �ɭs ���S �����& v������� Ԁ���� #ŀ���� Bŀ���� aŀ���� �� �� �ɀ���� �Ā���Ы �Ā� �� C� a� �� �� x�L\�Hڢ
�f �0��0��0��0��0��0ʎ� �h`H�Z��� � � ��! ��  ��	 ���
 �
 � �	 �  7Ĭ
 �r� ���
 ��h� ��� �
 �
 � �	 � � � ��  ��!  7�� � � � � � ��! ��  ��  7Ĭ �D� ��L� �� �ĭ
 � ��  �	 � � � ��!  �ĭ	 i�	 �  7ĭ � ��! ��  �ĭ 8�� �  7ĭ �\� ��L��z�h`xH�Z� 
���ڍ 轾ڍ �  � �! � � �J� ��� � JJ��- �� i� � i � � � � �Ȁ�� � � �
�! � �L\�z�hX`H� �  7ĩ�� h`H�Z�/���� ���� ��z�h` ������ �������� �� �� U� ?� ��` ������w �����p��� �� �� G� ?� �ɀW 	�� �P��� �� �ʩ� � �ɀ8 S�� �1��� �� �ʩ� � �ɀ ��� � �ʩ� � �ɀ���s `�g � �>�g ��I�� �g m m i)�0im� mo mp ��  "��� �ֈ� �� ��`H��o � �p  ?�h`H�f �� ��h`�Z�o ڮp ڮn ڭk �l  U� �ˠ �(mo � �,�(� ȱ(mp � ���  �����
Ș��̩��� ��n ��p ��o z�`H�Z�k �l  �ˠ �(mo � ȱ(mp �  "�����z�h`�Z�k �l  �ˠ �(mo � ȱ(mp �  �����	������� z�`�Z�o ڮp ڮn ڭk �l  G� �ˠ �(mo � �+�'� ȱ(mp � ���  �����	���ͩ��� ��n ��p ��o z�`�Z�o ڮp ڭk �l  �ˠ �(mo �0:� ȱ(mp �  �����	���ܩ��� ��p ��o z�`�Z�o ڮp � �ˠ �(mo �� ȱ(mp �  �����	���ܩ��� ��p ��o z�`�Z�o ڮp � �ˠ �(mo � ȱ(mp ��  �����	���ܩ��� ��p ��o z�`� ٜf �g  4� J� `� �� �� ��������0��� �� JȀ���� �� JȀ���� �� 4Ȁ����� �� 4Ȁ� ��`��� �� �2� �f  �`��� �� �2� �g  �`��� �� �d� � �٩� �n� � �٩� �x� � ��`��� �� �d� �� )�  $ڭ�  ڭ�  ک� �n� �� )�  $ڭ�  ڭ�  ک� �x� �� )�  $ڭ�  ڭ�  �`� �� �� �� �� �� �� �� �� �� � �d�� �� �� ����$�� �� �� �f �g �b�m `�` �a �b �c �d �e �h �i �j �k �n �s �� � � �v �� ��`H�  � �� ��h`ڭ  � �� ���`H ������ ��h`H ������h`H� h`ڮf �qۍ �`�Z� � �� ���z�`��� �� �D� �f  �`��� �� �� �b )�  $ڭa  ڭ`  �`��� �� �%� �� )�  $ڭ�  ڭ�  �`��� �� �_� �i )�  $ڭh  �`H ��mj mo mp m` mf mh )�0� �j h`H�Z�n H� �n �j 
����i� 轗�i�  �ʭj �l  d�h�n z�h`H�Z� H� H� � �
i� �


i� �a�  $���������h� h� z�h`H�Z�m H�q � �r � �a�m �k �l  d�h�m z�h`H�Z ������o �����o �����p  ?�z�h`H�Z�o �p  �ӭ �q � �r �k �l  d�z�h`H�Z� � � �  �ˠ �(
m � ȱ(


m � �m �  $�����z�h`H�Z�l 
���& ��' �n 
��&�( ȱ&�) z�h`H�Z�b �� 0N��a �� 0D��` �� 0:�b �� 0S��a �� 0I��` �� 0?�b �� 0M��a �� 0C��` �� 09��L u� �� �̩d� �� ���� ʩ�� �- �̩d� �� ������� � u� �̩d� �� ������� z�h`�� �� �� �� �� �� � �� �� ����`�� �� �� �� �� �� � �� �� ����`�` �� �a �� �b �� `�` �� �a �� �b �� `�` �� �a �� �b �� `H�Z�
�� �� � �Lfͩ � 4� J� `� �Ȉ�A� � �A8�7� �P� �ߍ& � �<�  �� $�������� �̀���� �̀��� j̀���� j���дz�h`Z�
��D�& ȹD�' ��� i7�&z ��`H�Z8�7� � �a�
� � ��A8�7� ��a� h`H�A8�7� � �a�	�0� ��Z8�7� ��a� h`H�Z��)	@�& � �ۙ0 ��0���h�. �N�/ � � ��ڍ* ȹ�ڍ+ � e� Ϲ0 �* ȹ0 �+ �� �Ω 3�:� ���0�� �. �. �C�. Z� �Aۙ0 ��0��z�:Ъ�ߍ& z�h`HZڭ. i�, �/ �- � � �m. �h�*�,������* i�* �+ i �+ �, i0�, �- i �- ����zh`HZڭ. �, �/ �- � � �m. �h�*�,������* i�* �+ i �+ �, i0�, �- i �- ����zh`HZک�� �� �. i�, �/ 8�@�- �- � �	�, 0�00�, 8�0�, �- � �- � �ڭ, i� �$�f )�JJJJ�  $ڭf )�  $��zh`H�Z�d �0b� ��  b� i� �� �� �� �ͭ� � ��� ٭c )�c �d �e �n �� �v �v ʈ� ��v �w �x �y  �� �� � �� 5� q�z�h`H�Z�t �u � � �
��v ���ȹv )��	H� � �h���ܭt � ��u � � /� 5�z�h`H�Z� �� �� �Т��� >������Z�
��v � �v � �
�� �� ȭ �� z�� �ψZ�
�� �� ș� z� �� �� �v �� �� �� ��z�h`H�Z�

��6�



���6��) �6��* �6��( z�h`H�Z�* z�h`H�Z� ڢ� >�����b�  �� �� 3Ѣ� >�����a�  �� �� 3������z�h`H�Z���  �� $�����z�h`�Z�P���� ���� ��z�`�n ��� �n `�n ��:�n `H�Z�k 

mn �� ��m` �` �a i �a �b i )�b �z�h`H�Z�k 

mn �� ��mc �c �d i �d �e i )�e �z�h`H��f i�f �h`H�f � ��8��f �h`H��g �0��g ��g i�g �h`H�g � ��8��g �(h`H��h i�h �i i �i �h`H�Z� �0�� � JJJ� � 
m � �� � �	� 
�� ��� � �v  �v z�h`H�Z� �0�� � JJJ� � 
m � �� � �	� 
�� ��� I�� �v - �v z�h`�Z� �0�� � JJJ� � 
m � �� � �	� 
�� ��� � �v - � ����� z�`H�Z� �0�� � JJJ� �� � �	� 
�� ��� � �t  �t z�h`�Z��0�� �JJJ� �� � �	� 
�� ��� � �t - � ����� z�`H�Z� ��  b� i� �� �˩J� �c� �  �ڊ�I�:� �� 3����� � �ө�� �  ��z�h`H�Z� � � �  ������m � ��a�  �� $���������z�h`H�Z�
i� �


i� z�h`H�Z b� iש�)��&  �ɩ� �� ��� � �� v���� �� �ɩߍ&  Y� ��z�h`� �� ��  b� iל � � � � � � � �� �� �ߍ& `�� ���Q�� ���.�� � b׭� �� � �  Y֭� � i׭� �� � �  ���� �� �� � ��� �� �� � �խ� ���.�� � b� i׭� �� � � � �  	��� �� �� � ��`�� �Ս� ȱՍ� ȱՍ� ȱՍ� ȱՍ� )
��(��� �(��� Ȍ� �� �� �� � �)�� ���� ���� � ��� � ��� ���� �� ��`�� ��� ȱ�� ȱ�� ȱ�� ȱ�� )
��(��� �(��� Ȍ� �� �� �� � �#� ��  b� i׭� �� � � �� �� � � `�� ��� ȱ�� ȱ�� ȱ�� ȱ�� )
��(��� �(��� Ȍ� �� �� �� � �)�� ���� ���� � ��� � ��� ���� �� ��`H�Z�� )?	@�� �� 4��-� �� �� �ܪ�� )@��J��� �� Ȍ� ������� �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� �骭� )@��J��� �� Ȍ� ������� �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� ������� �� �� �� � �� � �� z�h`� �� `� �� ``���� ���� ���� ���� �� �� ��� ��  � �� Y� �֩��� `���� ���� �� ���  �� 	ש��� `� ��� �!��� �� ���  �� 	ש��� `�"��� �#��� �� ���  �� 	ש��� `�$��� �%��� �� ���  �� 	ש��� `H�Z� � H� H�
� �� �  �h� h� z�h`H�Z� � H� H�
� �2� �  �h� h� z�h`H�Z� � H� H�
� �F� �  �h� h� z�h`� � � � � � � � � � � �( �) �* `� � ������ � `� � ɪ�� � � `Hڪ���




� ��) �& �h`H�Z ��
���ڍ$ ��ڍ% � �" �@�# � � �$�"��(���" i0�" �# i �# �$ i(�$ �% i �% ���Ωߍ& z�h`��� �� �� �  �٩�� �� �
� � �٩�� � @��0��� ��C��0��`H�Z� �@� � � � ����� ���z�h`H�Z
���ڍ ��ڍ � ��$��a��b��c��d�8�7�  $�Ȁ�z�h`H�Z�)�JJJJ�  $ڊ)�  $�z�h`xH�Z� �a��$��b��%��c��&��d��'���� ��� �� � �J� ��� � �- �� Ȳ- �� �� ��� � z�hX` GAME  OVER $PAUSE$LEVEL  :$HEIGHT :$G T C$ �C��ڠڦگڸڶ � �  � � �   @ `��9�򥫧d����9�򥫧d����9�򥫧d����9�򥫧d��֬֬ƭƭN�N�ƭƭ֬֬ƭƭN�N�ƭƭ֬֬ƭƭN�N�ƭƭN�>�>�N�.���.�N�>�>�N�.���.�N�>�>�N�.���.�F8-$$      		      f g        �� � �� � �� � �� �� �� �� �� �� �� �� � q� �� �� �� �� �� �� �� ��T�.�� �� � ?� ?� �    �� � �� � �� � �� �� �� �� �� �� q� � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �    q� d� _� d� � � �� � q� � �� � q� d� _� d� � �� K� T� _� T� _�    ���.����� �.�T�}����� ���}���������:��� 0�    ���.����� �.�T�}����� ���}���}��.�}�T�}� �   ��}����� �:�����\� ���}�������.�.���}�    �� �� ��    _� T� K� ?� ?� � ?� K� T� _� _� T� K� K� T� _� T � � _� T� K� ?� ?� � ?� K� T� _� _� T� K� K� T� T� _� � � _� @�    _� 2� 8� ?� G� K� T� _� � � _�    �� /2�   �
	�
�
�
	�	�

		���H���  Rݾ�/�  �ޣ�iߣ�  �߳߾���������    �      �    �   �  �  �   �      ��  � ��   �  �   � �   �   �  �  �� �   �      � �   �    �      �   �     B�J�R�Z�b�j�r�z��������������������������������������������
�
dnx� � �  0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            W� �}�