�7�b�����r�	!��������       �      �      �   �  �   �  �  �1  �  �1  � ; ��  � ; ��  � �� �� � ��0o3 � ��o� � ������ � ��7� � ����3 � ��o� � ���� � ����?� ������� ��V�� ���7�� ���7�� �����7�� �>�V�� �33_�� ?03�� 03 ?� 03 ��� ��������       � ��������          	!��������  0    �  �    �  0    �  �    � ��
   � �*   � �*   � �* � � �� � � �� �� 0 0 �
� ��� �*� �� �*� ��� �*� ��� �� ��� 0� #� ���� #����k�� +�33�{�� +����k�� �� ����� �����k�� �������� �������� �������� �����k� �������� ��     � ��������       � ��������          	!��������  �    �  �   �  �  � ���?? � ����� � ��� � � ��� �S� �� WU� ��WU� ���P� ����� � ���� � ���_U� ��� <L� ��� � � ���� � ���� � ï�� � �� � ���  ?<� �������� �����3� �����? � �������� ����� � �����33� ������ �����?� ��������       � ��������          	!��������   �   �   0   �   �   �   0   �   �   �   0   �   �   �   �   �   ;  �  ��<  � ����� � ���? � ������  ���? �  ���  � ���  � 3����0� ����� � ������ ����? �  ��� �� 3����?�� �33333�� �������� �:    �� �:  ��� �: 8�/�� ��0���� ������ � ��"�(��� ��������          (+  �                                     � <                                     ��  ��� �� ��������� ��3������  �� ���<�0 0��� � � 0 <� 0� �  �� � ��� <�0 0��� <� �0 <� 0� <�  �� � ��� ��0 0��� <�0�0 0� 0� <�0 0�  0 ��� �?0  � � �0 ��  � 0� �0  0�  0 ��� �<0  � � �0 �� � 0� �0  0�  0 ���� ��0  � ���? ��� 0���?  0�  0 ��� ��0  � �� �0  �� 0�� �0  0�  0 ��� ��3  � ���0 ?  <� 0���0  �� � ��� � ?  � ��� �?0 <� 0���  �� 0 ��� < ?  � � ?� <0 <� � ?�   �0 ���? <  � � ?� � �0 � � ?�   ��  ��� �� 0  ��<���������<��  � <                                      �                                                                                                                                                                                                                                                                                                                         ��           �   �  �     �? �?�� <            �   �  �     � �0                   �  �   � � �� <                  �  �     ��� <   ����?��� <<�� �    ��    <<� ��������?� �     ��    ��� ?0����� �     ���   ��� <0� ���� �     <�<�<    ��� �� ���� �     �� ���   ��� �� ����� �     � �0 0  ��� �� �0� �� �     ?� ?�0 0 < ��� �� �0  �� ��    ?� ?���? �� �?��? � �? �?���?��?  ���? �?0�      �  �      0�?                         � �0      0 0                         � �      �                          �? �      ��                                                                                                  %                                      ��                  ��              �                 �?             ��                 < 0             �                    �             �                     �             0    �?0��  �     �0 �  �?  ? 0    ��0�?�?  �?     �0 0  �� �? 0     ��� � �     �� <    ?  0     0 � � 0 �     ��       0 �  0 � � ���     �   ��   0    0 � � ���     �   ��   �    0 � � 0       �  �       �    0 � � � 0     �  �       ��  0 � � � �    < <  �   �    �  <�0 � � �<    �   0   <�    ��  ��0 � �  �    ��  0   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           9       ��                �UU=                \UU�           0    WUUU          0    WUUU      �   0   �UUUU     ��  0   �UUUU     ��  0   ��_�_    ��  0   ��WU�    ���  0   �UuuU]   ���   0   �U�U]  ����   0   �U]�U]  ���  0   �U�U]  ���  0   ����_�   ���  0   �����   ����  0    W�U   ���?  0    _UU�  ������  0    |UU�   0�p��� �    ���  ������? 0      ��� ���? <   �<�< ��0 ���? ������������ ���? ������������� ��� ������>�����  ��� ?�����
�����  ��� ����������   ��?  �����?����?   ��    ����?����   ��     ����?����            ���?���?            ���?���?            ���?���            ���?���            ������            ������            ��  ��            ��   �            �?    �            �?    �            �?    �            �?    �            �/    �            �o   �            �o   �            ��  9             �  9              � @              � @                �                �               l �                l �               �����?              �����              �����?             ������             ������        /                       ��?                _U�              �UUU              pUUU5              pUUU5              \UUU�              \UUU�              \UUU�             �_UUU�            p]UUU�5            p]UUU�5            p]UUU�5            ]�U����         ��_}U}����?�      ��_� W�����       ��W�W����? ��    ���������? ���   ����������� ����   �����_����������  ���_U�����? �����  ����������  ���� ��������   ����  ��� ���   �����  ��� ���   ��j��   ������   ����    ��? ���   ���*    �� ���   ���?    �   ��   ���?    �   ��  ����    �    �  ����   ��    �   ����   �� 0 @�    ���   <� 0 @�    ���   < 0 ��    ���  �  0 �     ��  �  l 0 �       �  <  l 0 �             �0 9              �0 9              �0@              �0@              �����            �����?            0�����3            ������?            ������?          � 0� 0�������zpk��Z���:���Z�@ki��z0����� 0        0 �* � Ⱦ(�#  ��� ��<+ 8��:, 8JU�, 8Z �, � � � � bD � � � �X % �HU! ����. �(0.  �<� 0� � �
 �2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �?��ʫʫʫ���? �                         ��    0    0   ��  �� �?�?���?0 ��?���������������������  ��?0 <��?< �  �? <   < ����?                     �   ��   ��   ��   ��    �?   �?    3    3�    3<    <    �    �?    ��<   �?3  �?3  ��??  ��  0��   �?   ?�  ���  �?�   ?�   �   ��   ��   ��   ��    �?   �?    3    3�    3<    <    �    �?    �    ?   �=   �   �3   ��    ?    30    �    �?    ��    �?    ��   ��?   ��   ��   ��    0�   ��    ��    <�    <�    �?    ��   <��   ���   ���  ���  ��   �  ���  ��   ���  �?�  ��    �?    ��   ��?   ��   ��   ��    0�   ��    ��    <�    <�    �?    ��    ��   ���   �|�   ���   ���    �    ��    �    0�    �    �                                                         ��    �           30  �30� ���� �������?��?  �? ��?�� �?003 �?��    ��                           ��    0    0   ��  ��  ?  ��  0  ?����������?�����?������ ��?�� ��?��  <    <   ??   ��    ��   ��?   ��    ��    �?    �?    �?    ��   �<   30�   33�   ��   �?�   ��   �?�   ?�?  ���?  �?�  �?�  �?�  �       ��   003   ��    ��   �?  �  �  � ���  0 �� ��� ��� ���  0  � �� �?�������� �� � ��� � �? ���   �?�?  �?�?  �?�  �       ��  003   ��    �                         ��   00 �00 ��0����0?��0��������0 � ���� ���� ����  ����  ��?0 <��?< �  �? <   < ����?                   \�ʁ8����6�������    ��� pUU��7����p��p��?��wT�����[��W���UU����:��>����� pUU\UU5\U�WU�WsU�SsU�S}U�SUU��U�\UU�\UU����� x�  x�  ��    ��� pUU\UU5\U�WU�WsU�S}U�SUU��_U� pU��U�\UU�����W\5��?���UU\UU5WU�5�U�՛U�՛U��kU}�kUUśU���UU5WUU5���? W-  W-  �/      ���UU\UU5WU�5�U�՛U�՛U}�kUU�kU���U �U�?WUU5����\5p��?�����pUU\UU5\�5W��[s��[3��[=|�WT�����[UU�WUU�����\5\5\5\5�?�? � ��: ��� ��� ��� ��� ��� ���  ?� ��<0<00��?�             � ��: ��� ��� ��� ��� ��� ���  ��  ��  ?<  �? ���0����     �����=��5��
���*���+���/���3����?�� �� ��   �  ��  �� �p=���5�����
���*���/���3����?�� �� ����?��  �    ��? |��\��נ�?ר�?��??��?�������� � �� �� ��  0  ���� |� \��W��נ�?ר�?��??��?����� �� ������0���0�?���� �   03  �� �UWpU���5���7��7\��5\�_5\?�5_��s���UU�?���         �   � �W �\5��\5��W���U��:W��:W��W���U��U� �� ��  ��  �� 0 ��  p� \5? \5�_կ_U�:_լ�_լ�_���sUsU����  �?  � ��?         �   ��   ��   ��   ��  ���  ���  ��;  ̣�3  ��  0�  +����ꫪ������W�:���W����W��~�\��W�\���W5p���W�?  �                                  ��   ���   ��:  ���  ���  �� ���  �>�� ��>�� ��>��  ����  ����  ���� ���������������:��꿪���zժ���_U��  WU   ��     ��   ���   ��:  ���  ���  �� ���  �«� ��«� ��ʫ�  ����  ��  ��� � �������������:��z�����z��������  p�    pU   \�    \    �                    �    ��   ��>   ���  ���>  ����   �*�  �*��  �*�. ���� ����  ����  ���� ����������������������W����U�� pU�   ���  �    ��   ��>   ���  ���>  ����   �*�  ���  ��. �꣮ ����  ����  ��>� ��� �������ꯪ��z����~����W��  W   �U    _5    p5    �?  ���������`����&�܅�.�p�����h�6�6�x�x���G����Ӫ_�%�뭱���� �U*
Z��*���*�z����ﯰ� �?  Ҍw�!��%�K���C�I�[�  ��?���<��?    ���0 << � � � � �< 0� ?��      ��  ��?   ��  �   <   <<   0   �   �   �   �   �   �<   00   <�   � � ? �  ��?         ��   ���  �  <    ��   �    0    <<    0<    �    �    �    �    �    �    �<    00    <�    �    �  � ?  �  ��?   �� <��<  ��?���������?    �����?�����������������?��?�� �?  ���WU�UU=|�5\U_�\U_�\U_�\U_�\u_�|�_�|�W=�UU�_� ��      �?  ���WU�UU=|��5\ue�\ue�\ue�\ue�\ue�|�e�|�_=�UU�_� ��  �?  ���WU�UU=|�w5\uu�\}u�\]U�\]U�\]}�|u}�|�=�UU�_� ��      �?  ���WU�UU=|�U5\uU�\uU�\uU�\uU�\uu�|uu�|�=�UU�_� ��      �?  ���WU�UU=|�5\uu�\uu�\uW�\uW�\uu�|uu�|�=�UU�_� ��      �?  ���WU�UU=|�_5\uu�\uu�\uu�\u]�\u]�|u��|�u=�UU�_� ��     ��Î�C���Ǐ ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              1d h h � � � � � � *5AUUUUh�����'B[w�������������4Pl�d ��?�wU�uU�uU�uU�uU�uUUuUU5��U��U��U��U��U��UUuUU5��WUU�WUU�WUU�WUU�WUU�WUuUU5�W}U�U}U�U}U�U}U�U}U�U}UuUU5�W��_U��_U��_U��_U��_U���UU5�WU��UU5���U�_U7�w]�WU�]�5W�UWU���5��UU]U�u]�7��UU]U�WU7�wUUuU��UU5�wUUuU��UU_U��UU5�wUUuU�}UUU�uUU5�wUUuUU��U�UU�UU�}UU_U�uUU5��UU]UU_�W__U__U_UU_U�uUU5��UU]U�W�Uu�Uu�U}UU_U�uUU5�W_UWU�W�U��U��U}UU_U��UU5�W]�UU�W�U��U��U}UU_U��UU5���U�W_�U��U��U}UU_U�_U7�w]�WU�_W�Uu�Uu�U}U�]�5W�UWUu�U�W}�W}�W}UU_U��5��UU]UuUU�W]�W]�WUUU�5��UU]U��U�_U�_U��WUU���5�wUUuUu��U�u]�7�wUUuUuU�U�WU7�wUUuU�UuU��UU5�wUUuU��U��UU5�wUUuU�uUU5��UU]U�uUU5�W_UWU�uUU5�W]�U�uUU5���U��UU5�w]�WU��UU5W�UW_��U_��U_��U���_���_UU7��UU]�WU_�WU_�WU_u}U�u}U�U�5��UU]uUUuuUUuuUUuUWUUWWUU_�7�wUUu]UU�]UU�]UU��U��U��W5�wUUuWU�WU�WU�wU�uU�uU5�wUUuWU�WU�WU�wU�uU�]U5UuUW�WU]U�]U�_�UuU_�Uu�U_UW_�]U��U�]U��WU�WU%�8AJUamx���������2Ol����.Qv���2Lf�����7Tm�����4Sp���� A`����Aa���	)	J	l	�	�	�	�	
=
b
�
�
�
�
@d����.Op����0Nk�����*Ig����/Sw����+AYgu}�������� � � �2Lh����\	U�� �\	U��
 �\���ת �\uU�uժ �\U��ת
 �\WU�ת* �\WU�ת� �\WU�ת� �\WUU��U�ת� �\WU�U�WUUת� �\WUu_UU]UUת� �\WU�U�uUUת� �\WU�U��UUת� �\WU�U��UUת� �\WUwU�WUת� �\WUwW�UUWUת� �� �\WUwW��UWUת� ��� �\WUw�UUWUת� �� ���� �\WUwuU�UWUת� �|= ����? �\WUw_U�WUת� ��\5 ���� �\WU�PU�WUת� ��WW5 ����� �\WUUuUUWUת� ��UW� ����� �\W�PU}UUWUת� ���U� �����? �\WT��_UWUת� ����? ���� �\WU���UUת� ���}� ���� �\WSU��U�UUת� ����_U  ���� �\WC��UU}UUת�  ��U  �? ��� �\W]�U_U_UUת� ��p�U  �?  ��� �\W�WWU�WUUת��� p��  �� ���� �\WUU��U�ת��  �U� ��? �?�? �\WU�ת� ��� 0�
 ������� �\WU�ת� �0�. ���� �\WU�ת� ���+ ���� �\WU�ת� ���� ��UU��? �\WU�ת� ���� �UU��� �\U��ת� ����  _U��� �\uU�uժ� ������W�U��? �\���ת� �����5\W��? �\	U�ժ� �����\\��? �\	U�ժ� ����
�\\�� ����/  ����=\=\u� � ���_
U��  ��+��\�\u�  ����_
U���  ��* �_�_U�  ����_���w��
 ��* �W�WU�  �\uU�W��
 뿫 ?T�UU�  �\U���
 ����CU�u5  �\WU�u��
 ���>TU]U�?  ����^WU�u��
 ���OU�UU  ��  \WU�u��
 ���CU��WU-  ��
 �\WU�u��
 ���U���U�  �� �\WU�u��
 ���@U���ϯ�*  �� �\WU�u��
 ���P���>���� �" �\WU�u��
 ���W����������  " �\WU�u�� �?����������  " �\W��U���Uu�:0 ����� � ������� �  �\W��WUUu�Wu�� ���?  <0������� �  �\W��_UU��_u�� �  ?����� "" �\���UU��u��0����?����� " �\���UU��u��3����?�?����� " �\���UU��u�3<������?���� �� �\� pUU�|u�00����?�� ��? �\70 pU� ��u������?�����;� ��� �\�pU���w� ���?��?��?���;�  �  ����\U����w�  ���? ?��?����  �?  ����WUU��\u� � ����<��?����   � \� _U�=|_u�?  �� �3��?����   � \��U��_Uu��  �? <������� � ���\WU�u��
  � ?���?��� � �0�\WU�u��
 �?������ � � � ��@U�u��
 �?������ � ��?  <� �@U�u��
 ��?������ � �� ���W��  UUu��
 ��?��? � ��  �3P�_��U  T��
 ��? ����� � �� ��@���U�WU����
 ��? �����  ���?���_U�W����
 ��� ��  �� ��_U�W��U��
 ��0���?��  �  � �_�WU�U�U�? 
 �� ���?��  �� � �_�W�_U�WUU?< �� �����  �� �_��_UU�U�?� �� ������?  �� ����U��UU�?� ��������?  �� �����_�U�� ? ������sU�  �� ���U�����W � �����sU� � ��*�? ���U����U �? �� ��_U� ���������W����@��� �� ��\U5 �\U�����W��UU ��� ��?��?WU� �\U�����_��U���?  �����?WU�� �\����������?T��?�?   �? �?WU�� �\uU���W���?  �?�?    �? �WU�� �\U��W�����  �?�  < �? �\U��� �\WU�U�����  � �  � �? �\U����\WU�@������� �  � �3 ����?�\WU�P�����?�� �  �  0�  �
���?�\WU����U���� �  �?  0 3 �
����\WU���U��� �  ��   3 �
����\WU��  ��� �  ��   3 ������\WU�յ������� ��  < ������\WU�յ������ � �   < � 0����\WU�յ�� ��<  � �   0 * 0����\WU�յ��  ��  0����   * 0����\WU�յ�� ��? 0�� �  �
 0���\WU�յ�� �����?? 0  �
 �?�\WU�յ�� �����?<0  � �<�\WU�յ�� ����?030  � � <�\WU�յ�� ��� �0  � � � <�\WU�յ�� ��� �3 � � � �<�\WU�յ�� �� �3 � � 0 �<�\WU�յ�� �? ?� � �  �<�\WU�յ�� �<�� � �  ��\WU�յ�� ���<� � ��\WU�յ�� ���<�� ��\WU�յ�� ���<< �� �\WU�յ�� ���0<0 �
  �\WU�յ��	 �<�� <�*  �\WU�յ�� ��� ��  � � 0 �\WU�յ�� � ��  �� � �\WU�յ�� � ��   �  �\WU�յ�� �� ��   �
  �\WU��WU��Wյ��	 � �    *  �\W��?\U�_յ�� �0 *  <    * 0 �\Wu�?p��pյ�� ����    0 � 0 �\W���su�pյ�� � �   0 � 0 �\W��0|u��pյ�� � ��   � �0 �\W��pu?0sյ�� �� �� � � �0 �\= p���p���� �  < �0 � �
0 �\u p5 p]��* �� � �0  �
0 �\� 0p �ߵ� ��? ��  �
 �\U 0p 0U�* ��� �
 �\U 0 �U� ���� ��33�������? ����� ��  ����� ����?��  ��� �� ���������  ����� ���  ����?����  ���  ���  ��  �� �����<��� �<<�<<< �<<< < <<<< ��<� � �<<�< � �?���?<<< � <�??<< � <��<�<�  ��������?�? ��?�� ?����	  ������ � ��� ����	  ������ �� �� ����	  �������   � ���� 	  �� ���  < < �< ����	  �� ��� � ��� ����	  �� �����?�? ��? ����	 	  �� �����?�	  �� �����?�? �? ���� �?  �� ��*p�N\�R5WT������R�:�R�:�J��J��J�  +:  ,  0  �     �    ?   �  ��_  �u�  ?pU5  �_U5  pUU  p�_�  _|U��?pU���?pU�W?\��W��? �WuU5 pU��� �_�j�  \���  WuU�  ��?   ��    ��  ���  ���  �   � �   p�   ��s   W]   \U�  \U�7  pUU  _� �U=�� _U�WpU�W�W5��: ���� \U]�; ��WU W�W� ��W5  WU]�  ����   �>   ���   ���  ���         �  �  � ����?���������������������?������?�����������?���?� �� ?���  � ��  < � < ����0���3 0 �   <  00�0�0�  �  0����00 < = �� �� p�pY�\U��0 0ww= 33ww��033�� ��?        �  �  � ����?���������������������?������?����?���>�����?� � ?���  � ��  < � < ����0���3 0 �   <  0�0��3�0 p} <��\I=?�_I����_Iͯ��pIëꬪI��:��sI�����հ��� ?��          ? �  �� �  ����� <���W�<�lU}U9���U��������������W��W{U}U��[}U}��[�U���Wk�U���_�U}U����U�U�?��V}�� �V}�>  �V}�>  �V}�>  �Z}�  �Z}�  �j}�  �k}�  ��}�   �}�    ��?    ��    ��           ? �  �� �  ����� <���W�<�lU}U9���U��������������W��W{}}}��[�U���[}U}��W[UUU��_k�}W����U�U�?��U}U� �W}�?  �}�?  ����?  ����  �U�  �U*  ��V�  ��Z�   ?j�    ��5    ��    ��  ��   ����?�����?<�?0�<�����?��WUU�?��UUU���U}� \W��  \���  W��?� ������?�_�����_�_?�UU�UU���_��?�W�_�;��� ���z����zU�U���UuU�:�_u���������?�ꪪ�� �ꫪ����������3<         ��   ����?�����?<�?0�<�����?��WUU�?��UUU���U}� \�W��  \��<�  W� � �����?�_�����_�_?�UU�UU���_��?�W�_�;��?���z=s���z5 p���5�\�:�7�ת�������?��^U�� ���U������������  ?�         ?     �� �� �,_U��8��UUU:�
_U����zU�� �_U��  \�UW5  W�UW� ��uU]W��_U�_��Up ��� � �� p���\ � �5\��U5\���W5pUU�UU�U��_U W�U��  \_}�5 �sU�U�p�� Ws\5? �\5\5   \5�?   �?       ?     �� �� �,_U��8��UUU:�
_U����zU�� �_U��  \�UW5  W�UW� ��uU]W��_U�_���U�s  � � � � �p � �p � �p��Up���WsUU�WU��U� WU�7W5 W���\5 W5�Ws5�U��W��pUs���\���  \_    ��  UU0      0   �  0 �  0   8� 0� 8 (0  �.?   0?��   ���  ��56�   �D�   ��3  �����        �/Y�  �-�  0.;?  �*<  �� ���3 �  �� �  0 0�  0   �  0   �  3    0 3  0       �  3   �0 �  _3 0  0W��  ��s�  ��s�08 �
3*4 ��� �gP�� pG@���?  ��0       ?W@���� �� /% �� � u� ?CQ���@��  0T�?0 ���00 �p1?� �0��0 3 0 3 �0   0  		

���k����#�;�K�o���ó��K�{�˴۴�G���õ?���϶߶�_�����#�3�w�����������Ѹݸ����.�F�X�p�y�������ʹ�����3�K�c�{�������D`x D`08xxxHHHH`HHH@HxHxx8`H8H(HXHPHxH`xHxHxHxHHxxxHx    �� x �x�    �� HxH(X
   � �0H`x (0(08@8@HPHPX`X`h   � � xHxpx   � �0H`x���0�H�`�x ((80PHxX`hHx0    ��P0P8�8@H	hPP`Ph�hPxh� x0`  	p 	 H X�X �   � �8 X (0h0 ` pHp�p �  `  x H`H P�P �`�@((h
0 h  `p` h�hxH� �  � (�(@h@8`8h`h�`�  �  �  � �  (p(00`0HX8`X`(hhh pxp  �  �    � �0hp(P8pXPpp�P   � �(X(@0X0@X@X�XXpX(`p`p`p���   � �  � H�888X8x8X(XhX�Xx8xXxxx  � �0`0 Pp`p �   � �0((8 HX h(x0�8�(�8xHpXhh`xX�PH@   � �0h�(�
8xHp   � �0H`x��0�H�`�x �  ((0088@@HXH`@h8p0x(@h8p`p0xhx   � �0H`xpp0pHp`px0h8PX0Xp   � �0H`p0pHp`00h088XX �8�Hx   � �   � �0H`x�p0pHp`�x0h   � �(@Xpp(p@pXpp0(
h(
���   � �H@X@(8h8`xP  �   ((0088@`@h8p0x(� ��� �(�0x8p@hXh`phxp�x���H`   � �   � �   � �  	X 	 `  x  0�0 @�@ `�` pxp �`� �0(�0h�0@�0P�0(H0BH0VH0hHp�8(�XH�0�X���h8�XP�8Hh�hp8X8XPpPphXhX�p�P808`8@8||     08p0p0�p0Xp0`80(80`X0(X0`x0(x0 h0h0�h0ph08�0�0��0X�0�00(00h00xp0p0�00p0 0(X0hX0`0x`P PPXP8P�Pp000�0`0`�`�xx||     #0(0X(08(0x(0� 0 00 0` 00`0``0p�0 � x88hXXXx xHhp(p���PHPP��h ( (hh�hhh0� 0 0�8080�P0P0�h0hP�P0�8080�P0P���||     (�8p8�hhPXP88P�P�00 HpH�``P�PH88h(((0��0�P� P P�HPH���0h 0( ||     -||     2||     7|P|�P|`|x`|(p|hp                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���آ t ���d���� � �����������  ��� � �� � �� �ύ& ��"  7ĩ�� d
�� ��L`�       ^�n�~�������������������.�>�N�^�n�~®¾�����������.�>�N�^�n�~ÎÞ�                                                                                                                                                                                    �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  HZ�H�@��m��������8��HJJH

�zh8����m�� ����ɪ�8��i0��i ����h�zh`H�i0��i ��_�����8������h`H�H�H�H�H������ k�h�h�h�h�h`�H�Z�ڮڦڦ� ��8��JJ�8���� � ����� ����h�h�h�h�z�h(`Hڭ  �� �������%���h`����������ow{}~���������������������H�  ����h`�H�Z�ڦڦڦڦ�
��`���`�� �â �  q�- �� q�- ��� Ā��iɠ���iɠ������h�h�h�h�h�z�h(`Hڪ)�JJJJ Ŋ) ��h`HZ� ��$�#�0i��:8�0��A08�7�i �Ȁ�zh`�H����� L��Z�H�H�H�H�H�H�H��H��Hi�H�i �H ��8��JJ�8�����m��i ��������?������6� ��ȭ��h�h�� �������� ��m��i ���hh� h�h��0�� �����������ݬ�������
�h���h�	��h�h�h�h�h�h�h�zh(`�� �2��.HZ�Z�Z� ���������
������� �h�h�zh`�H�Z�H�H�H�H�H�H �à �ȍ���-�i��i �� � y�����m��i � ����h�h�h�h�h�h�z�h(`� �#��H���hH�Z�ڦڠ �������Lv�L�L~���� �Ȁ����LYȥH�H�Z�
�������������	8������	�� ��������*�e��i ��e��	i �	� �������	���8����	��������
�8����������������8h���h������
�������	��������h�h�z�h`ڦ
����	��.������`H�� �� h`�  � `H�Z�H�H� H�H�H�H�H�H�H�H�H �Ì�JJ�NN� ����:����:�ȱ���:����:��8�����h�Hڭɀ�
��8�
���Hȱ�����he��e������� ��h�+� � � qʍ �� �3� m������ q�ڮ� y�����
������P��r� m�����m ����8� � �8� �	� �m ��H q� y�h��,���� qʍ �� �� � q�ڢ ��� �� ������ �L.�h�h�h�h�h�h�h�h�h� h�h�(z�h`Z���z�`Hڦ��	���Q����h`�ڮڮڍZ�)���=%ˑȱ�=(ˑ8����Z�JJ�����

������	��
�M��z�

�����JJ����z��ȭ�h�h�h��h`?���H�Z�H�H�H�F�H� �

�ȱ�z��Z�H��hHڍ ǭm����m����hhh�h�h�h�z�h`��d % 4 O B 
 z  0 
7 p 
   � � ���7�kĺ���ŀŕ������vǀȗȦȭ�q�y�,�                                                                                                                          x�d�# X � ���t���H���:�;�<�x����X � �� � 2� r� {� �Э= ��B�&�6�!�
����
�
�
�� �ꀜ ��í)|�|� G� �� �ϥ�
�	��
������
�
 �ĭ�
��d�5��
��L��0ͅ�1ͅ   �ϥ���L��N������9�:�;�;�c�X�H�  ����h`�H�H�H�	H����  �8��i�i�� ��ک �	������ � D� �֭  ��� Dͩ �	h �� v������  �h�	h�h� ��dh(``H�Z�  �խ�� �� �Ԁ 7� 7լ5���>��1 *� �� o�ڥ�� �� � e� � W� b� W� �� �d�耫����� ��z�h`H�Z�H��	H�Z�H���5� ;�����5 �Վ �բ �0� �խ�� �Ԁ� 7խ5���Q���I��ܭ5��� K���A *� �� o� o�ڥ�� �� � e� � W� b� W� �� �d�耐�5�����	���5�� �՜5h�z�h`H�@�� �ե@�A��@ �� g�h```H �� Kԭ���@4�@�������@4�@�� ���@ �ե@�Ah`H����5 �� 7խ5�������5����A�@ �� ��h` H�  �� Nͩ,4���� �� � e� � �� �d �֥�Ȑ ���� vϥ��8 �� � e� � W� b� W� �� �d�$����$��#����#d$� ��h`��C���D��E ��#�%��H�
H��
 {�h�h`H P �H �H(`H �H hH �H �� �H � H PH � H � � H � H h8 �8 �H @ H � H Px � H �� � H � H hX �X �HP� H �Hڢ	�
�Z�����t&���I�

��dЅ&�eЅ'�fЅ(�)�gЅ*��Ѕ+��Ѕ,��Ѕ-�.��Ѕ/��Ѕ0��Ѕ1��Ѕ2�3��Ѕ4 W��h`H W� ҥ��d �� W�h`H�Z�H�H��H��	�҅�������

m���&��'��(� ǈ�h��h�h�z�h`H�Z��H����

m���&�@��0� ���(�(�*�,�&�(�(::�(�)��&��'�'�*��&��'::�'�)��&��h��z�h`H�Z��H����

m���&�d�i��'�X8���'�O�i�(�E8���(�<���5���4 �յ&H�'H�(H��'��( �ѵ'��(�h�(h�'h�& �Հ��h��z�h`H�  ��Lm̩�������������h@H�Z�' )������ � 	�P�# �$ �% (z�hX@H�Z�H�H�	H�H�H�H�H�
�簍��
��'�� �(��!������� �	 iӢ �

�� �ȱ �ȱ �ȱ � ,� ������h�h�h�h�h�	h�h�z�h`ڢ?�=����`HڭmJJJ���m�������mJJJHJJJHm���h


��8h����h`H�Z�H�H t�hH�������>�>��
���� Ȁ�����i����h�h�z�h` @��Z tӬ�����9>z�Hh`H��HJJJ


��hH8�����hH8���h��h`HڭH�Hi�� "ԭ��>��� "ԭ�����hH�hH �ԍ������ ���i������h �Ԁh �Ԁh�h��h`8�`i`8�`i`H�Z�H�H��M�� "ԭ��9�8����� "ԭ�������i� �����i���h8���h�h�z�h`H�Z�H��H� �� @� �խ5���K��|�H�� "ԭ��@�i��i�� "ԭ�������� �����i���hh�h�hi�h�z�h`Hڭ	H�i��i� �Ŏ�� �Hڭ	H��	�@
��ȅ��Ʌ� �h�	�h`H�	H� �	�� �� v�h�	h`H�Z�	H��H ��d��@�

������� �� ��i٨��� �� �� �ր� �բ�@ �� �� �� �� �� �� ���	�� �բ�@ ��h��h�	z�h`H�Z �� � � o� o� o� �� � ��z�h`H�Hd����h�h`HڭH�H������� �����H���H� hJH,��9׀�$ �����h����= �ũ������	�cׅ�dׅ ǩ�	h�h��h`   �? � � 3033��?� �? ?�@�Hک,4��,4� ��Ld� �ۭ  )� ��Ldة,4�
����
��ɠ�(�)?����0�����"�Hmɓ�h�@-4�4�Ld�h���������� �0�

���}�}d�] p���V�  )��8-4JJJ���܍�4�� #܀1�8-4JJJ���


H��-4�4h4�4��܍�)�	��h`Hک,4�A�,4�@ ݭ�������� p���!�8-4JJJ���܍�4�� #܀ �� ��h`H����  �@-4�4JJJJJJ	4�4����܍�i��8�
�h`H�Z� �

���L�٩�<���ɠ�0����)?�����:����H}ɓ�h�L��h���������� �L�� �ٽ����h��'���$��%�H::�h�&��'�=�� ����  ���� ���� �ڜ���'�'�"�"�+�+���L��z�h`H�

��`=}�`�d�P ��އ�!�"�}��B�P �۩�6�ڽ�7���8�h`�H�HdB�}����  �~���� �	�w���� � �֩���  � �� �֩!���� � �֩���  � �� ������ � �֩���  � �� ������ � �� �֩���  � �� �� ��h�h��h`Zڮ��H��

��������Ρ��hH����hh���z`�Z��H� � �

�hH���}�D�~8��� ͢�4�})}~͢�&�8�ͣ��})}ͣ��
����  ��̟����zz�Hh`��m�8���Li��D��8��Ȱ��5��m����'����4��4�8������  ��� `H���m�� }�� ����(�h`H����)
�����m����m�� m�� m���(�h`Hک,4����J���L��H�� ���� ���� ���� �ڢ �������$��!h��)8���8�����i��"i�"�5��!���i�i�i�#�i�i�"�h``         2 dH�Z�H�H�,4�/��z� ��������
������������� ǀP��

���*ڢ ��������
������������ ǈʠ �

�������@-4�4h�h�z�h`H�Z�H�H��	� �

��}�B)H�~���hHm�hm�� �Ŋ�ڝ��})`JJJJ���������� ���̟����	h�h�z�h`H�Z�H�H� �	����

����H�~JJ

���h �� vǞ��٩�	h�h�z�h`H�Z �ե%� � ޭ
��U� �

��}�D�})`�`�2��<}�����,�=}�}�"ڊJJ����� I� � b߀	��� ���̟�� �ݥ%� � ��z�h`H�����4�R�~�~�~�>��|�d��]��Y�~�~�~���@�K��D��@���� �6�~�>��@�+� �$�� ����t��~���|�� ��� ��h`H�H�H�})`�@�X��� "ԭ��9�~�� "ԭ���})}�ڭ����� ���i������ɘ�� ��� J�h�h�h`H�Z�})`�`������K����E��<}��
�:ڊJJ�����ڊJJ�����"��,��,����� �,������ ��ȱ�� �z�h`H��� "ԭ���~�� "ԭ��e��,���})}~��~8�� ��\�i� ��6�`=}�Y�8�� ��@��,���~i��~8��~���5��,���~�~�%�~�~��`=}��8�0� �ڊJJ�t�h`H��,�����h`H��,�����h`H�,4�G�,4�@�8���4�i��)���!�i�� ݭ��)�	� �h`H�Z�(���d#d$d% 7� �� �Ү
���B
eB���
��g���h��� � ��}���}���}��}�̟�✞�����
H8��h����JJJ�


͟��B�B�:

���B�� �� �z�h`HڭH�H�6�i�8�8�8��Yڢ�8����8����7����� p������6����6�#��8JJJ


�8��6�6��
��6��6h�h�h�`HڭH�H�6� 
��������7��8���	 �h�h��h`H��|��#h`H�i�������� �05�
��0�=� �թ�@ڢ �� �� �� �� �������=0 �h`

��}��� ���B��B����=��H�Z�~������̟�W�

��}��~8�	0͢��i͢�ܽ8�	0ͣ��iͣ�ǜ���,���zZ��,�����
�����8z�h`H�}H�~H�H � L�C�}�D�~�E��i�������� �0d#d$d%h�h�~h�}�L�� �h�h�~h�}h`H�H�H��	�#�����D��E� �h�h�h`H�D���8��i�D�E���8��i�Eh`PASSWORD$PRESS  START$LEVEL  $GAME  OVER$TOP  SCORE$YOUR SCORE$��u�~����H� �	� ��������� � o�r�����d���� � ;� o�������� � ;� o� 7ĩ��T� � ;婀��  �d o�:��h`�H�H�H�H��������� �h�h�h�h�`Hک �2:������h`ڮH���H�9J
�9�����Hi���H�`8�H���H)�H����Hi��H8�)�HhH�˩�x�����P�9�i���� �à ����?ȑ(`� ��H�  �h`H� �h`H� �h`H�
������� ���h`H�Z 7ĩ���� � ��������� �ȩ �9�P���� � �� �� �ĭ� �E����
����&�ѭ9J��: ~�:����  ����9�� ��9��9��� ��9�ۢ������

m
����:����;����<���ۘ

�
��=����  �z�h`      I C $hvI�5CHڢ �: �������h`Hک��& �
JJJ
�� ��������� ǭ���	����n� ǩύ& �h`H� 7� /�H��� 橀��
�
�i��
i�*�i �ŭ
HJJ

�
�8JJ�

m
�h�
��:��;��<���F� �`� �h� ��Z� � �ĭ� ���h`H��� � 7� G詏�& ���<��
����� ǩ� o�:���ύ& � �� �h`Hڜ���� �X��� ��������� � ;�X��� �����h`H�Z��� � 7� G��������� � ����� �Ȝ�_���@ �� �� �խ  ��P��D�ɠ�E��@��֩�Ԣ�@ �� �� �� �� �� ���	���@ �� �� �� �� �� �խ�� Dͩ���  � �� �z�h`H���>��"���2�����&��
������������h`�������������������������������������������������������������������������������������������������������������������� �
���� ��������������������������������� �����
� ������� ���*��������������������������� �������������������������������������������������������������������������������������������������������������������Hک�� � 7� G詯�& � s� �� o� o� o� o� �� b� o� o� o� o� b�:� s� �� �� o� o� o� o� �� b� o� o� o� o� b�:� �� s� �� o� o� o� o� �� b� o� o� o� o� b�:٩ύ& �h`H�H�H��	�(��$������� �h�h�h`H�H�H��	�(��.������� �h�h�h`H�H�H��	���������)� ǩF� ǩ|� ǩ)� ǩ��� ǩ4� ǩX� ǩ|� ǩd��� ǩ4� ǩX� ǩ|� �h�h�h`H�H�H��	���������%� ǩB� ǩx� ǩ%� ǩ��� ǩ0� ǩT� ǩx� ǩ`��� ǩ0� ǩT� ǩx� �h�h�h` �v���3�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     L�L��L]�LF�L� �P�Q�R �� �� � � � � � � � �* d�d�� ����d�`�Q����y� ��r� �s�  A��y�y�t� O�R������ ��� ���  ��憥�Ł� ��P���J�Q����]� ��V� �W�  ��R����k� ��d� �e�  ���]�]�X� ���k�k�f� 
���� �� ]�`�S�T�VȱT�WȱT�XȱT�YȱT�Z)
�����[轑��\�Z)0�`ȱT�����ȄSd]d^�X� �L��_ i�� �
�T� �d_��Ȅ_dS���o�p�rȱp�sȱp�tȱp�uȱp�v)
�����w轑��x�v)0�{ȱp�����Ȅodydz�t� �� �Q� ��)��	���Rd| ��`�|�}�ȱ}��ȱ}��ȱ}��ȱ}��)
������轑�����)0��ȱ}�����Ȅ|d�d���� к� �R� ��)��@Ы���Qdo O񀠤a�b�dȱb�eȱb�fȱb�gȱb�h)
�����i轑��j�h)0�nȱb�����Ȅadkdl�f� й�m ��� �
�b� �dm��Ȅmda����
��=����=������Tȱ��U`��
��C����C������bȱ��c`H�Z�Y)?	@���Y;��%����^�[��Z)@��J������`�8��`��Z)0�`Ȅ^�[����^�Zd^��� z�h`H�Z�g)?	@���g;��%����l�i��h)@��J������n�8��n��h)0�nȄl�i����l�hdl��� z�h`H�Z�u)?	@���u;��%����z�w��v)@��J������{�8��{��v)0�{Ȅz�w����z�vdz��� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ƈ��d���� z�h`� `� `H�Z���������������)?
������轥���d� "�z�h`d��* d�`������ȱ���ȱ���ȱ���)
������轑�����)0��Ȅ�d�d���� �d�`H�Z�����L��������;��)����������)@��J��������8������)0��Ȅ������Ɛ��d���)����)����
�@����������( ��ŕ��* ��捥�Ō� "�z�h`H�Z�  i�  ��dSda��_�m �� 
� �� �� ����Pz�h`H�Z�Q� ��R� �d���)?Ŝ�D�� �>��
�����p����}轁��q����~dod|� �Q�R��)�����R �����Q O� ��z�h` �(�� ��� ��� �(�� ��� ��� �(�� ��� ��� (�� (�� q(�� P�� �(�� (�� �P�� �(�� �(�� �(�� ��� ��� �(�� (�� (�� �P�� �(�� �(�� ��� ��� �(�� (�� (�� �P��     � �
� �
~� �
}� �
|� �
{� �
z� �
y� �
x� �
w� �
v� �
u� �
t� �
s� �
r� �
q� �
q� �
� �
~� �
}� �
|� �
{� �
z� �
y� �
x� �
w� �
v� �
u� �
t� �
s� �
r� �
q� �
q�     � �
� �
� �
~� �
~� �
}� �
}� �
|� �
|� �
{� �
{� �
z� �
z� 
y� �
y� 
x� �
x� q
w� 
w� q
v� 
v� d
u� q
u� d
t� q
t� _
s� d
s� _
r� d
r� K
q� T
q� K
q� T
q�     � q�� <�� �(�� (�� �� �<�� �(�� (�� K�� ��� ��� ��� T�� ��� ��� ��� ?�� ��� ��� ��� K�� ��� ��� ��� _�� ��� ��� ��� �� ��� ��� ���     ��(� ������}(�}��}��.(�.��.�� �(�  (�� �(� �P� .(� �(��P� T(�(��.(�.��T��}(�  (�� �(�.P� T(��(���� ����(�� (� �(��P�      ��
�
��
~��
~��
}��
}��
|��
|��
{ �
{��
z��
z��
y��
y�}
x��
x��
w}
w��
w�}
v��
v�}
u��
u�}
t��
t }
s��
s�}
r��
r�}
r��
q�}
q�     �T
}
�T
~�}
~�T
}�}
}�T
|�}
|�T
{ }
{�T
z�}
z�T
y�}
y�T
x�}
x�T
w}
w�T
v�}
v�T
u�}
u�T
t�}
t�T
s }
s�T
r�}
r�T
q�}
q�T
q�}
q�     � �� �<��.(�  (�� ��<��T(�  (�� ��T��.��T�� �� T��.��T�� �}��T��}�� �� T��h��T����T��@��T�� �� T��@��T��     �.���� �(�� (�� ��� ��� �(�� (�� �� q�� d�� _��     � K
� K
� K
~� K
~� K
}� K
}� K
|� �
|� K
{� K
{� K
z� K
z� K
y� K
y� K
x� K
x� K
w� K
w� K
v� K
v� K
v� K
u� K
u� K
u� K
t� K
t� K
t� K
s� K
s� K
s� K
r� K
r� K
r� K
r� K
q� K
q� K
q� K
q� K
q� K
q�     � ��� ��� ��� �� _�� K��     � �
�� /d��     ���_�����_��     � �� d�� T�� C�� ;�� 2��     �     �
�

		�
	 �
�



	�
	

			 �
	
	 �
	� �
	�I�q�}�]�w��x�D�D�
���
���x�D�  ��b�b�(���(�����D�  ���  ���      "���4�R�"�|�|�|���������������*�2����������� % O  % O     % o  %                                                                                                                                                                                                                                                                                                    �� ���