��� � �[ �  ���D�P��  �ݩ �t  �ݩ��t �[  ��� �[ ���� ��˩�� �ĩ�� � �[ �  ���m�P��  �ݩ �t  �ݩ��t �[  ��� �[ ���� ��˩�� �ĩ��M  ���a �`�b �
�� ��� �*�� ����  �ܩ!�� � �[ �  ���h�P��  �ݩ �t  �ݩ��t �[  ��� �[ ���� �"�˩�� �� ���a �8�b �	�� � �� �+�� ����  �ܩ"�� � �[ �  ���h�P��  �ݩ �t  �ݩ��t �[  ��� �[ ���� �&�˩"�� �� ���a �U�b �	�� �!�� �,�� ����  �ܩ'�� � �[ �  ���3�P��  �ݩ �t  �ݩ��t �[  ��� �[ ���� �*�˩&�� �ĀP ���a �=�b �
�� � �� �-�� ����  �ܩ���  �� �ݩ�� ��� �	�a ���b �.�� ����  �ܜ� �  ���L7� ��  ��� ������V���U�:�jU�:�ZU��Ze��V�U�V�U�VUU��VUU��VUU��V�U��V�U>�Z��?������ ���  ��  ��  ��� ����𫪪����:�VU�:�UU��UU��UUU�j�U�j�V�j�U�UUU�UU��UU�:�VU�:𫪪���� ���  ��  ��  ��� �������Vj�?�Uj�>�Uj���UU���UU���UU���Uj��Uj��VY��VU��ZU�:�jU�:�������� ���  ��  ��  ��� ����������U�?�ZUU>�VUU��UUU�kUZ��k�Z��kUZ���UUU��VUU��ZUU���U�>����?�������� ���  ��  ��  ��� �����ZU��VU�:�UUU:��U�ꫪU�ꫪU�ꫪU�ꯪU����U����U����U����U�>����?������ ���  ��  ��  ��� ����𫪪����:���Z:���Z鯪�Z�VUU�UUU�UUU�VUU鯪�Z鿪�Z鼪�Z:����:𫪪���� ���  ��  ��  ��� ����������?��U�>��U����U����U����U����U�ꫪU�ꫪU�ꫪU��UUU:�VU�:�ZU����� ���  ��  ��  ��� ������������?����>k����k����kUU��kUUU�kUUU�kUU��k����k��������>����?�������� ���  ��  ��  ��� �����V���V��:�V��:�Z���Z���Z���Z���Z����Z����Z����VU���VU�>�VU�?������ ���  ��  ��  ��� ����𫪪����:���Z9�UUU�UUU�UUU�UU�ꯕ��ꯕ��ꯕ��꿕��꼖��:����:𫪪���� ���  ��  ��  ��� �������ZU�?�VU�>�VU����Z����Z����Z����Z�ꫪZ�ꫪZ�ꫪZ�ꬪZ�:��j�:��j����� ���  ��  ��  ��� ������������?����>���V����V����V����V��VUU�kUUU�kUUU�kUUU�l��V>����?�������� ���  ��  ��  ��� �����VU��VU�:�VU�:�Z���Z���ZUU�ZUU�ZUU��Z����V����VU���VU�>�VU�?������ ���  ��  ��  ��� ����𫪪����:�U�Z9�UUU�UUU�UUU�UUU鯕VZ鯕VZ鯕VZ鿕VZ鼖VZ:��V�:𫪪���� ���  ��  ��  ��� �������ZU�?�VU�>�VU����Z����Z���UU���UU��UU�ꫪZ�ꫪZ��VU�:�VU�:�ZU����� ���  ��  ��  ��� ������������?����>k��V�k��V�k��V�k��V�kUUU�kUUU�kUUU�kUUU�l��U>����?�������� ���  ��  ��  ��� �����VU��VU�:�VU�:�Z�U�Z�V�Z�V�Z�V�Z�V��Z�V��Z�U��VU���VU�>�VU�?������ ���  ��  ��  ��� ����𫪪����:���Z9�UUU�UUU�UUU�UUU鯕�Z鯕�Z�U�V�VUU�VUU:�jU�:𫪪���� ���  ��  ��  ��� �������jU�?�VU�>�VU���UZ����Z����Z����Z�꫕Z�꫕Z��UZ��VU�:�VU�:�jU����� ���  ��  ��  ��� ���������ZU�?�UU�>�UU��k��U�k��V�k��V�kUUU�kUUU�kUUU�kUUU�l��V>����?�������� ���  ��    � �      � �     � ��     ���    ���    ������   ������?   ������  �����   ��^UU�   ��WUU�   ��UUU�   ��UUU�:   �zU�U��  ��zU�Wժ��zU�Wժ: ��zU�Wժ �zU�U��  �zUUU�>   ��UUU�   ��UUU�   ��_Uի   �����:   �����:    �����:    쫾��;    <��: �    �  �                  � �     ���    ����:    ����� �  ������;  ������ ������� ������� ��~UUU� ��^UUU��  �^UUU�� �^U�U�� �^U�W��  �^U�U�: ��^UUU�: �^UUU�: ��^UUU�� ��^UUU�� ��^U_U���^U{U�� �^��U�:  ������: �������� ������� ������  ��Ϊ�   ���   0 ;                                    ;  �     ; �     � ���   �ϫ��?   ����� �������  ������  �������� �������? ��WUU�� ��UUU�� ��UUU�� �zUU����zUU��� �zUUU��  �zUUU��  �zUUU�� �zUUU��� �zUU��� �zUUU�:  �zUUU�:  ��UUU�: �������� �������> ������� ������   �ê��:     ��:     <�;     � <       �     0       0 0�  0   � ��  ?   ��� �:   �Ϋ��:   ����ά   ������   ������   ������   �������� ��W�_�� ���U�W�� ���U�Wժ ��zU�Wժ  �zUUUժ>  �zUUUժ���zUUUժ�: �zUUUժ�� �zUUU���  �zUUU��   �zU�U�>   �zU�U�:  ���U�W�:  ��������  �������� �ê����� ?𪪪��?    뫺�    �>�Ϋ    ���    � � �    0 0     �                     0  �?���  ��?�?��������  ����  �������� 3�  ����  �������� 3�  �?��  ��?��������?��  ����  ���� ���� 0  ����  ��0�� ��� �  �?���  �������?��                                                                                                                          0  �  �  �             <                0                 0  � � �             0      0             0  �  �               �  <  <  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          H���� ��� ��� ��� � �[ ���\ ��� �\ �b �[ �a  �ܭ\ �q�� ��  ���\ �� ���� �ө�] ���^ ��� �\ �\ �b �[ �a ��� ���  ���^ �^ �^ �b �] �a �� �� ���  �ܭ^ �D0� ��  �ݭ� �� � ����� ��� ��  �� �ݭ\ �b ��� �[ �a ���  �ܭ[ i�[ �a  �ܭ] �a ���  �ܭ] 8��] �a  �ܭ] �� �݀����M  �䜦 �� hL� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                H�Z��J  �䩀�� �	�a �(�b � �ݩ(�� �N�� � �a �O�b ���  �ܩ�� ��� ��� �$�a �P�b �K��  �ܢ  �ܽ���c��� 轠��a  �ܩ���  �� �� ���ة�a ��� ��� �M��  �ܠ#����  �݈��  ��� �݀ ��  �� ]� a�z�hL��  ��    ��   ��   ���  ���  ����  �Ϗ�  ������ �����?   ����  ����   �      <    ���  ��� ���?  ���� �Ϗ�?  ������ �����?   ����   ����   �      <                 �   �  �� <� ��? �  � �� �� �? �> �> �? ��? ��0 �3                                                                       <                                      �0                                      �0                                      �                                      �                                      ��                                      p?�                                    \�                                    \7                                      \�                                      _]�                                     s]U                                    suU                                   ���W5                                   ��UU5                                   ��UU�                         ����     0 WU�                        � 0 �  ?  0 �WU                      �?�U�]�  0  \U                      <���4�0     pU                    ��? ��U     pU5                   <��  PW��     �U�                 00�3� UWUW��    �UU��                0��u�����_ٗ=    �UUUU5                �LW�?]U�U�W�     WUUU�                ��� ]U�UU��_�    WUUUU               �? WU]U�UU����    �UUUU               0QuWW����UW�i7�     ��_�               0@���   ����=0       p�                �� W���?CP��0       �W               �UUW3  0W]�o�3        �                �W�UW3�0W]]�y                        ������3�"0�����                        ��WU3�*0WUW��                       0w]UWU3 0WU�i�?                       ��]UWU3�
0WUש�?                        ������3 0������                        <tUW�W3�*0W_���                        |uUWUW3  0Wwݗ��        �             ����_3  0WW_���       

 � �          �����W3�
0WW�����    ������           �U����3�*0����j��*     ��� ��*   *    �U]��U3�*0W�������*�����* ���*  �����]UWU3�0��u��������������*����*�����T�/_WU3 �0W�U����������������* �"�
����Uuj���3 
0���o�� �  ��� � �������������_�/T�U3 0WWV�����(� ���"
� �r��.W�W3 0WW����? "�  �  (""*   pu�W�U3 �W_U���? � 
� � �  � �  ( pu�J���3) �����? ?�   �    
     ���JUwU3  Wu�ٮ�? �;0 8    � �  " �p��TU�_3
�*WUg���? �<0�           <  pU�S]WU3(  ו֦��?��00       �   � <P��U3  0WU������0�        0   �U�����3*(0�������0�           ��W���U3
0W]�����?  3        0     �����U3�Z__Y���W� �        0��    �W���U�U3�0W�^��_U�0 �   �     ��0   �_�����U3 0����_UU0   < �     ��0  0�}UU���3 0���WUUU� � � 0      �� ��uUUU��3�0�UUUUU���  0      �  0�wUUUUUU3�0WUUUUU�  �  0    �3  0��_UUUUU3�0WUUUUU= �< 0    ���3  0��_UUUUU3�0WUUUU� 3 0    pU<   ���_UUU�����_UUU�  03        p��� ���UU�U�T]UU�   0�� 0     <Q   � ��W�U�T]U�              �����       ��U�T��                ���          �U1�T     �              �?           ��3��    �                             0�                                   0�     �                                   �0     �                             �0                      3�                                00  3�                                       0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      H� jݩ�b ��a � �ݩ@�� ��b � �a �(�� �p�� ���  �ܩ��b �	�a � �� �� �� �ݮ  ����� �hLA�   �3             �                      00                                    00�0�  �0�  �� �����  �     0�0�0  �0 ? 30  030 3   <     000�3 � �3 �  �? �?�?��       0000   3    �0  000 0       000�0 �  �3 �  �0� �?���  ?                                                                                                                                                                                                                                                    0 0            �                      0     �?       0                      ?0<� 00���   00 ����  �0��      �000  00 33  0�0 00 3   �00      000� �?�33�  000 �?�3  �3 ��?      300 0  030   000 0 30 3 00�     �00�� ��30�  �00 ��� �3 ��?�                                      <                                                                                                                                                                                                                    0    < 0 �  0             �            0    0 0 �  0          �  �     � �0�000�3 ��0�  ?�?��� ��   30 �03000< �  3��<����<��   �30 �0030000 � �� ���������   30�  303<000 �03 � �����   ��� �00��?��?  �3�  ??�? ��                                                                                                                                                                                                                                                   <�        0         0 �  �       0         0         0 0   �       0 �0� ��� 0�0<���3 0 �� ��?   0  �0 <�� �0 �0� 03< � <��  <��   0 �3 � � 00�30�?30 0 ��  ��   0 3  � 00300030 0 ��  ��    ���3 � �? 00�30��?�? 0 ?�  <?                                                                                                                                                                                                                                                      0�    �  0 0                0�         �     0                  0�     �00<� �  ?0<� ����   ?� ��<��  �0�  00?  �000   030  �  0��   �0�  00  000� �?�?�  ? 0���  �0�0 00  300 0 000   � 0���  �00�  �  �00�� �?���?� ����<                                                                  �                                                                                                                                                                                             �        �                          �  �        �              � ���  � ��  ��� ����      30  0 30 �  30��   030      �30 �? �30 �  �?0�  �?�?�      30� 30  30 �0 3 ��0 000      ��� ��? ��  �  � �?��                                                                                                                                                                                                                                                   �3      0       0         0         0      0       0 �      0         0��?  ?0�  ���03�00��3 ���    ��030  �0 00�0303< 003      3030  00� �?� �3 3030 00��    3030 30  303 3 3<30 000    �00���  �00�  ��?�0�0 ��?�? ���                                                                                                                                                                                                                                                       �           0�<                                   0                  ?�� �  00�00 00< 0  ��� ���       0  0030 030 0  030 ��<      �? � �?30 030 0  �?�? ���    30   03< 030 0  30�0  ��      ��?�������? ����  �?0�  �             �                                      �                                                                                                                                                                                                       �   0  00                               �   0  0                         �00������3 �3<�����00             �30� 3< 0<00 003030             ���?� �30 000�00�?�?             �0 �000 000 030�0  0             �00�� ��? �?����0��<                                       <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               jݩ�J  ��@�� ��� �_�� �`�� ��a �@�b  �ܜ� �����a ��b � �ݩ�a �#�b � �ݩ�a �2�b � �ݩ �L��        ��?                    ����     ��            ����     g          �����?    �e<          ������    �Y�          ������    l�           ������    g�  �        �������   g�T         ���wUU�   ��t        �WuUUu   ���U       �[UUUUU   ��W        [UUUUU   �꿿       �WU����    ���       ����� �     �Z       ����?��     �V       ��� ��     �V        ��?���3     �V        ���0�0     �U        �?�@p     �U        0?  �      �Q        ��  �      pA        �  �      pA        ��\  ��      p         ��X���      p  0        �@ ?�      0  0        �  �        0        �  0        0        �: ��3        �        �:   0      [  �        {�  ?�   �? [  �       �U�@\  �k  �       _U�  W�� k P     �UP� U�_  �k P     pU  ��� U  �n P     \PU��� T  @� P    �WU�W��� T   @� P    �jU���{    @� T    ��VU���{     T  T    �VUUU�_      U  P    k@UU \     T�  �   �V  P@0   UAUi   �   �   U @ @UUU   �   0       @UU�
T  �             VU��BU@�            ����PUUU�       @   ���*U�Z��       @U  $ ���JU����   �   @UU  � ��jUU����   �T   TUU  P��UU����   �U TU�U  @�������     0YPU�VW  YԪ����      0�UUU�UW  d����?       0�VUU��W  �����       0�ZU�j�W  ��           0��Z�V�_  ��           0����V�~  ��           0P���U��U ��           0@��ZU��UUU��           � ��VU��jUU��           � TjU䪫UU��           � PUU����U�:           ��TUA������           ��TU������            �TU  P�����            �TV  @�����         0   ��V  �����        �   ��V  骪?�            ��Z  ��C�      � <   ��j �>T�      00    ��j��CU�<     0�    �k� �kUU��     ��    ���� Ô�U�!�   � �  ����3����0   <� �  <���03��j0   ���  0����?0��Z0�  �������?00�0�� ?�  <�0��< ��� Ϗ  0�� 0< ��+����  0 � ��  0� ������30�0 8 �    � ����<��<?� � ��    ��0��0��? � ��     �?�/�<���� � �     0� �������03� �     0� 0��<�� � ���    0�����3;��< ����0  ���,0��?3�>� 0�<0  ����?�3<�0��  ���? ����?3��?+��?� �?��<0 ���<<���0��?��?� ����<�<�0� ����<� ������<�?�?< <�< �  0��<���03 ��3�   � ���? �03���0� � �   �   �? �03����0 0 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         
�ʃ��J�
�F�d�������܀���6�T�r�����́��&�D�b�������ڂ���4�R�p�����                         .   /       (               )                                                                                                  *   +                             ,  -                            !                                                 &             '     $     %                       "                  #                           �$�B�`�~�����؄���2�P�n�����ȅ��"�@�^�|�����ֆ��0�N�l�    $     !         %                                                            &             '                 ,            -.            / "              #                                                                                    (                     )                 *             +                                                                                                                              Ƈ�� �>�\�z�����Ԉ��.�L�j�����ĉ� ��<�Z�x�����Ҋ���,�*                          +                                         .           /                                                                                      &         '                   (                 )   $               %                                                   !   "           #                       ,              -                                                             1 ���������:�X�v�����Ќ��*�H�f�������ލ���8�V�t�����Ύ�                                        *,       !   (+-           )                                                                                                  0      1                                                                           &                '                   $               %                   .             /     "                    #                                                 F�d�������܏���6�T�r�����̐��&�D�b�������ڑ���4�R�p�����	








		
	












				         			            				  

 	 0    1				 	


	

    	



	    	  				 	   	    ,	    	    	  


		 	  	    	-
   .	    	     		 	 	 	 	     /	    	    		 	 	 	 


	      	    	   	 		 	 	 	    		(	 	 		 
 
 	    	







)




 	 		     	   	              	 		 	&	      	 			 






'



     	 		



 			                 	 		     		
  	 		   		  		




 	








 

 	 	 		 		      	             	 	 		 
		     	       	 	 		  

      	     	



		 	 		    	 	    		 	 			   


 




 		
!   



 
 			             	
            			$  	   		




%	


 	 		"




	

 

		      	    
 

#	    	    		  	        	     	    		
 
	 

   	    	  	 	  *		   	      		   


 	 
 	  +		   			       	   	   														  0     0        �  �	  X	  \%  G   � �p��t�`U���H�o*p�*m�	
VQ*
U\*Z�^-h�ܧX���Zk�'V�/�S�*��
�E�DU�T�(��;je?���/Xi�.F�.�jU<H�B�hU����T�~��?Tu��W��Zѿ�U��Y�/�go�)��;?  ,   � �����?���  �  p  �:  ��  �� ��e���pfY���p�e=�����eY߿����[��_���so}�s�^�s�_p�up��pgY�p�e=�����eY�W���W���k���m�ٟ��ٳ��ٳ��ٰmy6��z6��u6��z6p�]6pVW6pYW6pe�5�����e gY |�  �� �_�������� �   0  <�  3� � ?���000<�00��<���3���?3 g� �UU\VY5he�9W�U�g5w�[?������Wߧ���<0<<�0�<��<���33���?�����UU\VY5�Yf9WUU�[e��g�e�WUU՗UV�g�Y�WUU�\Ye5\f�5\UU5l�U6�e�pUU�VY����*���
 � �03 �? ��������:���:���:���:���:���:���:��� ����?���                                                                  � �_ �� �� �� �_	  �  k �� �� p� p�
 p^ ��    \  � �W= ���  � �? ��  �� `7 `7 �W  �  ��  p9 p7 p= ��  � �� �� p5 \?< |�� ��� ��0�  �� �� 0w 0w `� �?  ��  0[ 0w �z �z p� �� p�  �5  �:  |� �� ��  ��  � � ��	 ��	 ��  �   � �l �� �| �[ 0�  � �W 0\ <�5 = �� ��  �?  |�  _� ��  ��  |� � �o������=���1��Z? �� ��  �_ �_��\��� �_  � �  _= ���  �/  77 �_= ��� p�� p'V|'vL�z��^�U�  �? ��� ��� �5������� �?   �  _= ���  V%  _=  _= ��� ��[pWUpWup_�5��9�W�3 �?������ �5������� �?   �?  |�  _� X�  |�  |�  �����pU�p]�\_�l���W��� ��_ �_��\��� �_  �        �?� �� �� ������� ����� ����� ���������                  � ��� �������U�\UU^UU������ ��
                        �� �0  0      ��3_5W=\�Wp\��                         �� WU WU3 WU3 WU3 WU ^���� ��* ��         �  p  �  0  0    0  0  �:  �5  �5  �:  0 �� ��
 �*  �<<�<<�<<�<<� ���0��?�?    <  �� �W� pU� �< ��  �� �pU�Up�U�WU |U5�WU5��� ��  ��       <  ��< pU� T� ��� ��<�pU�Up�UpUU�U5�UU5��������?�?<   �?  �� �U <0  �  �� �U�U�pUWpU�\U= \U���� �  �      <  <� �U �0 �� <�� �U�U�pUWpUU\U�\UU������� � �03  ����0�:�:��:���:�̫�;3���������: ��: ���������? � �03  ����0�:�:����ꬪ�ꬪ�����갪�����: ��: ���������? 03  ���� ���0����:����3;�:������ꫪ�:������ ��: �������? 03  ���� ���0����:�������:���:���:��������� ��: ���?��� � �03 �? ��������:���ꬎ�ꬺ�ꬪ��33���:��� ���������? � �03 �? ��������:���:���:���:���:���:���:��� ����?��� � �03 �? ��������:���ꬺ�ꬺ�ꬺ�ꬪ�갪�:��� ���������? � �03 �? ��������:���:���:���:���:���:���:��� ����?��� �?  �� ��������������� ��  �� ��0;���;�:�;�:���뫾�����? �?  �� ��������������� ��  ��  ��  ��  �:  �: �����*<<<< �  � �� ��Q�`Ռ1 �\�*���  ������t��{'" � 0z@�  @      �� �z�
�5��ի�zի�_իzUի^Uի^}ի^�լzU5��W ��          �? �W�pUU\UU5\�_5W�������7������7���7�?����7\�5pUU�W�����? �? �W�pUU\UU5\UU5WUU�WUU�WUU�_UU�{UU��W�ۜ��6\�j5pUU�W�����? �? �W�pUU\U�7\U�?WU??WU??W��?W5�?W�?W��\U�?\UU5pUU�W�?��� �? �W�pUU\UU5\UU5WUU�WUU�WUU�WUU�W�_�W���\U�:\UU5pUU�W�?��� �? �W�pUU�_U5�U5��U���U��?W��?\��p������U5\UU5pUU�W�����? �? �W�pUU\UU5\UU5WUU�WUU�WUU�WUU�W�_���zլjU5\UU5pUU�W�����? �  \5  \5 �\5?W���W]u�W�W�W6��W5\�|7�=��WpYe\�W5\5\5\5\5����?���������?�      <   �  ��  �<     �� W]5�0��Qu��^�ՠWu����/���
��
         �  � �03��3��00�?ï����0��������? �? ��0                � 000�� �� �>���� �� ���� �� ���?� � �  H��a �K�b � �� w� jݩ�a �K�b � �� w� jݩ�a �K�b � �� w�h`���� �
 �����`H�Z�\ i
��1�W ���X �[ i��W� �)Ɋ�%���!�5�Ƀ��^����� �� ����  ��z�h`���� ��H�Z�\ i
��1�W ���X �[ 8���W� �%Ɉ�!����W�����5�� �� ����  ��z�h`���� ��H�Z�\ 8���1�W ���X �[ i��W� �������
�� �� ����  ��z�h`���� ��H�Z�\ i��1�W ���X �[ i��W� �)���%���!��������<�� �� ����  ��z�h`���� ��H�Z���� �� 
����W 轖�X �[ JJme �i �\ JJJJmf �j � �W�c�L��ͬ ����Ȁ�ȱW�i ��ȱW�j ��ȱW���� �/��{ �{ �
�@��{ �P�1� ���G�0��� i�� �8�2��� i
�� �)�3��� i�� �� ��@�� �� ����	�� �� ���� �$� ��  ,� �� �ȩ�� ���M  ��z�h` �݀� �݀�H�Z�� 
����W ���X �� �W�c�N�� � �/��+������ �F�0�)�� �Z�"�\��!�� �]��_���� �8��9��:��W�� �Ȁ�z�h`H��[ �p�\ �	�� �� ��� �I�� ��� � �� �� �� �� �g �h �i �j �k �l �m �n �o �p �q �{ �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� � �e ��f � ��� �� �� � �� ��  �h`�� � � B���� ����� ��� G�� ��`�/�� �� �� �� �� �� �0�� �� �� �� �1�� �2�� �� �3�� �8�� �� �� �� �� �9�� �� �:�� �� �� �� �� �� �� ��� `Hک/�� �� �� �� �� �0�� �� �� �� �1�� �2�� �� �3�� �� ��F�� �����h`H�Z�/�� �� �� �� �� �� �1�� �0�� �� �� �� �� �� �2�� �� ��8�� �������:�� �����z�h`Hک/�� �� �� �� �0�� �� �� �� �� �2�� �� �� �3�� �@�� ��Z�� ������\�� ������h`Hک/�� �� �� �� �� �@�� �� ��� �0�� �� �2�� �� �� �� �3�� �1�� ��]�� �������_�� ������h`H�Z���b ��a �  �ݩ(�i ��j ���b � �a �b �1�U ���V �a �UI��U��i �i � ��(�i ��j �j � ���zh`H��� ��� ��� ���b � �a �� �
0	8�
�� �� iP��  �ܩ�a �� �
0�	�� iP��  �ܜ� h` �� � *�`H�� �_ �� �`  ���� ����� ��� ��� �
�� �	�� h`���� ��H�� �_ �� �`  ���� ����� �0�� 8��� ��� �
�� ��� h`���� ��H�� �_ �� �`  ���� ����� ��� ��� �
�� �	�� h`���� ��H��[ 038��[ +��\ 0#8��\ �� � ��� ��� � �
�� �	�� h`�� �� ���� ��H�[ �_ ��\ 8��` 4i�` 0,���� �#�\ �` ��[ 8��_ �[ i�_ 0���� h`� �� ��H�Z�[ JJme �i �\ JJJJmf �j � �'��c�Sͬ �������'��i �?�'��j �6�� �����{ �	�$��{ ��� z�h�� ������  �� ��LQ�z�h`L��H�� i�[ 0 8�	�[ �� i�\ 08�$�\ ���� h`H� jݩ����a ��b � �ݩ�a �-�b � �ݩ�a �F�b � �ݩ�a �U�b � �ݩ�a �i�b � �ݩ�a �x�b � �ݩ��� �P ���� �� jݩ�a ��b � �ݩ�a �-�b � �ݩ�a �<�b � �ݩ�a �K�b � �ݩ�a �Z�b � �ݩ�a �i�b � �ݩ�a �x�b � �ݩ��� �< ���� ��� ��h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���ة��  ��� � �u � � �v � �ύ& ��" t ����W ��X �� � �W����X ��� j�X �� ��L �H�Z�� �
0�� �	0�	�� �� L��� � �
�����$�� ���)�� �w�� ɠ��� �k�� ɀ��� �_�� �`��� �S�� �� ����� � ��� �=�� �0�� 8��� �+�� � ��	�� �� ��� � ��� i�� �� ����� z�(h@H�Z�' )��S ��� �� �ޭT �# �$ �% (z�hX@                                                                                                                                                                                                             ���t �ȍT �#  �ީ ��L �� �ݩ��� �
 �݈� �� jݩ ��L �� �ݩ��� �� � �݈� �� �� j� -�� �J  �� ,� �� �� �� �� �� X� ���� ����� � �& jݩ ��L �� �� jݩ �  ]� a� � L/� jݩ �� �  ]� a� 8�LQ©  ��L �� �ݩ��� �P �ݮ  ����� �� �� j� ]� a� � L/�Hڮ  ���
����  �݀q���
���  $ŀc���
���  �ŀU�����  NƀI���
���  �ƀ;�� jݩ �  ]� a��hL/	���� ����	����
���  qǀ�� I��h`����  �݀�Hک���  jݩ2�b ��a � �ݩP�b ��a � �ݩs�b �	�a � �ݩ�� ��� �*�b �
�a ��� �/��  �� �� �ݮ  ����� �� �ݜ� �h`�*�b �
�a ��� �/��  �ܩH�b  �� �� �ݮ  ��
�H�b  �܀����  ��L �� ��L��xHڭ� �r �� �s ����  �� �� �� jݩ�b ��a � �ݩ<�b ��a � �ݩ�a �� i��  �ީP�b ��a � �ݩ�a �{ ��  �ީd�b ��a � �ݩd�b ��a �� ���� �݀� �ݩ�b ��a � �ݮ  ��� �� �� �ݭr �� �s �� � ��  j� ,� �� �� ���hX`H�� ��M '��� � �q��k �f � ��\ �0�5 ��� �� ����� �\ 8��\  �� �ȩ���  ���k �Ҁ.�. �ܩ�� � �� �����  ٭l �� �ܩ � ��� h` �ܩ��  �� �݀�H�� �	�M n��� � �q��k �f ���\ �`�5 ��� �� ���	�� �\ i�\  �� �ȩ���  ���k �Ҁ.�. �ܩ�� � �� ���	��  �حl �� �ܩ � ��� h` �ܩ	��  �� �݀�H�� ��G ؠ�� � �k��k �e � ��[ ��/ ��� �� �	���� �[  �� �ȩ���  ���k �؀.�. �ܩ�� � �� �	����  vڭl �� �ܩ � ��� h` �ܩ��  �� �݀�H�� ��G ���� � �k��k �e ���[ ��/ ��� �� ����� �[  �� �ȩ���  ���k �؀.�. �ܩ�� � �� �����  Xڭl �� �ܩ � ��� h` �ܩ��  �ܩ���  �݀�H�� � �O �ǭ� 
��<��Y �<��Z �� 
��Y� �/m[ �� � �$ȱYm\ �� Ɉ ��� ����  �� � �Ȁ��� �� �� h`H��� �� �a �� �b �� ���� ��� �� i4��  �܀��� ��� �� i4��  �ܜ� h`H�Z�� 
����W 轡�X �� JJme �i �� JJJJmf �j � �


��W�c�Tͬ ���ȱW�i ��ȱW�j ��ȱW�7��� � �3���M  ��ȱW�� ȱW�c���� � �ȱW�� ��  ,� �� ��z�h`��� � � �ʭ� � � �̭� � � �έ� � � �ϭ� � � ��` �� �� � ��  �`H�Z� �

�����c�L��ͬ ��� �0L�ɭe i
�n ȹ���e 0��n �8�e 

�� �f i	�n ȹ���f 0��n �8�f 



�� �;�� ȹ��� ����������ͺ �;�ͻ �4�ͼ �-�ͽ �&�; � ��� �� � � �ʜ �� �� z�h`�� �� ���e i
�n ȹ���e 0a�n \�f i	�n ȹ���f 0J�n Eȹ��� �����������#ͺ ��!ͻ ��ͼ ��ͽ �	�; �� =ʀ�L�H �ʭ �>�� � �7�� �_ �� �`  ح� � �δ � �� �;��<�� ��;��  �� ��h`� �1�� �_ �� �`  �׭� � �� � �� �=��>�� �ǩ=�� ���� ���� ͺ �-ͻ �(ͼ �#ͽ �; ��� �a �� Ʉ�b �� ��  ��`H�� �B� �ѭ� ���+�� Ϳ �,�� �'�� �"�A�� �_ �� �` ��  ��� �	�� �� �� h`�� Ϳ ���� ���� �� \ˀ�H �̭� �C0�E0b�G0L��L̭� �_ �� �`  �׭� � �-�� �$�� �B�&�� �� �$� �ѭ� ����� �� �� ��G�� ��� ��  �� !�h`�� �_ �� �`  ح� � �-�� � ��� �D�&�� �� �̩ �ѭ� ����� �� �� ���E�� ���� �� ���� �_ �� �`  Nح� � �8�� Ɂ�� �F�2�� �� �� �� �� L�˩ �ѭ� ����� �� �� L�˩A�� L���� �� �� �� �� L�˭� �_ �� �`  �ح� � �8�� � ��� �H�2�� �� �� �� �� L�˩ �ѭ� ����� �� �� L�˩C�� L���� �� �� �� �� L�˭� � ��a �� ɀ�b �� ��  ��`H�Z� �

��G��c�L��ͬ ���� �0L�ͭe i
�n ȹG��e 0��n �8�e 

�� �f i	�n ȹG��f 0��n �8�f 



�� �I�� ȹG�� ������������ �1��� �*��� �#��� ���� � ���� �	�� �� �� z�h`�� �� ���e i
�n ȹG��e 0a�n \�f i	�n ȹG��f 0J�n EȹG�� �����������#�� ��!�� ���� ���� �	��� �� H΀�L%�H �έ� �@�� �_ �� �`  �ح� � ��� �� �� �� �� �� �I��J�� ��I��  �� ��h`�� �:�� �_ �� �`  Nح� � ��� �� �� �� �� �� �I��J�� ���I�� ����� ���� � ��a �� Ʉ� ��b �� ��  ��`H�Z�h � �

��p��c�rͬ ���e i
�n ȹp��e 0��n �8�e 

�� �f i	�n ȹp��f 0��n �8�f 



�� �� �
+ȹp�� �� �B�� �=�� �8��?��� ��h �%�� �#�#ȹp���4 %Щ�� �h  �� %�LϜ� z�h`��� ������� �۩�� ����
 ѩ�� �� �Щ�� ���� �� �8�� �3�� �.�� Ɂ'��� �� �� �� �a �� �b ��� ���  �ܜ� `H��� � ���L�Э� i��b ��� ��� ��� �� ��� ��a  �܀4��/�a  �ܭ��� a������ ����a  �ܜ� h`���H��� �� i�
�b ��� ��� ��� �� ��� i�	�a  �܀'�	�$� �a  �ܭ	�#��� ��	�	�a  �ܜ� h`�$�	��H��� � ���L�ѭ� i��a ��� ��� ��� �� ��� i��b  �܀9�Ɉ�>�b  �ܭ��� a��Ʉ�� ���i��b  �ܜ� h`���������� ��H�Z
����W 软�X � �

��W�c�Wͬ ���e i
�n ȱW�e 0��n �8�e 

�_ �f i	�n ȱW�f 0��n �8�f 



�` ȱW�� ���� z�h`� �� ��H�Z� �

�����c�L��ͬ ���� �0L�ҭe i
�n ȹ���e 0��n �8�e 

�� �f i	�n ȹ���f 0��n �8�f 



�� �N�� ȹ��� �� ��� ��� � ���� � z�h`�� �� �� ����ȹ��� �� ��� ��� � ��L8�H �ӭ� �_ �� �` �� �[ 0�V ح� ����� �0:�� � �׭� ���6�� �$$�� �� �N�
�N��  �Ӏ�O��  �� {� ��h`�� �� �� ��� �\ 0�� �ح� ����� �� �� �� �� Nح� ��Ш�� �� �� �� ���� � ��a �� Ɂ�b �� ��  ��`H�� � �h�� �_ �� �`  �׭� ���R�� ��
�����A�� ��� ��� �� �a �� �b �?��  �ة���  �� �� �ܜ� �� ��  �� �� ��h`� � �	�  �� �ȭ� � �	��  �� �ʭ� � �	��  �� ͭ� � ���  �ϭ� � ���  ��`� � ��� � �δ  �� �ȭ� � �	��  �� �ʭ� � ��� �	��  �� ͭ� � ���  �ϭ� � ���  ��`�� ��� � ��� 8���  �� �ȭ� � ��� 8���  �� �ʭ� � ��� 8���  �� ͭ� � ��� 8���  �ϭ� � ��� 8���  ��`� � ��� i��  �� �ȭ� � ��� i��  �� �ʭ� � ��� i��  �� ͭ� � ��� i��  �ϭ� � ��� i��  ��`H�� � �L֭� �_ �� �`  �׭� ���o�� ��j�� ������������ ��� ��� ��� ��� �� �a �� �b �?��  �ة���  �� �� �ܜ� � �� ��  �� �� �� ��h`�� ��H�� � �f�� �_ �� �`  �׭� ���P�� ����	��
�� ��� ��� �� �a �� �b �?��  �ة���  �� �� �ܜ� �� ��  �� �� ��h`H�� � �L׭� �_ �� �`  �׭� ���l�� ��g�� ������������ ��� ��� ��� ��� �� �a �� �b �?��  �ة���  �� �� �ܜ� �� �� ��  �� ��  �h`�� ��H�� � �i�� �_ �� �`  �׭� ���S�� ��N�� ��	��
�� ��� ��� �� �a �� �b �?��  �ة���  �� �� �ܜ� �� �� ��  �� ��h`�� ��H��� ��� ���  �ܜ� h`�_ Ͳ $iͲ 0�` ͳ iͳ 0����  �ǜ� `� �� ��H�Z�` i��1�W ���X �_ i��W� �	� �� z�h`���� ��H�Z�` i��1�W ���X �_ 8���W� �	� �� z�h`���� ��H�Z�` i��1�W ���X �_ i��W� �	� �� z�h`���� ��H�Z�` 8���1�W ���X �_ i��W� �	� �� z�h`���� ��H��� ��� ���  �ܩ���  �ݩ��  �ܩ �H  q㜨 h`H�l �l ���l �f ��m  ,� ��h`H�l � ��l �f ��l �l ���l ��m  ,� !�h`H�Z��� � �d �f �p �� 
�� ��W � ��X �p 
��W�Y ȱW�Z � �c �e �o �o ��Y�� �d � �9�d0
8�d�0Lڜ� ���  �ۭc �$i�c �o �ŭd i�d �p ���m ���l 
��ʒ�� �ʒ�� ��l 
��ڒ�� �ڒ��  �ۭc �$�i�c �o Ll��p �d m� �d L?٭m ���l 
��Ғ�� �Ғ�� ��l 
��⒍� �⒍�  �ۭc �$�c i�c �o Ll� 0� ��z�h`H�l �l ���l �e ��m  �� \�h`H�l � ��l �e ��l �l ���l ��m  �� �h`H�Z��� � �c �e �o �f �p � �d �� 
�� ��W � ��X �p 
��W�Y ȱW�Z �o ��Y�� �c � �5�� ���  �ۭd ɀ��d i�d �p ���c �$i�c �o ��L{ۭm ���l 
��꒍� �꒍� ��l 
��򒍧 �򒍤  �ۭd ɐ��d i�d �p L���o �c m� �c L�� 0� ��z�h`H�Z�� �0$8���� 
����W m� �W �h ���i �X �
����W m� �W �h 轙�i �X �� �i �� �j �d �1�U ���8�>�V �c �W�U�W i�W �X i �X ��i �i � �୤ �i ��h i�h �W �j �j � бz�h`H�Z� �y ��z � �w �@�x � � �y-t �w��(���y i0�y �z i �z �w i0�w �x i �x �����z�hH��� ��� ��� �� �� �[ �a �\ �b  �ܜ� h`H� �t  �ܩ��t h`xHڭ� 
����W ���m� �X  ���hX`H�Z�� �i �� �j �b �1�U ���V �a �W�� �� ���� ��!���� U�� �� -t ��� Mt ��� QU�U�W i�W �X i �X ��i �i � Э�� �i ��j �j � Ѝ�i �j z�h`H�Z�W �@�X � � � �W����X ���z�h`�Z�� � ����� ���� ��z�`Hڭ  �����h`Hڪ���




�g ��)g �& �h`H���� ��b ��� ��� �[ �a  �ܜ� h`H�Z
������ 轱��� � ���$�'�a��[��d�8�7��  2�ȭ���ݩ���  �݀�z�h`xH�Z�� �[��%��a��$��d��&����W ���X ��g �b �1�U ���V �a �W-t �U�W ȲW-t �U�W ��g ���a �a z�hX`H�Z�)�JJJJ��  2ފ)��  2�z�h`� � � �  ]� a� � � � � � � � �* �G �O � ���H �S `� ���%�+ � ]�$ � �% �  ���+ �+ �& � 4� ���%�8 � a�1 � �2 �  ���8 �8 �3 � �� ���X� ���� � ]� � �	 �  �� ���� � a� � � �  .�� � �
 � ��� � � � �S ��� q� ��`� �� ȱ�	 ȱ�
 ȱ� ȱ� )
���� 轿� � )0� ȭO �	�����H Ȍ � � �
 � �L��  ��� �� � �� ��Ȍ � ���! �"�$ ȱ"�% ȱ"�& ȱ"�' ȱ"�( )
����) 轿�* �( )0�- ȱ"����H Ȍ! �+ �, �& � �� � � �M )����� �.  ��`�. �/�1 ȱ/�2 ȱ/�3 ȱ/�4 ȱ/�5 )
����6 轿�7 �5 )0�: ȱ/����H Ȍ. �8 �9 �3 � Ы� � � �M )��@К��� �!  4���� �� ȱ� ȱ� ȱ� ȱ� )
���� 轿� � )0�  ȭO �	�����H Ȍ � � � � Х�  ��� �� � �� ��Ȍ � ���J 
����K 轇�L �K� ȱK� `�J 
����K 轍�L �K� ȱK� `H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; � �8�� �� )0� Ȍ ����� � � �; � z�h`H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; �  �8��  �� )0�  Ȍ ����� � � �; � z�h`H�Z�' )?	@�; �' I��-; �; �, �)��( )@��J��; �; �- �8��- ��( )0�- Ȍ, �)����, �( �, �; � z�h`H�Z�4 )?	@�; �4 I��-; �; �9 �6��5 )@��J��; �; �: �8��: ��5 )0�: Ȍ9 �6����9 �5 �9 �; � z�h`� `� `�H ���S  q�`H�Z�H ���%�I ���H �O �I )?
��g�Q �g�R �P  ��z�h`�O �* �G `�P �Q�C ȱQ�= ȱQ�> ȱQ�D )
����@ 轿�A �D )0�E ȌP �? �B �C � ��S `H�Z�O ���L��= �F �C I�F )��F �B �@��D )@��J��F �F �E �8��E ��D )0�E ȌB �@����B �D �B �C )�; �I )����
�@����; �; �F �( �; �G ��* �G �? �? �> � ��z�h`H�Z�  ��  �� � �� �  �� � �� .� q��� z�h`H�Z� � �
� � ��N �M )?�N �Q�� �K�N 
����" ���/ 软�# ���0 �! �. � � � �M )�����  ��M ���  4� q�z�h` ��!� q�!� _
�!� d
�!� q�!� ��!� q�!� _
�!� d
�!� q�!� ��!� q�!� _
�!� d
�!� q�!� ��!� q�!� _
�!� d
�!� q�!� q�!� d�!� _
�!� G
�!� G�!� GP�!�     � K��� T��� _��� T��� d<�!� _
��� T
��� d<�!� q�!� d�!� _
�!� �
�!� ��!� �P�!� d
��� _
��� d<�!� d
��� _
��� d<�!� K
��� G
��� K<�!� K
��� G
��� K<�!�     � �(�#� �(�#� q(�3� q(�3� �(�#� �(�#� q(�3� q(�3� �(�#� �(�#� q(�3� q<�3� �<�!� �P���     � q(�3� q(�3� q(�3� q(�3� 
��� w
��� <�!� 
��� w
��� <�!� _
��� Y
��� _<�!� _
��� Y
��� _<�!�     � ��!� ��!� ��!� �<�!� ��!� q�!� d�!� _�!� ��!� �<�!� �!� q�!� <�!� ��!� ��!� ��!� �x�!�     � ��!� ��!� ��!� �<�!� ��!� ��!� �!� q�!� ��!� �<�!� ��!� ��!� �<�!� ��!� ��!� ��!� �x�!�     � KZ��� G�!� ?��!� ?�� ?�� ?�� ?��� K�!� _� � K�!� ?��!� �� �� �� _x�3� �� �� �� _<�3� �� �� �� _<�3� _<�3� _<�3� _<�3�     � _Z�!� T�!� K��!� K�!� K�!� K�!� K�!� _�!� �!� _�!� K��!� ��!� ��!� ��!� x�!� ��!� ��!� ��!� <�!� ��!� ��!� ��!� <�!� <�!� <�!� <�!�     �i��2     ��� /��     � ���� ���� ��� _��� K��� ?��� /���     � ���� ���� �������.���T���     � (��     �
	�
	�
�
�
	

�
	
	 �	�
	 �				�
	 ��������G���  ����  K�  ��  #�  ��  p�����p����������	���4�=�H�\���"\@�%h�ʕ�j���
�Z�����/!���(�h����(�h�.��Z�"��N�z�B�
n�6	�	�	6_�J���ʘ
�J���������
�J������(�h�(�x����(�h����(�h�����$&%�%���� �� �0�@�P�`�p�����ʓ
�J���ʔ
�iU ��J�
�J���ʓ
�J���ʔ
����G�p��     




c  
c	c
cc����R��,�        	   	 
         c 
	
	c 		

 c 	
c 

	


	c�����V�� /:  3/      :      2   /0 c0  / 02 /  00  / 	/2 c20 
3  3/ /0 :  / 00 c/2  / / 3/ 3/ / @/ 1/ c/@ /3 
/0 	3/ 0/ 2/ / c��������://3  :   20/cEEEEEEEEEEEEEEc02 3/30/:/ 00c2// //3/3//@/1c@/3/0//3/0/2/c      cD�[�r���  ����������   	
   ����������    $(,048< L KLKLKLKc���������(�7�G�U�a�m�x�~�������������������������!�&�LIFEaFORCE$AREA$DOLLAR$PAUSE$PLAY$EXPLAIN$PRESSaaSTART$VITALITYaaOVER$WELCOMEaTOaPLAY$PRESSaANYaKEY$TOaCONTINUE$DESINGEDaBY$PROGRAMMER$MUSIC$YINaYONGaQIANG$HUaXUaHUI$PICTURE$ZHANGaLI$BANaYONG$SPECIALaTHANKS$JIaYAaLING$POISONING$YES$NO$THEaEND$THANKaaaYOU$CONTINUE$END$CONGRATULATIONS$YOUaAREaAaVERITABLE$HERO$GAMEaaOVER$ 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p��������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  ��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                                                                                                                                                                                                                                                                                                                                                                                                                                                          S� �	�