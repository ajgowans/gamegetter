�(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �
                            �
       ���                          ��*       �j�
                          ��)       �j�
                          ���       �ZY
                          ���       �VY
                          ���       �VU
                          ���       �VU
                          `��       �VU
                          hU�    PU�VU	                          hU�     �VUY                         hU�      PUVUTUU                     XU�      @U U @                    �Z�             T                   �j�    P           P                  hi�    @        TU                   ji�          TP                     Ve�     @i   U                      Ve�
      �Y P                        Ve�
      �UU@V                         V��
      �jU�                     �  V�V*      �ZUU
                     p-  V�V*     ��VUU �?                  \�  V�V*     ��VUU: ��                 _�  VU�*     ��UU�9 ��                 W�  �U�*     ��UUU9 ��                 W���U�*     �UUU� l�                �V��VU�*     �UUU� l�                �V��VU��     ��UUU� lV~U              �V��ViU�     ���UU�\� @U             �U��V�U�     ��UU��Z   P            �U��V�U�    ��UU��k     U           �՗>�V�V�    �YUU����      P          p�U>�V�^�
    �UUU����       UUU        p�U>�UU^�
    �VU�j��Z@     @       p�U>�UU^�
    ��U�Z��jAA     TU        hUU�|UUZ�
    ��U�ZU�jU      P         hUU�UUZ�
    �UU�VU�ZU     @          hUU��UUY�
    �UU�VU�ZY   P           hUU��UU��
    �UU�UU�Z�UU              hUUU�UU��
    �UU�UU�Z�PUU             hUUU�UU�
    oUUeUU�Z�
                �UUU�UU�
   �[ZUUUU�Z�
                �UUUjUU��*   �[ZUUUU�Z�
                �UUUZUU��*   �ZZUUUU�j�
                �VUUZUU��*   �ZjUUUU�j�
                �VUUZUUU�*   ��jUUUU�j�
          UUT�VUUUZUUU�*   ��jUUUU�j�
         P T@�UUUUZUUU�*   ��jUUUU�jU
               TUUUjUUU�*   ��jUUUU�kU
               @UU�jUUU�*   ��jUUUU�[U
                UU�jUU��*   �VUUUU�[U*                @U�jUU���   �UUUUU�[U*         P         �UU�j�   ��VUUUU�[U)          T   P  ��VUUZ�  @��ZUUUU�[U)              �U�U��VUUY�  T ��UUUU�[U�
            @�U�U��VUUY�   ��VUVU�[U�*          P UU�U�U��ZUUe� P      U�ZU�&          @U  �V�U��ZUUe� P     �VUeZU��              �Z�U��jUU��     jUUUeZUe�              �Z�U�V�UU��   �jUUUUZUe�              �V�U�V�VU��P   �VUUUUiUU�             ���V�V�VU�� PU��UUUUiU��             �Z�V�VUZU��
 P�着jUUUiU��             �V�V�UUYU��
  ��VUZUUUiU�U             �U�W�UUUU��
  ��UU�UUUiU�V             �U�W�VUUU��*  ��UUUVUUiU�V            ��U�W�VUUUU�*  �UUUZUUiU�Z            �jU�V�VUUUU�*  �UUUjUUiU�Y
            ��UU^iUUUUU�*  �[UUUiUUiU�Y
            ��UUj�_UUUU�*  �ZUUUiVU�U�U
            ��UUY�_UUUU�*  �ZUUU�UU�U�U	            ��UUY�_UUUU�*  �ZUUU�VU�UUU	            ��UU��~UUUU�*  �ZUUU�ZU�UUU)            ��UU���UUUU��  �ZUUU�ZU�UUU)            ��VU���UUUU��  �ZUUUUjUUUUU)            ��VU�j�UUUU��  �ZUUUUiUUUUU%            ��VU�ZUUUUUU� ��ZUUUUiUUUUU%            �iVU�ZUUUUUU� ��ZUUUU�UUUUU%            �UVU�VUUUUU�� ��VUUUUeUUUUU�            �UU��VUUUUU�� ��UUUUUeUUUUU�            �UU��VUUUUU�� ��UUUUUUUUUUU�           �UU��VUUUUU�� ��UUUUUUUUUYU�           j�UU�VUUUUU�� ��VUUUUUUUUYU�          �jUUU�WUUUUU�� ��VUUUUUUUUjUU
          �jUUU�UUUUUU�� ��ZYUUUeUU�jU�
          �jUUU�eUUUUU�� ��[eUUU�UU�jU�*          �ZUUUieUUUU������[�UUUuUU��U��         ��jUUUYjUUUU������j�~UU�VU��U��
��   �
����VU���VUU�����꿪��ꫪU�����k��jU���V���jU��jU�����UUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUU��? WUU�?<\UU� pUU�? pUU��0pUUU��_UUU=? \UUU� WUUU���_UU�? ��UU�� ��WU����W]�����Wu���Wu  Wu���Wu�����U�U���WUU����WUU}���WUU�� UU5 � �UU �  WU�����WUUUUUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUU��? WUU�?<\UU� pUU�? pUU��0pUUU��_UUU=? \UUU� WUUU���_UU�? ��UU�� ��WU����WU�����WU���WU  WU���WU�����U�U���WUuU���WUuU� WUu�� Uu5 � �U]�����W'UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUUUUUUUUU_UUUU�WU_UU��\U_UU���\U_UU�� \U_UU��WU_UU�� W�_U��? W�WU�?<\�WU� p�WU�? p�WU��0p�WUU��_�WUU=? \�WUU� W�UUU�����UU�? ���UU�� ���UU�����U]������Uu���W�Uu  W�Uu���W�Uu����W}U�U���W}UU����W}UU}���W}UU�� UU5 � �_UU �  _UU�����_U'UUUUUUUUUUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUUUUUUUUU_UUUU�WU_UU��\U_UU���\U_UU�� \U_UU��WU_UU�� W�_U��? W�WU�?<\�WU� p�WU�? p�WU�� p�WUU��_�WUU=?0\�WUU� W�UUU�����UU�? ���UU�� ���UU�����UU������UU���W�UU  W�UU���W�UU����W}U�U���W}Uu����W}Uu}� W}Uu�� Uu5 � �_U]�����_UUUUU�_UUU��?pUUU���sUUU��pUUU �_UUU��\UUU�� \UUU�<�pUUU?< �UUU� �UUU���UUU=�UUU�� pUUU�? \U]U���WUuU� \UuU��pU�����_U�����_U�50��UU7�  �UU����WU]����UU����?_UU�?�pU����pU5 _� \U� |� WUUpU�UUU�_U}UUUUU�UUU��WUU�??WU��? WU� ��UU��?�UU���UU��WU�� \U�� \U��?\U��?�WUU� WUU��UuU��U�U� �U�U��W�����U��?��UU����WU��\U��?\UW��WU���WUu���_U���U5 _�U5 p�U� p�UU�_�UUUU�_UUU��?pUUU���sUUU��pUUU �_UUU��\UUU�� \UUU�<�pUUU?< �UUU� �UUU���UUU=�UUU�� pUUU�? \U]U���WUuU� \UuU���pUu���?_U���?�\U�5���sU�5� ��UU�\��WU}��? WU�����\U5���?pU5���pU5�� \U5pU� WU5\UU�UU�WUU}U	UUUUUU�_UUUUU��?pUUUUU���sUUUUU��pU_UUU �_UUUU��\U�UUU�� \U�WUU�<�pU�_UU?< �UUUU� �UU�UU���UU�WU=�UU�_U�� pUUUW�? \UUU�U���WUUU�W� \UUU�_��pUUUu���_UUUu����_UUUu50��UUU�5�  �UUU��<��WUU�U����UUUU����?_UUU}���pUUU� ?�pUUU5 �� \UUU� �� WUUUU�_�UUUUU�_}U
UUU�_UUUUUU��?pUUUUUU���sUUUUUU��pUUUUUU �_UUUUUU��\UUUUUU�� \UUUUUU�<�pUUUUUU?< �UUUUU� �UUU�U���UUU�WU=�UU�UU�� pUU�WUU�? \U�UUUU��WU�WUUW� \�UUU]��\�WUUUu����UUUUu���WUUUU]����UUUUU]�0�WUUUUW=��UUUUUW5��UUUUUW���UUUUU]����UUUUU�=���WUUUUU�5 _UUUUU 7 \UUUUU5 7 \UUUUU����WUUUUUUUU�_UUUUUUU��?pUUUU_UU���sUUU�_UU��pUUU�WUU �_UUU�UUU��\UUUUUU�� \UU�_UUU�<�pUU�WUUU?< �UU�UUUU� �UUUUUU���U�_UUUU=�U�WUUUU�� pU�UUUUW�? \UUUUU]���W�_UUUU]� \�WUUUUW���p�UUUU����?_UUUU���?��_UUUUu5����WUUUUu5� ��UUUUUu���WUUUU�u��? WUUUUU�����UUUUUU5���?WUUUUU5�?� \UUUUU5��� \UUUUU5p�7 WUUUUU5\���UUUUUU�W}UUUUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUUU�0pUUU?��UUU�< \UUU�� WU�U����Wu���\u��� \]��??W]�?��U]����WUu}��?WU������UU�?�WU���� WU5��3 WU��UU�W5pUU5�U�_UU5 WUUUU��UUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUUU�0pUuU?��_U�U�< \UUW�� WUU]����WU]��\U��� \U����?WU����UU��UUU5��_UU���U�����U��?�U��_��U}�WUpUUUUU=\UUUUU�WUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUuU�0pU�U?��_UUW�< \UUW�� WU�U���UU�U���UUu����Wu����0\�� �?�\U��?<�WU�����UU�����UUU��?UUU}��_UUU�0pUUUU��UUUU��UUUU�UUUU_�UUUUU��uUUUUUuU_UUUUUuUUUUUUU�UUUUUUU�_UUUUU�?��UUU�?���UU�?�?��UU�?���WU����W�������W5�?����W5���� �W5���  W5��� 0�_5����0�\�3�0 �\5�\3�\5�\=p�W5�W�_UU�W�\UUUUUU5\UUUUUU�WUUUUU�WUUU�� \UUU�� pUUUU�UUUU��_UUU?��UU�����UU�����UU� ��U� �<��U����UW�=���UWU����UU���_�UU5��WuUU �_uUU���UU�|UWU |UUU UUU�UUU5 �UUU5��_UUU�� \UUU��_UUU���WUUU��UUUU�_UUUUUUUU�WUUUUUU5\UUUUUU5��WUU�W��7\�_|5�\5��5�\53 ���W53��3\�3 ��\�0  ��\�� ���\������\������?W������U�����wUU�?���_UU����_UUU�_��WUUUUU��UUUUUUU_UUUUUUU]UUUUU�U]UUUUU]_WUUUUUW�UUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUUU�0pUUU?��_UUU�< \UUW�� WUU]����WU]��\U��� \U���?W�� ���U�� ��UU�U�UUUW���WUU]���_UU���?UUUU���_UUU�?�pUUU��pUUU� 0pUUUU\UUUU��W&
UUUUUUU�WUUUUUU��\UUUUUU���\UUUUUU�� \UUUUUU���WUUUUUU=�WUUUUUU� WUUUUUU<<\UUUUUU�? pUUUUU��� pUUUUU�3�3pUUUU��=��_UUUUU��\UUUU�_�� WUUUU�w���UUUUU�u��WUUUU]��?WUUU�_]���UUUU�Wu�?�UUUU�U���UUUUUU����UU�_UU���WU�WU�?�� WU�jU5��= WU?�U�s�U��V�_5pU�jU�W�_U� �U5�UUUU?��V�UUUU �UUUUUUU �jUUUUUU	��ZUUUUUU� 
hUUUUUUU��UUUUUUU) �ZUUUUUU�
 hUUUUUUU�*�ZUUUUUUU��UUUUU-UUU�|UUUUUUUUU	|UUUUUUUU�|UUUUUUUU% |UUUUUUUU	 |UUUUUUUU
�UUUUUUU���UUUUUUU%� �UUUUUUU	( �UUUUUUU	*�UUUUUUU�

�WUUUUUU�	��WUUUUU�`���WUUUUU�h���WUUUUU%X�j�WUUUUU%��Y�WUUUUU%��U�WUU�WU���U�_��\U��UUU_���\Ui�UUU_�� \UYUUUU_��WUYUUUU_�� WUUUUUU_�? WUUUUUU?<\UUUUUU} pUUUUUU��? pUUUUUU�0pUUUUUU���_UUUUUU�3 \UUUUUU��� WUUUUUU����UUUUUUU���WUUUUUU���?WUUUUUU����UUUUUUU��?�UUUUUUU���UUUUUUUU����UUUUUUU���WUUUUU�?�� WUUUUU5��= WUUUUU�s�UUUUUU�_5pUUUUUU�W�_UUUUUU5�UUUUUUUUU�UUUU.UUUUU�VUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUUU)�UUUUUUUUU� ZUUUUUUU�

�UUUUUUUU)� ZUUUUUUU�
`UUUUUUU�
  UUUUUUUU� �UUUUUUU�
�UUUUUUUU* UUUUUUUU��_UUUUUUU��WUUUUUUUU*�UUUUU�WUU�UUU��\UU�_UUU���\UU�WUUU�� \UU�UUUU��WUUUUUU�� WU�_UUUU�? WU�WUUUU�<\U�UUUUU? pUUUUUU<0p�_UUU�U��_�WUUUUW?��P�UUUUU]�< _UUUUU]����_UUUUUW����WUUUUUW��?�UUUUU�U���|UUUUU�U����UUUUU�U��WUUUUU��� WUUUUU����UUUUUUU���UUUUUUU���_UUUUUUU���pUUUUUUUU��UUUUUUUU�pUUUUUUUUU\UUUUUUUUUWUUUUUUUUU�UUUUUUUUU�UUU��WUU�??WU��? WU� ��UU���UU����UU��WU���\U�� \U��? \U��?�WUU� WUU��UUU��UUU� �UUU��W�������?�������������� �������_U��?WU����WUuU��|UuU�?�U�U��UUWUpUUUU�_UUUU�_UU��?pUU���sUU��pUU��_UU�� \UU�?�\UU�<0pUU?<��UU� �UU��UU=�UU���pUU�? \UUU��WUU� \UU��\UU��?pU��?�_U5���_}5���_�5�  ��������U�����W_�����U���
UUUUUUU�WUUUUUU��\UUUUUU���\UUUUUU�� \UUUUUU��WUUUUUU�� WUUUUU��? WUUUUU�<\UUUUU� pUUUUU�?0pUUUUUU���UUUUU�?��PUUUU]���_UUUUu����WUUUUu5��WUUUU�_��\UUUU�W�??pUUUU�U���_UUUUU���_UUU��U���_UUU��U���WUUU�UW5 �UUUUU]���WUU�_U����_UU�WUU���UU�UU����UUUU5 _� W�_UU5 \5 \�WUU�p5 \�UUUU�_��W.UUU�|UUUUUUUUU	|UUUUUUUU�|UUUUUUUU% |UUUUUUUU	 |UUUUUUUU
�UUUUUUU���UUUUUUU%� �UUUUUUU	( �UUUUUUU	*�UUUUUUU�

�WUUUUUU�	��WUUUUU�`���WUUUUU�h���WUUUUU%X�j�WUUUUU%��Y�WUUUUU%��U�WUU�WU���U�_��\U��UUU_���\Ui�UUU_�� \UYUUUU_��WUYUUUU_�� WUUUUUU_�? WUUUUUU?<\UUUUUU} pUUUUUU��? pUUUUUU�0pUUUUUU���_UUUUUU�3 \UUUUUU��� WUUUUUU����UUUUUUU��? WUUUUU����\UUUUUU����sUUUUUU�����WUUUUU����\UUUU�U5  \UUUU�U���<\UUUU�U����WUUUUU����_UUUUUU}��UUUUUU����UUUUUU5 _� WUUUUU5 \5 \UUUUU�p5 \UUUUUU�_��W.UUUU�jUUUUUUUUU��ZUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUU�
�UUUUUUUU�� ZUUUUUUU�
�UUUUUUUU*� VUUUUUU��  PUUUUUUU�
 _UUUUUUU� �_UUUUUUU��WUUUUUUU�
�UUUUUUUU) UUUU�_UU��_UU��?pUU��WUU���sUUU�UUU��pUUUUUU �_UU�_UUU��\UU�WUUU�� \UU�UUUU�<�pUUUUUU?< �U�_UUUU� �U�WUUUU���U�UUUUU?�UUUUUU�� p�_UUUUU��\�WUUUUU���W�UUUUUU�� �UUUUUW��?0pUUUUU]���3pUUUUU]����pUUUUUu���_UUUUUu���\UUUUU��  \UUUUUU����WUUUUUU���UUUUUUU����UUUUUUU���WUUUUU� |�\UUUUU� p� pUUUUUU�� pUUUUUU�U�_UUUUU,UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU_UUUUUUU_UUUUUUU_UUUUUU�_UUUUUU�WUUUUUU�WUUUU�U�WUU��W�UUU�??W�UU��? W�UU� ��U}UU��?�U}UU���UUU��W_UU�� \_UU�� �_UU��?�WUU��?��WUU�� �WUUU���UUuU��WU�U� �WU����WUu=����UUu��?sUUu���sUU�5< ��UUU�����_UU=����pUU����?�UU3�?��UU�����UU0��UU�  �UU�    UUU����UU'UUUUUUUU�UUUUUUUU��WUUUUUUU�??WUUUUUUU�? WUUUUUUU���UUUUUUUU<�UUUUUUU��UUUUUUU�?WUUUUUU��? \UUUUUU��? \UUUUUU���\UUUUUU��WUUUUU�_=� WUUUUU�W�?�UUUUUU�]��UUUUUU]���}UUUU�_W���UUUU�WW����UUUU�U]���UUUUU�5 �UUU�_UU���UUU�WU�����_UU�UU���?pUUUU����?�UկVU3�?��U��ZU�����U� hU0��U?�VU�  ���ZU�    �jUU����U� �ZUUUUUUU  �VUUUUUU� 
�UUUUUUUU
��VUUUUUUU% 
ZUUUUUUU���UUUUUUUU� �VUUUUUUUU��UUUUUUUUU�ZUUUUU/UUUUUU�UUUUUU� ZUUUU�  PUUU� � �UU� � �UU
�
  �U��Z�
�U�ZU�� |UZUUU
 |UUUUU) |UUUUU�
|UUUUUU
_UUUUU�*_UUUUUU�_UUUUUU�_UUUUUU�WUUUUUU�WUUUU�U�WUU��W�WUU�??W�UU��? W�UU� ��U�UU��?�U�UU���U}UU��W}UU�� \}UU�� \UU��?\_Uu��?�W_U��� W_U�U���_UuU���WU]U����WU]����WU]�����WUu� ���UU������UUU�����UUU����3_UU����pU�0�?�pU�<�?0pU�0�?�pU�� �?pUU�  \UU=   �WUU����UU+UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�UUUUU�U�_U�U5��U�U���W�U���W�U��?\�U? �_������5�����������������5���������?�U�����U��?��U? ��������������5?��_�5�?�s��0|���?�����?p����30< �����0���  ��    U����U UUUUUUU�UUUUUUU�UU�UUUU��WU�_U���_U�WU���_U�UU��pUUU�  �_UU����WUU�����UU����?UU5����_UU5����\UU5����\UU���?�WUUU��?�UUUU����WUUU5���WUUU����WUUU�?�WUUU����UUU�����UUU����UUUU?���UU������UU����WU��� WU? �?0WU�0�WU�?   WU�    �UUU����_UU'	U�WUUUUUUU�_UUUUUUU	UUUUUUU�UUUUUUU�WUUUUU� �_UUUUU��UUUUU%�UUUUU%� �WUUUU	����_UU���U?��UU�hVU���WU�hVU���WU�ZUU��?\UbZUU?�_UbYUU���_UiUU����UiUU5����UeUU�?�?WeUU����WeUU���WUUU5��� WUUU���� WUUUU����UUUUU��?�WUUUU? ��_UUU����UUU���<�UUU5�?�s�UUU5<0|UUUU��?��_UUU=���?pUUU����UUU0< �UUU� ���UUU0��UUU�  �UUU=    |UUU�����W.UUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WUUUU�WU�_�WU5���WU����WU����WU��?�WU? ��WU���?W����?\5����\���_���W���W5����W�����WU����WU=  �WU����W�����W�?���W5�?��W50|U��?��_��?p����30< �����0���  ��    U����U+UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU_UUUUUUU_UUUUUUU_UUUUUU�_UUUUUU�WUUUUUU�WUUUUUU�WUUUUUU�UUUUUUU�UUUU�_U�UU��?pU}UU���sU}UU��pUUU �_U_UU��\U_UU�� \�_UU�<�p�WUU?< ��WUU� ��WUU���UUU=���UUU��0p�UUu�? \}UU����WUU��? �_UUu��?0pUUu��pUU]��?_UU]���UUUu �}UU������WUU����?\U�0?���pU��� sU�0��pU��� pU� < � pUU?   �_UU����UUUUU�UUUUUUUU��WUUUUUUU�??WUUUUUU��? WUUUUUU� ��UUUUUU����UUUUU������UUUUU�_��WUUU��U���\UUU�_U�� \UU��UU��? \UU�_UU��?�WU��UUUU�WU�_UUUU��U��UUUUU��U�_UUUU]� ���UUUUUW�?��_UUUUU����UUUUUU����_UUUUUU����sUUUUUU�����wUUUUU� �3�UUUUU� ��WUUUU���WUUUU���<WUUUU��WUUUU   � WUUUU�   �UUUUUU����WUUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUU��? WUU�?<\UU� pUU�? pUU�� pUUU��_UUU=?\UU]� WUUu���UUUu� �WU]��\U]���\U� ���WU� �?UU]��_Uu�����U�����W5���3\5��?�\5� <\5�< �\5  < \�   �WU����_UUUUUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�? WUU��3WUU�?\UU�3pUU�? pUU�� pUUU��_UUU=?\UUU� WUUU���UUUu� WUU]�� WUU]��\UU]���UU]����UUu����U���0W5��?0\5��?0\5���?�\5�?�?\5   �\�   �WU����_U}}����z�^�WUU}��}0?�                                                                                                                                                                              �(                                        TQEDUTTUQED ET          DA DDUUTTEDU             ����                           ����*                           ������                        ��  �*  @         TUUEUUDUUEUUE �*TeU���  TUEQTUETUEQTU            ��BUeU�*        @              @  �*TUeUU��"   @                  @ ��BUUeUU��   @   @               @ ��TUUeUU�*      @     UEEPUAUUUU�*UUAeUU�*AAUUAUUU@UEE       @   �JUU eTU��     @                 �JUUAeUU��                     @  �RUUUeUUU�    @              @   �VUUUeUUU�      @      PUUAUUUUE�RA e@� QQEUUUUPUUA  P   @      �V �*e�J�          P   @  @     �VA�*e�J�  @       @   @  @     �RU�*e�JU�  @       @   @        �VUJe�RU�  @        @ QUUUUTUUUP�VUJe�RU�TUUUTUUQU  @    @   �RU�*e�JU�             @    @   �VU e@U�             @    @   �VAUUeUU�             @     @   �R UUeUU�           PUAUUUUUU  �VAUUeUU�  TUUUUPPUA           �VUUPeTU�  @                    �RU@ePU�  @     @               �VUUPeTU�                          �VUUUeUUU�                             �����������              ���������������BUUUUUUU����������������              �@UUUUUUU(                              @UUUUU                UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                 UUUUU                                  UUUUU                                  UUUUU                 UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                  UUUUUUUUUUUUUUUUUUUUUU                              UUUUUUUUUU                              UUUUUUUUUU@UUUUUUUUUUUUUUUUU            UUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@                UUUUUUUUUUUUUUUUUUUUU@                          @UUUUUUUUUU@                          @UUUUUUUUUU@                          @UUUUUUUUUU@ ��  ���
  ���*          @UUUUUUUUUU@           ����  ��� @UUUUUUUUUU@              �  � � @UUUUUUUUUU@  ���  ���
  �   �  � � @UUUUUUUUUU@  VUU  XUU	  `*  ���� � @UUUUUUUUUU@  VUU  XUU	  `%  �UU� � @UUUUUUUUUU@ �VUU���ZUU���j%  �UU� � @UUUUUUUUUU@  VUU  XUU	  `����UU�
� @UUUUUUUUUU@  VUU  XUU	  `%  �UU�� @UUUUUUUUUU@ �*���  ���
  �%  �UU�� @UUUUUUUUUU@               *  ������ @UUUUUUUUUU@ ��������������       � @UUUUUUUUUU@               �������
� @UUUUUUUUUU@ �*                    � @UUUUUUUUUU@ V%                    �� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ �*                    X� @UUUUUUUUUU@                      �� @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@ �*                    � @UUUUUUUUUU@                      �� @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@ �*                    � @UUUUUUUUUU@ V%                    �� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ V%                    X� @UUUUUUUUUU@ �*                    �� @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@                      � @UUUUUUUUUU@               ����  � @UUUUUUUUUU@               �     � @UUUUUUUUUU@               �     � @UUUUUUUUUU@               �   ���
� @UUUUUUUUUU@               �   VUU	� @UUUUUUUUUU@               �   VUU	� @UUUUUUUUUU@               ����VUU�� @UUUUUUUUUU@ �*             �   VUU	� @UUUUUUUUUU@               �   VUU	� @UUUUUUUUUU@               �   ���
� @UUUUUUUUUU@                       � @UUUUUUUUUU@ �*                     � @UUUUUUUUUU@ V%                     � @UUUUUUUUUU@ V%             DUTUQQ� @UUUUUUUUUU@ V%              @  @ @ � @UUUUUUUUUU@ V%             'UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUUUUUUUUU_UUUU�WU_UU��\U_UU���\U_UU�� \U_UU��WU_UU�� W�_U��? W�WU�?<\�WU� p�WU�? p�WU��0p�WUU��_�WUU=? \�WUU� W�UUU�����UU�? ���UU�� ���UU�����U]������Uu���W�Uu  W�Uu���W�Uu����W}U�U���W}UU����W}UU}���W}UU�� UU5 � �_UU �  _UU�����_U'UUUUUUUUUUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUU}UUUUUUUUUUUUUU_UUUU�WU_UU��\U_UU���\U_UU�� \U_UU��WU_UU�� W�_U��? W�WU�?<\�WU� p�WU�? p�WU�� p�WUU��_�WUU=?0\�WUU� W�UUU�����UU�? ���UU�� ���UU�����UU������UU���W�UU  W�UU���W�UU����W}U�U���W}Uu����W}Uu}� W}Uu�� Uu5 � �_U]�����_UUUUU�_UUU��?pUUU���sUUU��pUUU �_UUU��\UUU�� \UUU�<�pUUU?< �UUU� �UUU���UUU=�UUU�� pUUU�? \U]U���WUuU� \UuU��pU�����_U�����_U�50��UU7�  �UU����WU]����UU����?_UU�?�pU����pU5 _� \U� |� WUUpU�UUU�_U}UUUUU�UUU��WUU�??WU��? WU� ��UU��?�UU���UU��WU�� \U�� \U��?\U��?�WUU� WUU��UuU��U�U� �U�U��W�����U��?��UU����WU��\U��?\UW��WU���WUu���_U���U5 _�U5 p�U� p�UU�_�UUUU�_UUU��?pUUU���sUUU��pUUU �_UUU��\UUU�� \UUU�<�pUUU?< �UUU� �UUU���UUU=�UUU�� pUUU�? \U]U���WUuU� \UuU���pUu���?_U���?�\U�5���sU�5� ��UU�\��WU}��? WU�����\U5���?pU5���pU5�� \U5pU� WU5\UU�UU�WUU}U	UUUUUU�_UUUUU��?pUUUUU���sUUUUU��pU_UUU �_UUUU��\U�UUU�� \U�WUU�<�pU�_UU?< �UUUU� �UU�UU���UU�WU=�UU�_U�� pUUUW�? \UUU�U���WUUU�W� \UUU�_��pUUUu���_UUUu����_UUUu50��UUU�5�  �UUU��<��WUU�U����UUUU����?_UUU}���pUUU� ?�pUUU5 �� \UUU� �� WUUUU�_�UUUUU�_}U
UUU�_UUUUUU��?pUUUUUU���sUUUUUU��pUUUUUU �_UUUUUU��\UUUUUU�� \UUUUUU�<�pUUUUUU?< �UUUUU� �UUU�U���UUU�WU=�UU�UU�� pUU�WUU�? \U�UUUU��WU�WUUW� \�UUU]��\�WUUUu����UUUUu���WUUUU]����UUUUU]�0�WUUUUW=��UUUUUW5��UUUUUW���UUUUU]����UUUUU�=���WUUUUU�5 _UUUUU 7 \UUUUU5 7 \UUUUU����WUUUUUUUU�_UUUUUUU��?pUUUU_UU���sUUU�_UU��pUUU�WUU �_UUU�UUU��\UUUUUU�� \UU�_UUU�<�pUU�WUUU?< �UU�UUUU� �UUUUUU���U�_UUUU=�U�WUUUU�� pU�UUUUW�? \UUUUU]���W�_UUUU]� \�WUUUUW���p�UUUU����?_UUUU���?��_UUUUu5����WUUUUu5� ��UUUUUu���WUUUU�u��? WUUUUU�����UUUUUU5���?WUUUUU5�?� \UUUUU5��� \UUUUU5p�7 WUUUUU5\���UUUUUU�W}UUUUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUUU�0pUUU?��UUU�< \UUU�� WU�U����Wu���\u��� \]��??W]�?��U]����WUu}��?WU������UU�?�WU���� WU5��3 WU��UU�W5pUU5�U�_UU5 WUUUU��UUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUUU�0pUuU?��_U�U�< \UUW�� WUU]����WU]��\U��� \U����?WU����UU��UUU5��_UU���U�����U��?�U��_��U}�WUpUUUUU=\UUUUU�WUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUuU�0pU�U?��_UUW�< \UUW�� WU�U���UU�U���UUu����Wu����0\�� �?�\U��?<�WU�����UU�����UUU��?UUU}��_UUU�0pUUUU��UUUU��UUUU�UUUU_�UUUUU��uUUUUUuU_UUUUUuUUUUUUU�UUUUUUU�_UUUUU�?��UUU�?���UU�?�?��UU�?���WU����W�������W5�?����W5���� �W5���  W5��� 0�_5����0�\�3�0 �\5�\3�\5�\=p�W5�W�_UU�W�\UUUUUU5\UUUUUU�WUUUUU�WUUU�� \UUU�� pUUUU�UUUU��_UUU?��UU�����UU�����UU� ��U� �<��U����UW�=���UWU����UU���_�UU5��WuUU �_uUU���UU�|UWU |UUU UUU�UUU5 �UUU5��_UUU�� \UUU��_UUU���WUUU��UUUU�_UUUUUUUU�WUUUUUU5\UUUUUU5��WUU�W��7\�_|5�\5��5�\53 ���W53��3\�3 ��\�0  ��\�� ���\������\������?W������U�����wUU�?���_UU����_UUU�_��WUUUUU��UUUUUUU_UUUUUUU]UUUUU�U]UUUUU]_WUUUUUW�UUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUUU�? WUUU�<\UUU? pUUU< pUUU�0pUUU?��_UUU�< \UUW�� WUU]����WU]��\U��� \U���?W�� ���U�� ��UU�U�UUUW���WUU]���_UU���?UUUU���_UUU�?�pUUU��pUUU� 0pUUUU\UUUU��W&
UUUUUUU�WUUUUUU��\UUUUUU���\UUUUUU�� \UUUUUU���WUUUUUU=�WUUUUUU� WUUUUUU<<\UUUUUU�? pUUUUU��� pUUUUU�3�3pUUUU��=��_UUUUU��\UUUU�_�� WUUUU�w���UUUUU�u��WUUUU]��?WUUU�_]���UUUU�Wu�?�UUUU�U���UUUUUU����UU�_UU���WU�WU�?�� WU�jU5��= WU?�U�s�U��V�_5pU�jU�W�_U� �U5�UUUU?��V�UUUU �UUUUUUU �jUUUUUU	��ZUUUUUU� 
hUUUUUUU��UUUUUUU) �ZUUUUUU�
 hUUUUUUU�*�ZUUUUUUU��UUUUU-UUU�|UUUUUUUUU	|UUUUUUUU�|UUUUUUUU% |UUUUUUUU	 |UUUUUUUU
�UUUUUUU���UUUUUUU%� �UUUUUUU	( �UUUUUUU	*�UUUUUUU�

�WUUUUUU�	��WUUUUU�`���WUUUUU�h���WUUUUU%X�j�WUUUUU%��Y�WUUUUU%��U�WUU�WU���U�_��\U��UUU_���\Ui�UUU_�� \UYUUUU_��WUYUUUU_�� WUUUUUU_�? WUUUUUU?<\UUUUUU} pUUUUUU��? pUUUUUU�0pUUUUUU���_UUUUUU�3 \UUUUUU��� WUUUUUU����UUUUUUU���WUUUUUU���?WUUUUUU����UUUUUUU��?�UUUUUUU���UUUUUUUU����UUUUUUU���WUUUUU�?�� WUUUUU5��= WUUUUU�s�UUUUUU�_5pUUUUUU�W�_UUUUUU5�UUUUUUUUU�UUUU.UUUUU�VUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUUU)�UUUUUUUUU� ZUUUUUUU�

�UUUUUUUU)� ZUUUUUUU�
`UUUUUUU�
  UUUUUUUU� �UUUUUUU�
�UUUUUUUU* UUUUUUUU��_UUUUUUU��WUUUUUUUU*�UUUUU�WUU�UUU��\UU�_UUU���\UU�WUUU�� \UU�UUUU��WUUUUUU�� WU�_UUUU�? WU�WUUUU�<\U�UUUUU? pUUUUUU<0p�_UUU�U��_�WUUUUW?��P�UUUUU]�< _UUUUU]����_UUUUUW����WUUUUUW��?�UUUUU�U���|UUUUU�U����UUUUU�U��WUUUUU��� WUUUUU����UUUUUUU���UUUUUUU���_UUUUUUU���pUUUUUUUU��UUUUUUUU�pUUUUUUUUU\UUUUUUUUUWUUUUUUUUU�UUUUUUUUU�UUU��WUU�??WU��? WU� ��UU���UU����UU��WU���\U�� \U��? \U��?�WUU� WUU��UUU��UUU� �UUU��W�������?�������������� �������_U��?WU����WUuU��|UuU�?�U�U��UUWUpUUUU�_UUUU�_UU��?pUU���sUU��pUU��_UU�� \UU�?�\UU�<0pUU?<��UU� �UU��UU=�UU���pUU�? \UUU��WUU� \UU��\UU��?pU��?�_U5���_}5���_�5�  ��������U�����W_�����U���
UUUUUUU�WUUUUUU��\UUUUUU���\UUUUUU�� \UUUUUU��WUUUUUU�� WUUUUU��? WUUUUU�<\UUUUU� pUUUUU�?0pUUUUUU���UUUUU�?��PUUUU]���_UUUUu����WUUUUu5��WUUUU�_��\UUUU�W�??pUUUU�U���_UUUUU���_UUU��U���_UUU��U���WUUU�UW5 �UUUUU]���WUU�_U����_UU�WUU���UU�UU����UUUU5 _� W�_UU5 \5 \�WUU�p5 \�UUUU�_��W.UUU�|UUUUUUUUU	|UUUUUUUU�|UUUUUUUU% |UUUUUUUU	 |UUUUUUUU
�UUUUUUU���UUUUUUU%� �UUUUUUU	( �UUUUUUU	*�UUUUUUU�

�WUUUUUU�	��WUUUUU�`���WUUUUU�h���WUUUUU%X�j�WUUUUU%��Y�WUUUUU%��U�WUU�WU���U�_��\U��UUU_���\Ui�UUU_�� \UYUUUU_��WUYUUUU_�� WUUUUUU_�? WUUUUUU?<\UUUUUU} pUUUUUU��? pUUUUUU�0pUUUUUU���_UUUUUU�3 \UUUUUU��� WUUUUUU����UUUUUUU��? WUUUUU����\UUUUUU����sUUUUUU�����WUUUUU����\UUUU�U5  \UUUU�U���<\UUUU�U����WUUUUU����_UUUUUU}��UUUUUU����UUUUUU5 _� WUUUUU5 \5 \UUUUU�p5 \UUUUUU�_��W.UUUU�jUUUUUUUUU��ZUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUUU)�UUUUUUUUU�ZUUUUUUUU�
�UUUUUUUU�� ZUUUUUUU�
�UUUUUUUU*� VUUUUUU��  PUUUUUUU�
 _UUUUUUU� �_UUUUUUU��WUUUUUUU�
�UUUUUUUU) UUUU�_UU��_UU��?pUU��WUU���sUUU�UUU��pUUUUUU �_UU�_UUU��\UU�WUUU�� \UU�UUUU�<�pUUUUUU?< �U�_UUUU� �U�WUUUU���U�UUUUU?�UUUUUU�� p�_UUUUU��\�WUUUUU���W�UUUUUU�� �UUUUUW��?0pUUUUU]���3pUUUUU]����pUUUUUu���_UUUUUu���\UUUUU��  \UUUUUU����WUUUUUU���UUUUUUU����UUUUUUU���WUUUUU� |�\UUUUU� p� pUUUUUU�� pUUUUUU�U�_UUUUU.UUU�|UUUUUUUUU	|UUUUUUUU�|UUUUUUUU% |UUUUUUUU	 |UUUUUUUU
�UUUUUUU���UUUUUUU%� �UUUUUUU	( �UUUUUUU	*�UUUUUUU�

�WUUUUUU�	��WUUUUU�`���WUUUUU�h���WUUUUU%X�j�WUUUUU%��Y�WUUUUU%��U�WUU�WU���U�_��\U��UUU_���\Ui�UUU_�� \UYUUUU_��WUYUUUU_�� WUUUUUU_�? WUUUUUU?<\UUUUUU} pUUUUUU��? pUUUUUU�0pUUUUUU���_UUUUUU�3 \UUUUUU��� WUUUUUU����UUUUUUU��? WUUUUU����\UUUUUU����sUUUUUU�����WUUUUU����\UUUU�U5  \UUUU�U���<\UUUU�U����WUUUUU����_UUUUUU}��UUUUUU����UUUUUU5 _� WUUUUU5 \5 \UUUUU�p5 \UUUUUU�_��W0UUUUU�jUUUUUUUUU��ZUUUUUUUU�
`UUUUUUUUU��VUUUUUUUU	
hUUUUUUUU%��UUUUUUUU��ZUUUUUUU�
`UUUUUUU�
(�UUUUUUUU)  VUUUUUUU
  TUUUUUU� �_UUUUUU�� �_UUUUUUU*��UUUUUUU�
�_UUUUUUUU��UUUUUUUUU�_UUUUUUUU��UUUUUUUU��_UUUUUU���UUUUUUU�?�_UUUUUUU���WUUUUUUU��WUUUUUUU?� WUUUUUU�3� WUUUUUU��0<\UUUUUU��? pUUUUU�?<� pUUUUU��?�0pUUUU�����_UUUU�WW�? \UUUUUU]�? WUUUUUU]���UUUUUUUW�� WUUUUUUW��\UUUUU�U���sUUUUU�U����WUUUUUW���\UUUUU]7  \UUUUU����\UUUUUU����WUUUUU����UUUUUU5���UUUUUU�__UUUUUU�� \UUUUUU�� pUUUUUU� W�UUUUUUU�U�UUUUUUU�WUU��\UU���\UU�� \UU��WUU�� WU��? WU�?<\_� �p�? 0���<�����pU??��_W����W]����Uu���Uu���_U]���_UW����UW���W]5  W����WU����U����U5���U���_U�5 WUp5 \U5�� pU�U�_U 	UU  PUUUUU��CUUUUU   @UUUU���OUUU     @UU�?��OU ��00 @U����03�TU ��00 @UU�?��OUU     @UU�����?PU      TU�����?UU       TU�������T        T������PU       UUU����?UUU      UUU�����@UUU      TUUU�����TUUU     TUUU���CUUUUU    PUUUU���SUUUU   PUUUUU��PUUUUUU  UUUUUUUUPUUUU 	UUU  PUUUUU���PUUUU   @UUUU����UUU     @UU�����OUU  PU��3��SU  PU�����OUU     @UU��?��SUU      TUU�����T       T����3�CU        U��?���?UU       UU�?��?TUUU      UUU��?�?UU      UU����CUUU     UUUUU��??UUUU    UUUU����PUUUU   TUUUUU?UUUUUUU  UUUUUUUUUUU UUU   UUUU��?UUUU   TUUU��?�PUU     @UU�?�OUU ��00 @U���03�O ��00 @�?��T      TU�����?UU     @U������O      @�?��?�?T      PU �����SU     PU�����CUU     PU�����SU     PU�?�?TUU    PUUU���SUUU   PUUU�?�UUUU  @UUUUU �PUUUUU PUUUUUUPUUU UU@UUU  TUU��PUU  @UU�?�U    T���T00P�33��S00@����O    @�����O    @�����O    @�����O    @�����C    P����P    T���?TU    UU���OUU  @UU��PUU  TUU�<TUUU  UUUU�CUUUUPUU0UUU)_UUUUUUUUUU_UUUUUUUUU� _UUUUUUUUU	 _UUUUUUUUU _UUUUUUUU��_UUUUUUUU%� _UUUUUUUU	( UUUUUUUU
|UUUUUUUU�
|UUUUUUU���|UU�UUUU�h� |UU]UUUU%��(~�_�_UUU%��+��5�U]U	����  � _UU�&j��  < \�U�%j�    \UU��e��    |]UbeU��  �?�uUZeuU� ����uUVUU��������UVUU���� �UUU� �3 �? �UUUU���0 |UUUU���0 \UUUU����� pUUUU����  pUUUuU�?� �UUU�_����UUU5����� �]UU� ��?� �WUUU ��0  WUUU ���  \UUU �0  \UUU<���  \UUu50<��? \UU��0<���? WUU�<0����� WUU� � �� WUUU0�����WUUU0��?<�UUUU0���� �WUUU����� WUUU5 ��� WUUU� � 0�UUUU�� ��UUUUU< �pUUUUU5�� �?\U0UUUUU��UUUUUUUUU�jUUUUUUUUU*�UUUUUUUUU�ZUUUUUUUU%(�UUUUUUUU��VUUUUUUU�
hUUUUUUUU
(�UUUUUUU�*� VUUUUUUU�  XUUUUU]U)  PUUUUU��
  �UU�__��UU�?|5� �W��? � /�UU     ��WUU5     �UUU�    �WUUUU5  ��?WUU�U���\UU5_���? pUU5� �?� pUU�  ��? \UU�  �  WUUU �  WUUU5����0 \UUU�� � \UUU����� \UU}����� �UU�� ?�?�uUU�<� 0��UU 0��  �UU= 0��� �UU5 �� �UU� ��?0 �UUU���� pUUU����pUUU���30pUU�0�  <0\UU7 ����30\UU  ����\UU5  ���� \UU� ����� pUU� 0�?< pUUU0�0 pUUU=0 � _UUU�� �UUUUU���@UUU&	U]UUUUUUUUuU�UUUU��_U�WUUUU�W�UU�U |5�WUUW= � WU�\5   |U�p5    pU���  ��UU�5�� WU��� WU ��  \U �� \U ��  \]��?  \u=�?<p��� �0p���? 0�p���<�p<����0p5  ??��\5 ����\� ���� p� 0���? pW0��� pu��� p����� p�����0  �5 �����5  ���� �5 ����? ��0���? �U��� \U=�0  _U500 �UU�0�� 0�UUU�? �U}}����z�^�WUU                                                                                                                                                                                                                                                                                                                     �(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �
                                      ��                                     ��U�
                                   �jUU*                                   �ZU�*                                   �ZU��                                   �VU��                                   �UUU�                                   �UUU�                                U  �UUU�                             TUAU�UUU�
                            T   U�UUUZ
                                 �VU�Z	            �*             @     �VU�V%           �j��            @  UU  PU�V�           �ZiU&           @ @   ZUU�U�           �ZiU�           @ P@ �ZUUeU�          �ZiU�           @ @�jUUUU�          �ViU�              P�ZUUUU�          �ViU�           @  PU�VUUUU�          �ZYU�
            UUUV�VUUUU�          �ZYU�
              eV�UUUUV�          �VUU�
              hU�UUUUZ�          �VUU�
              jUiUUUUZ�          �VUU�
              jUZUUUU^U.          �VUU�* �            jUZUUUU^U.          �VUUU*�j� U         jUZUUUU]U:         ��VUUU)�V�R U        jUZUUUU]U:         U�VUUU)�UU         jUZUUUUUU:       @U �V TU)�VU-         jUZUUUUUU:         �  PU)�ZU�P@       ZUZUUUUeU:      @     PUU��ZU�       ZYZUUUUi�:      @    UUU��VU        ZYVUUUU��>          @UUU�hUU  @      �ZYVUUUUj�>       P  XUUU�ZU @P      �ZYUUUUUj�6        UUUUUUU�jU    P      �VYUUUUUj�         �j�UUU
            �VZUUUUUi��        �ZiUUU�*  T       �VVUUUUU��ZP       �ZYUUU�j�@�@     ���VUUUUU��Z        �VYUUU�j�V�UU      �i�VUU            �VVUUU�j�V�       �e�V�UU%            �VVUU��j�V�       ���U�UUU�
   @       ��VUU��j�V�       ��UU�UUU��  @       ��VU�j�j�V�       ��UU�UUUU�  P       ��VU�U�j�U�       �jUUiUUUU�ZU        ��ZU�U�j���       �jUUjUUUU���U        ��ZUiU�j�e�
       �jU�jUUUUU��         ��VUYU�j�[�*       �jU�jUUUUUU�         ��UUUU�j�Z�*       �jU�jUUUUUU�         ��UUUU�j�V�*       �jU�jUUUUUU�         ��UUUU���UU*       �jU�ZUUUUUU�         �jUUUUU��UU*       �fU�ZUUUUUU�         �jUUUUU�VUU*       �fU�ZUUUUUU�         �jUUUUU�VUU)       �eU�VUUUUUU�        �ZUUUUU�ZUU)       �UU�UUUUUUU�        �ZUUUUU�ZUU)      ��UUiUUUUUUU�        �ZUUUUU�ZUU�      ��UUiUUUUUUU�
       ��ZUUUUU�ZUU�     ��UUYUUUUUUU�
       ��ZVUUUU�ZUU�     �ZUUYUUUUUUU�
       ���VUUUU�ZUU�     �ZUUYUUUUUUU�
       ���VUUUU�ZUU�     �ZUUYUUUUUUU�
       ���VUUUU�ZUU�     �ZUUYUUUUUUU�
       ���UUUUU�ZUU�
     �VUUjUUUUUUU�
       ���UUUUU�ZUUU*     �VUUjUUUUUUU�)       �V�VUUUUUjUUU*     �VUUZUUUUUUU�)       �V�ZUUUUU�UUU)    ��UUUZUUUUUUU�)       �V�ZUUUUU�VUU%    �ZUUUZUUUUUUU��       �V�ZUUUUU�VUU�    �jUUUZUUUUUUUU�       �Z�ZUUUUU�VUU�   ���UU�ZUUUUUUUU�
     ��j�VUUUUU�VUU�   ���UU�VUUUVUVUU�*     ��Z�VUUUUU�VUU�  ���jU�VUU�ZUiUU���   ���V�UUUUUU�VUU�� �������VU��U������������V�VUUUUU�jUUU���                   ��������jUUU���Z�����UUUUUUUU�WUUUUUUU��\UUUUUUU���\UUUUUUU�� \UUUUUUU��WUUUUUUU�� WUUUUUUU�? WUUUUUUU�<<\UUUUUUU?< pUUUUUUU� pUUUUUUU�3pUUUUUUU���_UUUUU�U�\UUUUUU�� WUUUUU����UUUUU��W�� WUUU��W]?�?\UU��WU]���WU��WUU]���WU�WUUUu���UUUUUUu����UUUUUU�5  �UUUUUU����?_UUUUU����pUUUUU��?�?�UUUUU�0 �UUUUU��UUUUU�  ��UUUUU�    |UUUUUU����WUUUU�UUUUUUUU��WUUUUUUU�??WUUU��UU�? WUU���UU��UU���UUU�?�U���UUU������UUUU�?���UUUUU���UUUUUU���\UUUUU�����\UUUUUU����WUUUUU�}�� WUUUUUu�??�UUUUUUu�?�UUUUUU]�?��UUUUUU]���WUUUUU]����UUUUUUu����UUUUUU�U���UUUUUUU �_UUUUUU���?pUUUUUU�����WUUUUU����?\UUUU�0����pUUUU5�� sUUUU5�� <�pUUUU� ? �pUUUUU    _UUUUU�����UUUUUUUUU�UUU��WUU�??WU��? WU� ��UU��?�UU���UU��WU�� \U��? \U��� \u���<W����<W�U??�Uu���Uu��3�U]���W]����Uu����Uu����U�U WU���W�����\5����p������� �<0 ������    |U����W$	UU��UUUUUU �WUUUUU3  \UUUU�<  pUUUU5? 0�UUUU5  ��UUUU ��UUUU ��UUU� � ��UUU5 ��UUU�� ��UUUU?�0 \UUUU�0 WUUU�W�?�UUUU�U��sUUUUUU��_UUUUUU��WUUUUU� �UUUUUU5 \UUUUUU _UUUUUU WUUU}UU?�U�U�UU�U�W�W��_��_�_��_��_�_��W�?��_��W������ W������ \�����Up5��pU�\� 7pU?�W��?\U��W��?WU���UU��UU�?|UU��UUU�WUU�U$	UUU��_UUUUU� �WUUU�   �_UUU? ��UU�� 0�?WU� ��?\U  p�\U � p�pU5� \� pU�� �W� pUU?�WU�pUUpUU�\UU7\U��?WU��W���UUuUU� �UU]U�� �_UUUU=��UUUU��_UUUU5 ��UUUUU �_UUUUU |UUUUUU?�WUUUUU��|UUUUUU��WUUUUUU��UU�UUU5�UU�WUU5�UU _UU5 W� �UU5�W� ��UU��_���UU������?_�U���p�U� �_U�U= �WU�U�\UU��_UU�WUUU�W$UUUUUU��WUUUUUUUU� \UUUUUUUU�? pUUUUUUUU�� �UUUUUUUU�� WUUUUUU��� \UUUUUU���? \UUUUUU5�� pUUUUUU5�_� pUUUUUU WU|UUUUU� �UU�UUU�� �U��UUU=   pU��UU�3 pU��_UU?  \U�_UU 3 �W� �WUU   |U5 �UUU � \U pUUU=� WU \UUU�< �U� WUUUU�UU��UUUUU_UU��pUUUUU�UUU��_UUUU�UUUU��WUUUUuUUU���UUUUU]UUU��UU�WUUUUU� \U� |UUUUU� \U��UUUUU� pU��WUUUU� ����WUUUUU�?���_UUUUU��W�UUUUU��pUUUUUUU��\UU}UUUUUU?�WUU}UUUUUU��UUUu$	UUUUUUUUUUUUUUU�_UUUUUUU��UUUUUU���WUUUUU��\UUUUU �pUUUU� ?pUUUU��?�UUUU�?|�UUUU�?W5�UUUU��U5�UUU���U5�UUU U��U��  \��U5   W��U3 ����_�  ?? �W? 3 � �U   � |U �� _U ?���UU=� ���_UU��UUUUUU�_UUUUUU��WUUUUU���WUU�_Uu�WU��U] WU��WU \U�? _U |U�?�_U5 �����U� ��WU�UU��UU�UU��pUU�UU��\UU�UUU��WUU�$	UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUU� _UUUUUU �UUUUUU �WUUUU�  �_UUUU� ��_UUUU�?��pUUUU��U?pUUUU��U5�UUUU��U5�UUU�|��UU�� ���UU�� 0�?pUU�? 0�?\UU ��WU��  ��WUU=   UUUU3 �UUUU�  pUUUU= 3pUUUU  \UUUU � W�_UU ?�U5�WU�� �_ UU��� ��WU7���_�_��W��U�uUU�\UU]UUU�WUU�$	U�_�W��UUU�| _UU ��  �UU�� 0 �WUs� � �\U]5  ���pUU�  ��?pUU�? pU?�UU� \U�U� �WU�U_?_UU?��U��UU�?psUpUU��p\U5\U� �_WU�W� �WUUUU� |UUUU��? _UUUU�?�UUUU� ��\UUUU5 ��WUUUU �_UUUUU? �UUUUU���WUUUUU��UUUUUU��_�UUUU�W5�WUUU�W _UUU�U�UUU � ��UUU � ��UUU5 ��?_�U5 ���p�U� �U�UU�U�UU=�_U5�_UU��WU��W$	U}UUUU�UUU�_�U� U� � � �U�0 <<  �W���   �\UW   ��pUU5  ��?pUU�  \U?�U��  WU�U�� �UU��5 |UU?�UW�WU�?p�U\UU��pu��WU��_U5pU� �WU�_U� �UUUU��? UUUU�?�WUUU���_UUUU5 �UUUUU �WUUUUU? |UUUUU��WUUUUU���UUUUUU��UUUUUU��_UU�_UU�WU��UU WU��WU \U�?�_U \U�?�_U5 �����U� ��_U�UU��UU�UU��pUU�UU��\UU�UUU��WUU�$UUUUUU��WUUUUUUUUU \UUUUUUUU�? pUUUUUUUU�� �UUUUUUUU�� WUUUUUU��� \UUUUUU���? \UU�WUU5��� pUU|�_�� pUU�p _U|UU� ��  WU�UUs� �U��UUs pU��UU]5   \U��_UUU�   WU�WUUUU �U� �WUUUU pU5 �UUUUU pU pUUUU� \U \UUUUW W� WUUU�U�U��UUUUuUpU��pUUUU_UpU��_UUUUU� \U��WUUUU�< WU��UUUUU��U��UU�WU5 _U� \U� |U��UU� \U��UU}UU� pU��WUUUU� ����WUUUUU�?���_UUUUU��U�UUUUU��pUUUUUUU��\UU}UUUUUU?�WUU}UUUUUU��UUUuUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUU��_UUUUUUUUUUUUUUUUU�UUUUUUUUUU�UUUU� ��UUUUUUUUU��_UUU5 ��WUUUUUUU�   �WUU= ��\UUUUUUU? �_UU� �?pUUUUUU�� 0�U�� ��UUUUUU� 0��U���U WUU�_U  0��W��_U \U��U � ���\��WU5 |U��W5� \�?���UU� �U�?�_�� �W�?  UUU��W�?�_U?�WU�  \UUU������UpUU�  WUUU���_UU7\UUU �UUUU�� �UU���WUUU5 pUUUUU pUU�uUUUUU�\UUUUU= \UU�]UUUUUU�WUUUUU��WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_�W��UUUUUUUUUUUUUUU�| _UUUUUUUUUUUUUU ��  �UUUUUUUUUUUUUU�� 0 �WUUUUUUUUUUUUUs� � �_UUUUUUUUUUUUU]5  ���UUUUUUUUUUUUUU�  ���sUUUUUUUUUUUUUU�? pU��UUUUUUUUUUUUUU� \U�UUUUUUUUUUUUU� �W� �UUUUUUUUUUUUU_?_U� �UUUUUUUUUUUU�U��UU5 pU��WUUUUUUUUwUpUU= \U��UUUUUUUU]U5\UU� W� ��UUU�WUUUWU�WU���U ��WU� |UUUUUUUU��U? ��_U5 �UUUUUUUU��_�� ��pU �WUUUUUUU��W����?p� �_UUUUUUU��_�����?��U]UUUUU�����_U ��|��U_UUUUU�� �WU= ��W= �_UUUUU��  �UU5  �U5 �WUUUUU�  \UU� U���WUUUUUU �WUUU=�UUU��UUUUUUU��UUUU�UUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUU�UUUUUUUUUUUUUU���U=�_UUUUUUUUUUUUU5 <�� |UUUUUUUUUUUUU5   �UUUUUUUUUUUUU5��<  �?WUUUUUUUUUUUU�U   �?\UUUUUUUUUUUUUU  ��\UUUUUUUUUUUUUU5  W�pUUUUUUUUUUUUU�? �UUpUUUUUUUUUUUUU}5 pUUpUU��UUUUUUUU�_ _U� pU���UUUUUUU�U�UU� \U���WUUUUUUu� WUU�\�  ��_UUUUUU]7�UU��W  ��UU�_UUU\UU���U? ����U��UUU�WUU��_��_��W� WUUUUUU��W���UU? \�? _UUUUUU��_��UU ��?�UUUUUU�����_UU5 ����UUUUUU�� �WUU�  �_U�UUUUUU��  �UUUU �UU�UUUUUU�  \UUUU= pUU�WUUUUUU �WUUUU�\UU�WUUUUUU��UUUUUU�WUUU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUU�UUUUUUUUUUUUUU5��U=�_UUUUUUUUUUUUU �� |UUUUUUUUUUUUU   �UUUUUUUUUUUUU��  �?WUUUUUUUUUUUU�500  �?\UUUUUUUUUUUUu�   ��\UUUUUUUUUUUUUU  W�pUUUUUUUUUUUUUU �U�pUU�UUUUUUUUUU pU�pUU�WUUUUUUUUU pU5 pU� �UUUUUUUU� \U= \U ��WUUUUUUU] \U� \�  ��_U�WUUU}W W��W� ����UUU�U�U���U������5��UUU}U�U��_���_��?��WUUU]pU��W���WU� ��_UUU� \U��_��UU� ��pU]U3�WU��� �_UU5  |?�U_� |UU��  WUU�  W �_UWUU��  �UUUU�U5 �WU�UUU�  \UUUU=|U���WUUUUUU �WUUUU�WUU��UUUUUUU��UUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUUUU5��UUUUUUUUUUUUUUUU ��_UUUUUUUUUUUUUU  �UUUUUUUUUUUUUU��  UUUUUUUUUUUUU�5   �_UUUUUUUUUUUUu��  �UUUUUUUUUUUUUU  ��UUUUUUUUUUUUUU � �?WUUUUUUUUUUUUU p��?\UUUUUUUUUUUUU p��\UUUUUUUUUUUU� \U� pUUUUUUUUUUUU] \U= pUUUUUUUUUUU}W WU pUU��UUUUUUU�U�UU \U���UUUUUU}U�UU= pU���WUUUUUU]pUU�\U ��_UUUUUU� \U��?W�  ��UU�_UU3�WU���U� ���U��U� |UU���U�?���W� WUWUU��U��_U? \�? _U�UUU������WU ��?�UUUUU�����UU5 ����UUUUU��? �UU�  �_U�UUUUU�� �_UUU �UU�UUUUUU?  �UUUU= pUU�UUUUUU�  |UUUU�\UU�UUUUUUU��WUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUU�?�_UUUUUUUUUUUUUUUUU?  |UUUUUUUUUUUUUUUU�   �UUUUUUUUUUUUUU��  �?WUUUUUUUUUUUUU=    �?\UUUUUUUUUUUU�3 ��\UUUUUUUUUUUU?  W�pUUUUUUUUUUUU 3 �U�pUU�UUUUUUUU   |U�pUU�WUUUUUUU � \U5 pU� �UUUUUUU=� WU= \U ��WUUUUUU�< �UU� \�  ��_U�WUUUU�UU��W� ����UUUU_UU���U������5��UUUU�UUU��_�����?��WUU�UUUU��W���WU� ��_UUuUUUU��_��UU� ��pU]]UUUU��� �_UU5  |?�U_UUUUU��  WUU�  W �_UUUUU��  �UUUU�U5 �WUUUUU�  \UUUU=|U���WUUUUUU �WUUUU�WUU��UUUUUUU��UUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUUU��_UUUUUUUUUUUUUUUUUU�UUUUUUUUUUU�UUUU� ��UUUUUUUUUU��_UUU5 ��WUUUUUUUU�   �WUU= ��\UUUUUUUU?  �_UU� �?pUUUUUUU�� 0�U�� ��UUUUUUU  0��U���U WUU�_UU�0��W��_U \U��UU � ���\��WU5 |U��WU5 < \�?���UU� �U�?�_U���W�?  UUU��W�?�_UU?�WU�  \UUU������UUpUU�  WUUU���_UUU7\UUU �UUUU�� �UU�U��WUUU5 pUUUUU pUU�UuUUUUU�\UUUUU= \UU�U]UUUUUU�WUUUUU��WUUUU.UUUUUU�_�W��UUUUUUUU�| _UUUUUUU ��  �UUUUUUU�� 0 �WUUUUUUs� � �\UUUUUU]5  ���pUUUUUUU�  ��?pUUUUU�W�? p�?�UUU��\_� \U�UUU����U�WU�UUU�� \_U��UUU��W��UU�pUUU�? WpUU��pUU��3W5\U���_UU�?\�WU��WUU�3pUU�  UUU�? pU�� _UUU�� pU���UUUUU��_����\UUUUU=? ����WUUUUU� 7 ��_UUUUUU���  |UUUUUU�� ���WUUUUUU�����sUUUUUUU�? �?�_UUUUUU�� �� UUUUUU�� �� |UUUUUU��  �� |UUUUUU��  �� _UUUUUUU�? �?��UUUUUU������ WUUUUU5�� �? _UUWUU�� �� |U�WUU��  ��|U�UUU��  ��U�UUU?�� ���_�UU���� ���W5UU�? �������\UU� ���� �? WUU� ��?  ���UUU� ��  ��pUUU�? ��  ��\UUUU� ��  ��WUUUU�?��?  �UUUUU���� ��UUUUUUU������_UUUUU/UUUUUU_UUUUUUUUUUU���U�WUUUUUU5 <�� |UUUUUU5  �WUUUUU5��< �_UUUUU�U  �_UUUUU�U  ��UUUU�U5  ��sUUU���U? �W��UU�����5 pU=�UU���_ _U�UU5 �U�U�pUU��p� _U�pUU���s5�UU�?\UU�� �\U���WUU�� �WU=��UUU=� WU��UU�7��WU? �_UU��U�� �WUU������|UUU� p=��?WUUU����_���UUUUU�? � ��WUUUUU��?��_UUUUUU�����UUUUUU����?�UUUUUU��  �� WUUUUU��  �� WUUUUU�?  �� WUUUUU��  �?�UUUUUU�� �_UUUUU�����pUUUUU�� ��UUUU� ��  �? WUUU� �?  �� WUUU� ��  �� �_UU��� ���5pUU���� �?|�UU� �������WU�  �� � �_U� ���  ���_U� ��?  �sUU�? ��  �U}U�� ��?  �_U�U����� ��WUUUU�����_UUUUUU������UUUUU5UUUUUU�_UUUUUUUUUUUU5��UUUUUUUUUU �UUUUUUUUUU WUUUUUUUUU��\UUUUUUUUU�500pUUUUUUUUUu�  �UUUUUUUUUUU  _UUUUUUUUUU  �UUUUUUUUUU  �_UUUUUUUUU  �UUUUUUUU� 0��UUUUUUUU] ��?WUUUUUU}W ��\UUUUU��U W�pUUU��U�UUpUUU�??W]pUU�UU��? W� \U��UU� ��U3�WU��UU���� |UU�?pUU���UWUU��pUU��0W�UU���_UU��\UU���WUU�� \U�� ��UUU��?�_��� �UU�U�? W��? �WUUW�����?�_UUU_�� �?UUUU����� ��UUUUU���  �?�_UUUUU�����?��UUUUUUU��� _UUUUUU��� ��\UUUUUU5�? ��\UUUUUU5�? ��\UUUUUU5�� ���WUUUUUU����?�UUUUUU5 ������UUUUUU �� ��WUUUUU ��  ��_UUWUU �?  ��U�WUU �   �U�UU���?  ��U�UU�����  ��_�UU��?�����W5UU��  ��  �\UU�� ��?  < WUU�� ��  ��UUU�� ��  �pUUU��? ��?  �\UUUU�� ���  �WUUUU�� ��?�UUUUUU�������WUUUU�_�z������z�_                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �(                                       DUTQEUT          @UTUQQQEUT             ����     @  @   @               @    ����*       @       @    ��     @    ������    @  @   @   @          @   ��  �*   @  @   @   @     TUUEU  �*TeU���  EQUQUEUA @       ��BUeU�*               ��@         �*TUeUU��"             @ XU@      ��BUUeUU��            @  XU       ��TUUeUU�*            @ XUPEUTEE �*UUAeUU�* QUUPUAQQEEUXU    @    �JUU eTU��  @  @        XU   @    �JUUAeUU��    @   @         XU   @    �RUUUeUUU�  @           XU   @    �VUUUeUUU�   @           XUUTUUA  �RA e@� UUUUTUU@APUU ��       �V �*e�J�          @            �VA�*e�J�         @             �RU�*e�JU�         @           �VUJe�RU�              PEUUEQ  �VUJe�RU�PUUUQUUATEEQPUUD  @      �RU�*e�JU�  @  E      @     @       �VU e@U�  @  D            @       �VAUUeUU�  @  @      @            �R UUeUU�  @       @    DEUUUEUE �VAUUeUU�UUUUE TU@UEU     @@   �VUUPeTU�                  @@   �RU@ePU�      @          @@    �VUUPeTU�        @       ��         �VUUUeUUU�                            �����������                  ����������BUUUUUUU�������������������
          �@UUUUUUU(                  ��          @UUUUU                   XUUUUUUUUUUUUUUUUUUUUUUUUUUUU        XU            UUUUU          @        XU            UUUUU          @        XU            UUUUU          @        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        ��UUUUUUUUUUUUUUUUUUUUUUUUUUUU@         UUUUUUUUUUUUUUUUUUUUUUUUUUUU@         UUUUUUUUUUUUUUUUUUUUUUUUUUUU@         UUUUUUUUUUUUUUUUUUUUUUUUUUUU@         UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ ��*  ��
 UUUUUUUUUUUUUUUUUUUUUUUUUUUU@     �   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@     �   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@  ����   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@  `UU�   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@  `UU�   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ �jUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUU@  `UU�   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ �*`UU�   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@  ����   UUUUUUUUUUUUUUUUUUUUUUUUUUUU@         UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ ��������UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ �*       UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%       UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%       UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%       UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ �*                        PUUUUUUUUUU@                          PUUUUUUUUUU@ �*  ����                 PUUUUUUUUUU@     �   UUUUUUUUUUUUUUUUPUUUUUUUUUU@     �   UUUUUUUUUUUUUUUUPUUUUUUUUUU@  ����                   PUUUUUUUUUU@  `UU�                   PUUUUUUUUUU@  `UU�                   PUUUUUUUUUU@ ��jUU��
                 PUUUUUUUUUU@  `UU�    ����  ���
   PUUUUUUUUUU@  `UU�    �          PUUUUUUUUUU@  ����    �          PUUUUUUUUUU@        ���   ���  ��
 PUUUUUUUUUU@       ��UU�   VUU  XU	 PUUUUUUUUUU@        UU�   VUU  XU	 PUUUUUUUUUU@ UTU UU����VUU���ZU	 PUUUUUUUUUU@ @  @   UU�   VUU  XU	 PUUUUUUUUUU@    @  ��UU�   VUU  ��
 PUUUUUUUUUU@ @  @  XU���   ���  �  PUUUUUUUUUU@ @  @  XU            �  PUUUUUUUUUU@ BEQUXU**�����������  PUUUUUUUUUU@       XU            �  PUUUUUUUUUU@       XU            �  PUUUUUUUUUU@       XU            �  PUUUUUUUUUU@       XU            �  PUUUUUUUUUU@ F@UETXU            �  PUUUUUUUUUU@     ��            �  PUUUUUUUUUU@                   �  PUUUUUUUUUU@                   �  PUUUUUUUUUU@                   �  PUUUUUUUUUU@ PUUA             ��
 PUUUUUUUUUU@    P               �  PUUUUUUUUUU@   @               �  PUUUUUUUUUU@   @               �  PUUUUUUUUUU@   @               ��
 PUUUUUUUUUU@ TQU             �U	 PUUUUUUUUUU@                  �U	 PUUUUUUUUUU@                  �U	 PUUUUUUUUUU@                  �U	 PUUUUUUUUUU@     ��            �U	 PUUUUUUUUUU@ BPUA              �U	 PUUUUUUUUUU@                   �U	 PUUUUUUUUUU@                  �U	 PUUUUUUUUUU@      ��            ��
 PUUUUUUUUUU@       XU            �  PUUUUUUUUUU@       XU            �  PUUUUUUUUUU@ �������ZU            �  PUUUUUUUUUU@        XU            �  PUUUUUUUUUU@        XU            �  PUUUUUUUUUU@        XU            �  PUUUUUUUUUU@        XU            �  PUUUUUUUUUU@        XU            �  PUUUUUUUUUU@        ��            �  PUUUUUUUUUU@                     �  PUUUUUUUUUU@UUUUUUU              �  PUUUUUUUUUU@UUUUUUU              �  PUUUUUUUUUU                      ��
 PUUUUUUUUUU                ����� �  PUUUUUUUUUU                (   ��  PUUUUUUUUUUUUUUUUU        ZTU
�  PUUUUUUUUUUUUUUUUU        �T%UI	��
 PUUUUUUUUUUUUUUUUU        �P%T		�U	 PUUUUUUUUUUUUUUUUU        �P%T
	�U	 PUUUUUUUUUUUUUUUUU        �Q)T
	�U	 PUUUUUUUUUUUUUUUUU        �Pi�
	�U	 PUUUUUUUUUUUUUUUUU ��      �Q*�	�U	 PUUUUUUUUUUUUUUUUU        �Qj�
	�U	 PUUUUUUUUUUUUUUUUU        �Qj�	�U	 PUUUUUUUUUUUUUUUUU        �Qj�	�U	 PUUUUUUUUUUUUUUUUU ��      �Qj�	��
 PUUUUUUUUUUUUUUUUU XU      �Qj�	�  PUUUUUUUUUUUUUUUUU XU      �Qj�	�  PUUUUUUUUUUUUUUUUU XU      �Qj�	�  PUUUUUUUUUUUUUUUUU XU      �Qj�	�  PUUUUUUUUUUUUUUUUU XU      �Qj�	�  PUUUUUUUUUUUUUUUUU XU      �Qj�	�  PUUUUUUUUUUUUUUUUU XU      �Qj�
�  PUUUUUUUUUUUUUUUUU XU      �Qj���  PUUUUUUUUUU         ��      �Qj�� �  PUUUUUUUUUU                ����* �  PUUUUUUUUUU          �(   P@UUUUUUUUUU@      @    ����*  @   P@UUUUUUUUUU@          ������      P@UUUUUUUUUU@         ��  �* @   P@UUUUUUUUUU@ QTUQTUE  �*TeU��� P   P@UUUUUUUUUU@   @      ��BUeU�*    P@UUUUUUUUUU@           �*TUeUU��" �* P@UUUUUUUUUU@ @       ��BUUeUU��    P@UUUUUUUUUU@ @       ��TUUeUU�*   P@UUUUUUUUUU@ BUQ @ �*UUAeUU�*   P@UUUUUUUUUU@  PU@  �JUU eTU���* P@UUUUUUUUUU@         �JUUAeUU�� U% P@UUUUUUUUUU@       @  �RUUUeUUU�U% P@UUUUUUUUUU@     @  �VUUUeUUU� U% P@UUUUUUUUUU@ TUA P �RA e@�U% P@UUUUUUUUUU@    @Q  �V �*e�J�U% P@UUUUUUUUUU@  @      �VA�*e�J�U% P@UUUUUUUUUU@  @      �RU�*e�JU�U% P@UUUUUUUUUU@  @  @    �VUJe�RU�U% P@UUUUUUUUUU@  ETUU �VUJe�RU��* P@UUUUUUUUUU@     @  �RU�*e�JU�   P@UUUUUUUUUU@         �VU e@U�   P@UUUUUUUUUU@          �VAUUeUU�   P@UUUUUUUUUU@         �R UUeUU�   P@UUUUUUUUUU@ QQPU Q �VAUUeUU�   P@UUUUUUUUUU@  @     �VUUPeTU�   P@UUUUUUUUUU@  @      �RU@ePU�   P@UUUUUUUUUU@         �VUUPeTU�   P@UUUUUUUUUU@          �VUUUeUUU�    P@UUUUUUUUUU@          �����������   P@UUUUUUUUUU@ �����������BUUUUU��   P@UUUUUUUUUU@           �@UUUUU(    P@UUUUUUUUUU@            @UUUUU  �* P@UUUUUUUUUU@            @UUUUU     P@UUUUUUUUUU@            @UUUUU     P@UUUUUUUUUU@            @UUUUU     P@UUUUUUUUUU@            @UUUUU  �* P@UUUUUUUUUU@            @UUUUU  U% P@UUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUU                UUUUU   U% P@UUUUUUUUUU                UUUUU   U% P@UUUUUUUUUU                UUUUU   U% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�* P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�* P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�* P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�* P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUU          P@UUUUUUUUUUUUUUUUUUUUUUUUUUU          P@UUUUUUUUUUUUUUUUUUUUUUUUUUU          P@UUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUU         P                 @UUUUUUUUUU         P                 @UUUUUUUUUU         P                 @UUUUUUUUUU      �* PUUUUUUUUUUUUUUUUU@UUUUUUUUUU ����   PUUUUUUUUUUUUUUUUU@UUUUUUUUUU                         P@UUUUUUUUUU                         P@UUUUUUUUUU     ��*                  P@UUUUUUUUUU     VU%                  P@UUUUUUUUUU ����VU%����  ���*  ���* P@UUUUUUUUUU     VU%�          �    P@UUUUUUUUUU     VU%�          �    P@UUUUUUUUUU     VU��   ���
  ����    P@UUUUUUUUUU �� �UU�   VUU	  `UU�    P@UUUUUUUUUU `U  UU�   VUU	  `UU�    P@UUUUUUUUUU `U���UU����VUU���jUU��  P@UUUUUUUUUU `U  UU�   VUU	  `UU�   P@UUUUUUUUUU `U  ZU�   VUU	  `UU�   P@UUUUUUUUUU `U  ���   ���
  ����   P@UUUUUUUUUU `U                   �* P@UUUUUUUUUU ��  �����������������  P@UUUUUUUUUU                        P@UUUUUUUUUU                        P@UUUUUUUUUU                      �* P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      �* P@UUUUUUUUUU ��                     P@UUUUUUUUUU                        P@UUUUUUUUUU                        P@UUUUUUUUUU                        P@UUUUUUUUUU ��                     P@UUUUUUUUUU `U                     P@UUUUUUUUUU `U                     P@UUUUUUUUUU `U                     P@UUUUUUUUUU `U                     P@UUUUUUUUUU `U                     P@UUUUUUUUUU `U                     P@UUUUUUUUUU ��                     P@UUUUUUUUUU                      �* P@UUUUUUUUUU                        P@UUUUUUUUUU                        P@UUUUUUUUUU                        P@UUUUUUUUUU                      �* P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU ��                   V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      �* P@UUUUUUUUUU ��            �����    P@UUUUUUUUUU `U            (   �   P@UUUUUUUUUU `U            ZTU
   P@UUUUUUUUUU `U            �T%UI	   P@UUUUUUUUUU `U  &
UUUUUUWUUUUUUUUU}UUUUUUU�W�WUUUUUU|UUUu�� �5�UUUU  �WUUU   0 WUUU�     WUUUU  �\UUU� ��?0�UUW? ���3 WU�  ��0 W_=   � \�  �� \�U ��  W�W �<�0�U�_5 ?< ��UU5 � � WU� ��� W�� <�? WU� �� 0�uU�? �? p]U� ���\sU�� �sU5���00pU� ���� pUU3���� \UU300��? \U�00�  � pU�����pU� ���� \U5 ����?pU� <�?�0pUU����0\UU=0 �� WUU�� �� �UUUU0?�pUUUU�<<UU$UUUUU]UUUUUUUU�U�_UUUUUU�5�UUUUUW �� _UUUu�   <\UUUU=     p]UUU�  ��UUUUU5��?0�]UUU����3 WUUU= ��0 WUU�  � \UU�  �� \UUu ��  \UUU� �<�0 pUUUU?< � pU}UU� � p�U� ��� ��WU <�? �UU �� 0 �WU� �?  �UU7   ����UU� � ��UU� ���pUUU0��?� pUUU�0���? �UUU5��� �UUU���UUU<��� pUU� ?��? \UU� ����? �UUu����� �UUU?0���pUUU��0 pUUU� 3 _UUUU�0 3 �UUUUUU����CUUU%UUUUUWUUUUUUUUUUU]UUUUUUUU�_��UUUUUUU�<�U_UUUUU]  � pUUUU��   0 �UUUUU�      wUUUUU  �? \UUUUU ��� pUUUU������ �UU}U� ��� �UUU 0 �?  W�_u ��0  W�W� ��0  W�UU ���� �UUU� ��  |�_UUU<� _�WUU�<�p�UUU� ��� �UUU5 ��� �_UUU= � 0 �WUUU0��� �WUUU0�? 0 ?WUUU������UUU� ���<��UUU5����3�pUUU�������?�UUU�����? WUUU� 3�? WUUU���� �UUUU|���UUUU� ����UUUU� ��0pUUU��� �� 0�UUUUU�� � |UUUUU�0��WUUUUU���PUUUU$	UUUU�_UUUUUU��_UUUUU  �UUUW�    _UuU    \UU�     p]UU  ���UUU5 ���]UU �??WU�  �? WU  �� \�   �?� \5  ��� \� �?pU= � pU� � pU� �?\U5 �?�WU  ? \�  �?� p7 0 0�?�p� �� ��� ��?��U�������U����?�U5����� pU0�� pU0����?pU�����p�  ��??�pu ���pU= �0\U� � \U�< �WUU=�� �WUU��?<U$	UUUU�_UUUUUU��_UUUUU  �UUUW�    _UuU    \�U�     pUU   ��uU� �� WUU��� _U���  WU= ���UU �� �U�  �?  W] �< _U5 ? 0 \U� < 0 \� �00 \=0 ?�� p5� �<  p� ��  p� ����p� ��pU��� \U����?\U���� \� ��  p 0�� p5 ���??�5 ������� �?�?��� ����pU<� 0pU5    <\U� ��WUU�\ �UUUU�W�_U'
UUUUU]UUUUUWWUU]UUUUUU_UWwUUUUU��_U�WUUUU� �UUUUU� ��UUU�U p�UUUUU � WuU�U5    UU�U5  �p]U����UU�p����UUU���  WU��� WUU ��  _U� �?  \UU �< �Uu= ? 0 WUu5 < 0��U�5 �00��U� ?�� �U �<  �U5 ��  �U5� ���  �U�� ���  |U�0����\UU3����0\UW�� �?�\U� ��?<�|U= ����� pU ����� pU5  ��?? pU�  <�� pU�  �00 pUU  �� \UU  �� \UU� �??�WUUU�   �UUUUU�� �|UU%
UUUUUuUUUUUUUUUUUUUUU]UUUuUUUUU5U]�WWUUU��U7_UUUUU�W=�UUUUU ��WUUUW= � WUUuU5   \�UUU    �UU�W �0�uUU�5 0< WUU? � WUU     �]U  <   �WU ��  <WW ���? W]= ��?��_�� ����<��� �����\5����� ���5<0�������5 �������� ���<���� ��?  ��� ��3 ��U��<03�U���< 3sU� ��sU=� �pU5�� � \U5��?   \U  0 �WU�  �0< �UUU  � \UUU�?�_�_UUUU��U�WUU'
UU�UU�UUUUUU]UUUUUUUUU}UU�UUUUUU�Uu�_]UUUU�U�|UUUUU�_��WUUUU �7 _UUU]�  7 \UU�U�  < pUWUU5    �WUU}5���  �UU��00  \UU5�00  \UU� �� ? p]U�  ?��pWU� �����\]� ����? \u��0��? _U]<�����U]3�?�0\Us����?��U�<��?��U  ���0�U  ���0�U  �� �U  ���U5  ?��0�U� ����pU� � � pU��  � pUU �� pUU� �� pUU �� _UU� �? �WUU� ��pUUU� ��� |UUU��?�WUUUU?� _UUUUU�  �WUU(
UUUUUuUUUUUUUUUUUUUUU]UUUuUUUUUuU]�WWUUU��U7_UUUUU�W=�UUUUU ��WUUUW= � WUUuU5   \�UUU    �UU�W    �uUU�5     WUU?    WUU   �0 �]U   ���WU � ��0WW?0�� ?0W]��0� ?0_��� 0<�3����0<?�0\5��0 �??0�5<�  ��?0�5 �<��?0�� ?���?0�� ?������� ? ����U??���� �U<����? pU�����? pU= �?�� pU5   �� \U5    <  \U    0 �WU�  �0 �UUU 0< \UUU���_UUUU=  �UUUUU� < UUUUU���]UUUUUU�W_UUU&	U]UUUUUUUU5U�UUUUU��U�_UUUU�W=�UUUU �5�WUUW= �5 WUuU5   \�UU�    �U�W�  ��uU�5�� WU��� WU ��  \U�� \U ��  |W �?  p]= �< p�� ? 0 \�� < 0 W5� �00 W5< ?�� \5  �<  \� ��  \� ����p� ��pW��� pU���?p]�� ��� pu�� ��  ��� �  �5 ��� �� ��� �����?? �U  ����U  �?�0pU5  ��0pU� � 00\UU�? _UUU����W�_��;�;�;�;������x+x�x�~-^�\�^=^�_�W�_��;�;�;�;�����+�x+z�z�|-^�^�|=��WW}��U��V) Z* j. n��n��o��k��Z��V��U�jU�ZU�VU�VU�UU�UUeUU��U��V) Z* j��n��o��o��k��Z��Z��V��U��UUjUUjUUZUUYU��U��V�Z��j��o��o��o��k��j��Z��ZU�ZU�ZU�VU�VU�VU�VUUV
p � ��r���  �� �@ p /�@� �@� D@L�LB@ %S! ����@�BL�@Q$@$@���B$S�B  �@�`tBp�,�(                                                                ����@ @��@��@��B������@@��@$@""�@/r�@ �@@  @`�������@O��� ��
U]UU�V��k��~��Y�A^�U^��^ժWU�UUUUUU�U���W���_���^�>�z���z���z���^U��UU�WUU�_UU�zUU�_UU�zUU�_UU�zUU�VUUUUUUUUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �(      ��        UUU��ZiUh)@U�
                �
       UUU�PU�ZU�Z�            ��  ��      U�UUT���VU�             �Z����*     @UWUUWU�  X�               @UU����     @UWUUU�
                      _���    @UiUUU�                        TU�*    PUeUU��                           T�
   PU�VU�
                            U�  PUUZ��                            P�*  PUUj�
                             @U� XUU��                              U�* [UU��                              PU��kUUժ                                U��oU�+                                TU��UTU              P                PU��UPU           TUU@                U��UAU          @    U               TUjUEU          @     P               PUiUT          U     @               @UYUT         @  U  P                UUUU          P   UP                TUUUU          @   @U                 TUUUU           T  @                  PUUUU            PUUU                   @UUQQ                                   @UUPA                                  @UT                                  @UT                                   U U                                    U                                    U                                    U                                    U                                    U                                   U                                   U         �                       @U        �*                        @U   �
  ��                        @UU  �Z���Z                         @AUU  �U���j                         @EUE �Z@U�VU                           EUUE  �UU@U                            UUE  j                               @UUE �Z                               @UUQ �V                               @UUQ �U                                @UTUQ j                                PUUUP�Z                           �*   PUUUԯV                          ���*  PUUUիV                         ��V�� PUUU��U                         �ZUU��`UWU�ZU                         �j @U�*`�U�VU                        ��Z   TU��UT�V                         �    U�jUT�U                               P�ZAUP�U                               @UVTUQ�U                                UUUpAUU                                TUU�EQU                                PUE��                                 @UE�=                                 �uAUT�                                 �wQTT�                                 �PT�                                 �OPT�                          PU     �OAU=                         T @U    �OAQ                                �_EP                        @     A  �WAP                            P   �WDQT        ��               UT @  �VDTT       ����             P@      �RDPTU      ������           @E       �BPTU     ���U ��
            T   T    JTU    ��jU  ��
   �          P    :UEU    �ZU    �� �*        PUU     <@AU  ��U       ����                 <UQAU  �V        ��*                  <UUPU  j                              0TTU �Z   @                         0UU �V   U                         0T�U��jUU  T                          �TUu��ZUUUUU                          �EUu��VUUUU                           �EU\壪U_UUU                            �U\��jUU                               �U\��ZU                                UU\��VU                               @UU\�jU                                @UUT�ZU                                @UUW�UU                                @U�U�U             T                   PU�U�U            T                   PUUUeU           @ P    ���
          PUUUUU           P     �jU��          PUUUU                XUU����
 ��
   PTUUU                  PU���������  PPUUU   P    @U          TU�������* pAUUU   TU    T           PUUUUUU���|AEUU    U                TUUUUUU���EU    U  @              @UUPUU��  U    U  @                    TU��U  U    T  @                     UU��U  U    T @U                     @U��W@U     T @                     U��[ U     T                        TU�Z@U     TT                        PU�j@     TTU                        @U�jP     TP                       @U��P     U               U        U�ZP    @EU P             PP        UUZP    @EUU @T                   UUV@    @EUU  A                     TUUU@    @EUU                        TUUUE    @UU             T          TUUUE    @UU                        TUUUU    @UU             @            TUUUU    @UU                         TUUUU    @UU                         TUUUU    @UU                    @   TUUUU    @UE    T               PU   TUUUU    @EUE  @U               PE  UUUUU    @AUE  @Q      @       PEU  VUUUU    @AUE  @T       @      PEU  VUUUU    @AUE  PP        U      PEU  VUUUU    @AUE  PT              PEU�VUEUQ    @AUE  PT              PU�VUDUQ    @AUU  PT               PU�VUDUA    @@UU  PT               PU�V@UA    PTUU  TT               PUT�V@eA    UEU  UT               PUP�V@eA    UU  T               PUP�VP�AU    UU @T               PUP�VP�U   @UU @UU               PUP�VT�U   @AUU @UU              PUP�UT�U   @AUU @UEU             PUQU�U U�
T   @QUUT @UEU             UUEU�U U�T   PQUUP @UEU       PU    UU�U UU*T   PQUUQ @AUEU      @UU   U�j UUjT @UQUUQ PAUEU      TUU  @UU�j@UU�P PTQUUQ TDUEU      T  @UU�Z@UU�R TPQUUQ TUUU     @UUU TU��VPUU�Z TPUUUU TTUUU     PUUQUUAU��U PUU��PTUUUUU UUUUUQU PUUUUUUUUUU��j PUU��ZUUUUUUUUUUUUUUUUUUU�(                                                                                                                                                                                                                                                              �*                                      ��
                                      ��*                                      ��                                      ��
                                      �%                                      ��                                       �
                              PUU     h
                             @U      h)                             T   TU   ��    ��
                          @  ��  _��                     PU         V
 ����                           @   V	 p��                               Z	 |+                        T  U     X	 W                        @U        X	��                          UU      X9��                                    X�_�                                    h�V%                                    h�U*                                    `U�
                                    `EU                                    `EU                                    hEU                                     hUT                                     hT                                     �UT                            ��      �UT                             ����  �UP                             �������VQ                               oUU�*�VP                                 T���VP                                  ���V@                                  P��VA                                  @��VA                                   ��VP                                   T��                                   Ti�                                   TYU�                                    TUU�                                    PUU                                    PUQ   ��  �*                          PUT   �����                           TUU   �U���                           TUU  �ZU��U                            UEU  �VPZ                           @UEU   jU                              @UDU  �Z                               PTU  �V                    �  �*     PU  �V         T          �*  ���
   PU  �        P@U        �����U��  PU  j       @            ���UUU�
  PU �Z                     UUPU�*  `U� �Z           @             TU�  `U� �V      P  PU U              U� �UUe�V                         TU� ��U���U          @               @U��Vu��jU       @    @ @              U�>�VU��ZU           @@U               TU��VU��V        T  PU                PU��VU�ZU         U                   U��UU�UU           UU                  TU�\dU                                @UUUpQU                                 UUAAQU                                 UUPUU                                  t}PU                                  �]U                                  �_U                                  �WU                                  �PU                                   �PT                                    T            ��                      ]           ��                       ]      ��  �                       U     ���� ��                        UPU    ��UU�
�                        TQT�    �UUUU��                        TT�  �ZU @UU                        TT�  �V   P                         PU�  �U                               PU�. �V                     �
        @U�* �U                     ��       @U�*�ZU                       �*       @UT�)�V                       ��  ��*   UTU��U                        �* ���  UUU�ZU                        ����U�*  TUU�VU                          ��VUU�  TUU�Z                           TUP� TUU�V                           @ @�
 PUU�T                               U* PUUU                               T� PUUEU                               P�`UEQU                                @��UEP                                 U
�VT                                 U*�VT                                 U��jUP                                 U���UP                                 T��UA                    PU          TU��uA                   T           TU�iQE                  T  @U        PUUiQ                 @  @UU        @UUYP             �*  @   T   TU       UUYTU      �    ��   @       @      UU�P     ��� ��j     PU           TU5T     �U�*���U    P     @      PU    �ZU���jU      U    @       @UUA  ��jUUU��U        T  U        @UUQU4  ��VU@UU         @U            UUQQ� ��ZUU  P            UU          PUQ@� �VUU                             @UQ@���UUU                              @U@��ZU                               @U@��U                                @U@�ZU                                @U@�ZU                                 @UQ �V                                 @UQQV                                 PUQ QU                                 PUQ TU                                 PUAU�                                  PU�                                  P@�                                  PTT�                    *   �
        PUPU�                    �
 ���*       XUAE�                     �������*      XUAP�                      ��Z P��
  � XUEU�                      @�  ���  �
 h�UU=                           ��
����j�UU                            ��������UWU                             �������UWU                             ����VZ�ZWU                              ��ZVU�ZWU                              ��jiU�Z[U                               ���UUZ]U                 $UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUU�_��UUUUUUUUUUU��?��UUUUUUUUUU�  ���<UUUUUUUUU  ������WUUUUUUU3����?���|UUUUUU��  ���?�����WUUUU�0��������UUU�?��� ?�����_UU?  �� 0�<��UU  �0�   ?<<��WU <�3 ?  <00��\U 7��3 � 0  �� |U����0 �?     WUU� �   �\��U�pU� �  � \��U5\�� 7 ?� �? p�W�W ��?  � pUWU U��   ���W�_U� �UU����� ? |�_U3�UU��\U5�? ��sU�UU5� WU��0 �pUpUU �UUU� 7pU�_UU |UUU�� <pUUUU�  �WUUU�� 0\UUUU5  pUUUUU� �_UUUU5 �_UUUUU� �_UUUU5 |UUUUUUU5 �WUUUU5 WUUUUUUU \UUUUU5�UUUUUUU�  WUUUUU5�UUUUUUU�  WUUUUU�pUUUUUUU� �UUUUUUU_UUUUUUUU�UU$UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUU��UUUUUUUUUUUUUU���UUUUUUUUUUUUU��<�WUUUUUUUUUUU������WUUUUUUUUUU���?����UUUUUUUUU���?����UUUUUUUU������WUUUUUU� 0 ?��\UUUUU�  � 0�0pUUUUU3��  <?<<��UUUU��  ��0<00��UUUU�0��<�? 0  �?WUU����0��     \UU?  �? 0�   �pUU?   ?< 0�  � |UU  �0 � �? 0�UU  <���  � ��WU  ��p����� �?\U�� �\� pU� � pU5   W�  \U=�? 0�U� � �U� WU�����UU�_pU�UUU�0 �WUU�_� |UUU�  �WUUUUU5 �WUUU�  WUUUUU5 pUUUUU�  \UUUUU5 \UUUUUU=  pUUUUU5 pUUUUUU�? �UUUUU� �UUUUUUU� �UUUUU� �UUUUUUU� �UUUUUU�UUUUUUUU�UUUUUU5pUUUUUUUUpUUUUUU�_UUUUUUUU�_$UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��_UUUUUUUUUUUUUUU?��UUUUUUUUUUUUUU�<��_UUUUUUUUUUUUU����UUUUUUUUUUUUU����UUUUUUUUUUUU���?WUUUUUUUUUUU� ?<\UUUUUUUUUUU�?<0\UUUUUUUUUU� <?�0�\UUUUUUUUUU� 0<� �UUUUUUUUUU�? 0  �UUUUUUUUU���   ��UUUUUUUUU5 �  < WUUUUUU�� �? � \UUUUUU=�� < � �UUUUU����0 � ��WUUU�  0�� �? ��?\UUU3 �� < ���pUU��  ��0 ��\=�UU�0���  ��� \��UU?�� ? �< pU�W�   ?�  �� 0 �U�W?  ��   �< �  ��W  <�3     �<  �W  ��3 0    �   \ ��3 < 0 �   p�� 0 ?�< �    �5   ���� <    �� �  W��� 7   �U�_�U��������?pUU�UUU���U�U�_                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �(    @   � @UUUUUUUUUU@ V%              @  @ @ � @UUUUUUUUUU@ V%              @  @   � @UUUUUUUUUU@ V%             QTEQUU� @UUUUUUUUUU@ V%���*   ����  @     � @UUUUUUUUUU@ V%        �  @      � @UUUUUUUUUU@ V%        �         � @UUUUUUUUUU@ V�  ����  ���@      � @UUUUUUUUUU@ VU  `UUU  �UUEUUAQQE� @UUUUUUUUUU@ VU  `UUU  �UU @    � @UUUUUUUUUU@ VU���jUUU����UU @     � @UUUUUUUUUU@ VU  `UUU  �UU      � @UUUUUUUUUU@ VU  `UUU  �UU       � @UUUUUUUUUU@ ��  ����  ���TUU@� @UUUUUUUUUU@                     � @UUUUUUUUUU@                    � @UUUUUUUUUU@                    � @UUUUUUUUUU@  UDTQUP           � @UUUUUUUUUU@          ��UATEUEU� @UUUUUUUUUU@          ��� @     � @UUUUUUUUUU@          ��� @      � @UUUUUUUUUU@         ��  @     � @UUUUUUUUUU@ @QEUUT  �*Te       � @UUUUUUUUUU@        ��BUe@TU@E � @UUUUUUUUUU@          �*TUe      � @UUUUUUUUUU@        ��BUUe      � @UUUUUUUUUU@         ��TUUe       � @UUUUUUUUUU@ UUEE �*UUAe        � @UUUUUUUUUU@       �JUU e        � @UUUUUUUUUU@        �JUUAe��������� @UUUUUUUUUU@        �RUUUe          @UUUUUUUUUU@        �VUUUe          @UUUUUUUUUU@ PUUU �RA e          @UUUUUUUUUU@     P@  �V �*e          @UUUUUUUUUU@    @@  �VA�*e          @UUUUUUUUUU@    @@  �RU�*e          @UUUUUUUUUU@    @   �VUJe          @UUUUUUUUUU@ PTQU �VUJeUUUUUUUUUUUUUUUUUUUUU@       �RU�*eUUUUUUUUUUUUUUUUUUUUU@       �VU e            UUUUUUUUUU@        �VAUUe            UUUUUUUUUU@       �R UUe            UUUUUUUUUU@  PU �VAUUeUUUUUUUUUUUUUUUUUUUUUU@        �VUUPeUUUUUUUUUUUUUUUUUUUUUU@       �RU@eUUUUUUUUUUUUUUUUUUUUUU@        �VUUPeUUUUUUUUUUUUUUUUUUUUUU@         �VUUUeUUUUUUUUUUUUUUUUUUUUUU@         ������UUUUUUUUUUUUUUUUUUUUUU@ ����������BUUUUUUUUUUUUUUUUUUUUUUUUU@          �@UUUUUUUUUUUUUUUUUUUUUUUUU@           @UUUUUUUUUUUUUUUUUUUUUUUUU@           @UUUUUUUUUUUUUUUUUUUUUUUUU@           @UUUUUUUUUUUUUUUUUUUUUUUUU@           @UUUUUUUUUUUUUUUUUUUUUUUUU@           @UUUUUUUUUUUUUUUUUUUUUUUUU@           @UUUUUUUUUUUUUUUUUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU               UUUUUUUUUUUUUUUUUUUUUUUUU               UUUUUUUUUUUUUUUUUUUUUUUUU               UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU       PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU       PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU       PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU       PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ����
 PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU �    PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU �    PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��    PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�    PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� �  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� �  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� �  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�� �  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   �  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����                                     �                                     �                                     ��
 TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   �  TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   �                                      �                                      ��
                                     �U	                                     �U����   ���
  ����   ���
  ����   ��   �U�  �          �          �       �U�  �          �          �       �U�  ����  ���*  ����  ���*  ����    �U�  �UUU  XUU%  �UUU  XUU%  �UUU    �U�  �UUU  XUU%  �UUU  XUU%  �UUU    �U����UUU���ZUU����UUU���ZUU����UUU��   �U�  �UUU  XUU%  �UUU  XUU%  �UUU    �U�  �UUU  XUU%  �UUU  XUU%  �UUU    ���  ����  ���*  ����  ���*  ����    �                                       �������������������*����������������*                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �(            �  PUUUUUUUUUU                      ��
 PUUUUUUUUUU@UUUUUUU              �  PUUUUUUUUUU@UUUUUUU   ���
  �����  PUUUUUUUUUU@                  �  PUUUUUUUUUU@                  ��
 PUUUUUUUUUU@         �  ���*   ��U	 PUUUUUUUUUU@ ��*  ��
 U  XUU%   VUU	 PUUUUUUUUUU@     �   U  XUU%   VUU	 PUUUUUUUUUU@     �   U���ZUU����VUU	 PUUUUUUUUUU@  ����   U  XUU%   VUU	 PUUUUUUUUUU@  `UU�   U  XUU%   VUU	 PUUUUUUUUUU@  `UU�   �  ���*   ���
 PUUUUUUUUUU@ �jUU����               PUUUUUUUUUU@  `UU�                  PUUUUUUUUUU@ �*`UU�                  PUUUUUUUUUU@  ����       UQETQEU  PUUUUUUUUUU@         ��          PUUUUUUUUUU@ ���������*          PUUUUUUUUUU@ �*       ���          PUUUUUUUUUU@ V%        �*        PUUUUUUUUUU@ V%       U��� @EUUU  PUUUUUUUUUU@ V%       U�*    @    PUUUUUUUUUU@ �*       UU��"         PUUUUUUUUUU@         UU��         PUUUUUUUUUU@ �*  ����UU�*        PUUUUUUUUUU@     �   UU�*PTUU  PUUUUUUUUUU@     �   TU��      PUUUUUUUUUU@  ����   UU��        PUUUUUUUUUU@  `UU�   UUU�       PUUUUUUUUUU@  `UU�   UUU�         PUUUUUUUUUU@ ��jUU��
 @�@P@UUT PUUUUUUUUUU@  `UU�  �J�    @  PUUUUUUUUUU@  `UU�  �J�      PUUUUUUUUUU@  ����  �JU�      PUUUUUUUUUU@        �RU�       PUUUUUUUUUU@        �RU�@QDUTU  PUUUUUUUUUU@        �JU�        PUUUUUUUUUU@ UTU @U�        PUUUUUUUUUU@ @  @  ��UU�        PUUUUUUUUUU@    @   UU�    @    PUUUUUUUUUU@ @  @   UU� T@@U  PUUUUUUUUUU@ @  @   TU�       PUUUUUUUUUU@ BEQU��PU�  @     PUUUUUUUUUU@       XUTU�   @     PUUUUUUUUUU@       XUUUU�          PUUUUUUUUUU@       XU�����         PUUUUUUUUUU@       XUUU����������
 PUUUUUUUUUU@ FPUAQTXUUU(           PUUUUUUUUUU@  @   XUUU            PUUUUUUUUUU@  @    XUUU            PUUUUUUUUUU@      XUUU            PUUUUUUUUUU@      ��UU            PUUUUUUUUUU@ TUUP UU            PUUUUUUUUUU@      UU            PUUUUUUUUUU@     UUUUUUUUUUUUUUUPUUUUUUUUUU@     UUUUUUUUUUUUUUUPUUUUUUUUUU@      UU              PUUUUUUUUUU@ TATEU UU              PUUUUUUUUUU@ @      UU              PUUUUUUUUUU@ @      UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ @      UUUUUUUUUUUUUUUUUUUUUUUUUUUU@       UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ BTU@  UUUUUUUUUUUUUUUUUUUUUUUUUUUU@       UUUUUUUUUUUUUUUUUUUUUUUUUUUU@     ��UUUUUUUUUUUUUUUUUUUUUUUUUUUU@       UUUUUUUUUUUUUUUUUUUUUUUUUUUU@        UUUUUUUUUUUUUUUUUUUUUUUUUUUU@        UUUUUUUUUUUUUUUUUUUUUUUUUUUU@ ���������UUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@        XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@UUUUUUU XUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@UUUUUUU ��UUUUUUUUUUUUUUUUUUUUUUUUUUUU          UUUUUUUUUUUUUUUUUUUUUUUUUUUU          UUUUUUUUUUUUUUUUUUUUUUUUUUUU          UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ��            @UUUUUUUUUU��UUUUUUUUUU XU            @UUUUUUUUUU��ZUUUUUUUUU XU            @UUUUUUUUUU�	��UUUUUUUU XUUUUUUUUUUUUU@UUUUUUUUU��� �UUUUUUUU XUUUUUUUUUUUUU@UUUUUUUUU�`���UUUUUUUU XU           P@UUUUUUUUU�hUU�UUU�ZUUU XU           P@UUUUUUUUU�XU�ZUU��X    XU           P@UUUUUUUUU�X�
�VU% X    XU           P@UUUUUUUUU�X� �ZU%�X    ���
  ���*   P@UUUUUUUUU��*���U��ZAUUU           P@UUUUUUUUU�����U�jUAUUU           P@UUUUUUUUU%�
����*`UA      ���
  ��* P@UUUUUUUUU��� �
�bUA      XUU	  `U% P@UUUUUUUUUU�
����jUA      XUU	  `U% P@UUUUUUUUUU�����VUA     �ZUU���jU% P@UUUUUUUUUU�*����jUUA   �
  XUU	  `U% P@UUUUUUUUUUU� �
�UjUA      XUU	  `�* P@UUUUUUUUUUU�
(���bUA      ���
  �  P@UUUUUUUUUUUj�
�`UA ��
            P@UUUUUUUUUUUb) ���bUA VU	  ���*����  P@UUUUUUUUUUUb%��
hjUA VU	            P@UUUUUUUUUUUj����jUUA VU���          P@UUUUUUUUUUU�Z	�UUUUA VU	            P@UUUUUUUUUUU���jUUUUA �j	            P@UUUUUUUUUUU� �UUUUUA �
            P@UUUUUUUUUUU���UUUUUA               P@UUUUUUUUU         @ ����          P@UUUUUUUUU         @               P@UUUUUUUUU         @               P@UUUUUUUUUTUUUUUUUUU             �* P@UUUUUUUUUTUUUUUUUUU               P@UUUUUUUUU                         P@UUUUUUUUU           �*             P@UUUUUUUUU                       �* P@UUUUUUUUU                       V% P@UUUUUUUUU ���   ���
            V% P@UUUUUUUUU   �     �*           V% P@UUUUUUUUU   �     V%           V% P@UUUUUUUUU   ����  �V%           V% P@UUUUUUUUU   �UUU  XU%           V% P@UUUUUUUUU   �UUU  XU%           V% P@UUUUUUUUU   �UUU���ZU%           V% P@UUUUUUUUU   �UUU  XU%           �* P@UUUUUUUUU   �UUU  XU%             P@UUUUUUUUU   ����  ��*             P@UUUUUUUUU                         P@UUUUUUUUU   �*�������*             P@UUUUUUUUU ��                      P@UUUUUUUUU               '	UUUUUUU�UUUUWUUU�UUUU}U�U�UUUU�_�W�UUU�5|5\�UUUW=p�p�UU��|=p�UUs5 �p�W��5   \�\� 7  �p?\U���?\U�??�<pU��? <pU� �� <�]=��?� <pW5��� ?\5��_�7�� W�� w ��?\� ��?�\�  � �W �� w}�����?w�=� ��0��3�? ��0� �� ��0������?p��� | � �5�������<����\50�����\��0�����WU����sUU7�<��sUU5 < �_UU < �WUUU�����WU'	UUUUUU�UUUUUWUU�UUUUU}U��UUUUU�_��UUUU�5|5�UUUUW=p��UUU��|=�UUUs5 ���W��5   ��\� 7  ��\U���\U�??�pU��? �pU� ����]=��?��pW5����\5��_�7�� W�� w ��?\� ��?�\�  � �W �� w}�����?w�=� ��0��3�? ��0� �� ��0������?p��� | � �5���� ?��<��� <\50���� <\��0��� �WU��� |UU7�<�|UU5 < �UU <  |UUU�����U/UUUUUUU�UUUUUUUUUU� �UUUUUUUU�   _UUUUUuU   �UUUUUW�    �UUUUUU     �UUUUU�   �\UUUUUU���UUUUU� ���pUUUUU �� pUUUU�  ����UUU�  <��UUUU  � �UUUU=  << WUUU� �? 0 WUUUU��� 0 WUUUU�?�30�UUUUU3�?��pUUUU�����pUUUU= ?�� �UUUu�?���  WUUU�3�� WUUU���? \UUU5?���  \UUU�0�?�  \UUU����  \UUU�  ���� \UUU?  ���WUU� �?�� WUU�7 0��< WUU�5 �3� WUU� �00�UUկU���UU��V�0�   pUU� X��? �_UU?�VU ��UU��ZU��WUUUU�jUUUUUUUU� �ZUUUUUUUU  �VUUUUUUU� 
�UUUUUUUUU
��VUUUUUUUU% 
ZUUUUUUUU���UUUUUUUUU� �VUUUUUUUUU��UUUUUUUUUU�ZUUUUUU0UUU�|UUUUUUUUUU	|UUUUUUUUU�|UUUUUUUUU% |UUUUUUUUU	 |UUUUUUUUU
�UUUUUUUU���UUUUUUUU%� �UUUUUUUU	( �UUUUUUUU	*���UUUUUU�

�3 �WUUUU�	��  �WUU�`���   |UW�h���   �WU%X�*�    WW%���    |W%���   ��U���U �?0�U��UU��?0 Wi�UU5���3 WYUUU=?��0 WYUU�< � \UUU= <�� \UUu <��  \Uu�  <�<�0 WUUW �<< ��UUUU� ��� ��UUUUU300��� WUUU� 0��? \UW� 3�� 0 \UU=  ��� pUu  ���� pUU  ��� pUU  0��� pUU5  0��� pUU  ���< \UU   ?�� \UU�   ����\UUU  ���\UUU5  ���WUUU� ���� WUUU� 0��0 WUUUU0�?���UUUUU=0  ?�UUUUU��   pUUUUUU�  _UUUUUU= ���UUUUUUU��_UUUU.UUUUUU�VUUUUUUUUUU)�UUUUUUUUUU�ZUUUUUUUUUU)�UUUUUUUUUU�ZUUUUUUUUUU)�UUUUUUUUUU� ZUUUUUUUU�

�UUUUUUUUU)� ZWUuUUUUU�
`UU��UUU�
  uUU�UUU� ��_U �_U�
���_  �UU* U�   _U��_U   � p��WU ���U*�UW �?? W�UU5 �?  \�_U]� ��  \�WU�� �?�  p�UU<���  pUU �? �_UU�  �WUU50� �UUU���?� UUU���?0 �UUU5?��sUUU5 �?� �pUUU�� ��� ?pUUU�� ���\UUU�0 ��?�\UUU70����� \UUU50�� �? \UUU������ pUUU ���3� pUUU� ����0 pUUU�  ��� pUUUU ��? pUUUU  �0 pUUUU5  �  \UUUU� �  \UUUUU?  �  WUUUUU�  < �WUUUUUU?   |UUUUUUU� �WUUUU(UUUUUUUuUUUUUUUUUU�UUUUUUUUUU�WUUUUUUUUU5WUUUUUWU�_5_UUUUUuU=�5�UUUUU���� WUUUU5<  < \WUUU�     p]UUu�    pUU�U  � p�UU5_����UU5� �??��UU� ��?  �UU� � ��  pUUU��?�  �UUU���  �UUu=�� �UU���   �UU5��� pUU57��?� pUU57���0  \UU5�<�� \UU5 �<��  �UU5����  wUU���?��UU����� �UU]?���� �UU����� �UU�3���� �UU�0 ���  pUU?�  0  pU�? ����  pU�7 <��� \U������ \UU0���? \�_U=�?� W�WU�  �U�UU��  �U}UUU ���PU0UUU)_UUUUUUUUUU_UUUUUUUUU� _UUUUUUUUU	 _UUUUUUUUU _UUUUUUUU��_UUUUUUUU%� _UUUUUUUU	( UUUUUUUU
|UUUUUUUU�
|UUUUUUU���|UUU]UUU�h� |UUU�UUu%��(~U�__UU%��*�U=�5�Uu	������� Wu�&j��=  < \]�%jU�    p]��eU�     psbeUU�  � p�ZeUU�����VUU]��?? �VUUw���?  �UUU��� ��  @UUUU���?�  �UUUU����  �UUUU��� �UU���  �UUU�5��  pUUU�5�? pUUU7??� \UUU5��  \UUU5 ��?�  �UUU5 <��?  wUUU� ��� ��UUU� ��� �UUU]����?� �UUUu3�����UUU�0���?�UUU0��?<pUUU  �� pUUU5����  pUUU50��� \UUU�3���� \UUUU�3���? \UUUU�?� WUUUU5  �UUUUU��  �UUUUUU ���PU0UUUUUU�VUUUUUUUUUU)�UUUUUUUUUU�ZUUUUUUUUUU)�UUUUUUUUUU�ZUUUUUUUUUU)�UUUUUUUUUU� ZUUUUUUUU�

�UUUUUUUUU)� ZUUUUUUUU�
`UUUUUWUU�
  UUUUU}UUU� �UUU�W�WU�
�UUU|UU* u�� �5�UU��_U   W��WU     \U*�UU�     \U�UUU �? �_�_UU� ��� �s�WUW?���� �p�UU� ���  pUU= 0 �?  �_UU� ��0  �WUUU��0  �UUUU����  UUU]5��  �UUU]5<� �_UUUs<��\UUU���� ?WUUU����WUUU ��0��uUUU ����]UUU5��0?psUUU50������pUUU�0������pUUU�0����� pUUU3����< pUUU���0 \UUU � <0 \UUU |��� \UUU ����  WUUU� ���� WUUUU��� WUUUU��0�UUUUU� �pUUUUU5? �pUUUUU�� �?TUUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUU��? WUU�?<\UU� pUU�? pUU��0pUUU��_UUU=? \UUU� WUUU���_UU�? ��UU�� ��WU����W]�����Wu���Wu  Wu���Wu�����U�U���WUU����WUU}���WUU�� UU5 � �UU �  WU�����WUUUUUUUUUUU�WUUU��\UUU���\UUU�� \UUU��WUUU�� WUU��? WUU�?<\UU� pUU�? pUU��0pUUU��_UUU=? \UUU� WUUU���_UU�? ��UU�� ��WU����WU�����WU���WU  WU���WU�����U�U���WUuU���WUuU� WUu�� Uu5 � �U]�����W                                                                                                                                                                                                                                                                                                                                                                                                                                                  �(                TUU�T                                 PUU�U                                 @UU�U                                   UUUBU                                   TUUA                                   PUU@                                   @UU            �                     @UU           �*                      @UU          ��                       @UUT         ��
                       @EUUP        ��V                       @EUUP   ��� ��U                        UUQ  �V���jU                         UUQ ��UU��V                          TUA �jUUUU                           TPUE% �VU                              TPUU���U                               TPUU��ZU                                PAUU��U                                PEUU�jU                                @UU�ZU                                @UU�VU                                 @UU�UU                                 @U@U                                 @UTPU                                 @UTTU                        ��*      @UTTU                      ������    PUUUU                      ��*@UU����* `UU U                     ��   @U����
�UU@U                            TUUU���VUPU                              UU���VUPU                               UU��ZUTU                                PUU�jT                                 TU�jU                                  U�Z�                                  P�Z�                                  @�YU�                                  @�UU�                                   UUU�                                    TU�                                    TU�         �*                         PU�         �                         PU�     �
��*                          PUU�     ����                          PEU    ���Z�
                          TEU    �ZUUU*                          TEU   ��UU U�                          TEU   �ZU  @�                         TEU   �V   U*                         UAU  ��U    P�* @                     UAU  �V     U�               @U     U@U  jU     T�j            PUUU     UPU �ZU       @U                 TU   TU �Z                           @  UUU �V                     T       @EUUU jU                        TU  @ @EUU��ZU                     @   T@  @UEU��Z                      U    U   @UU��V                      P       PUT��U                       @UUU    PUP�jU                                PUU@�ZU                                 TUUA�ZU         TU                     TU�V        P @                    TTQEWV           U                   UUU]V            P                   E\U]U       T                       @QUpUuU             P                  @P@AQuU       @                       @UQEuU        U  @U                   PUTEU        P @                    PUu         @UU                     pUu                                 pU4U                                 p4PU                  �   �
         p5PU                  �
 ���*        ��PTU                    ���U��
       �E�PTU                    �UUUU��       �U�UU                   PU  PU�      �U�UU                         T�*       WPUU                        @U�      WQU                         U�*      _UAU                         PU�      \UQU                         @U�* �  \UQPT                          T�����  \QPP                          @U����
 \ATP                           U��U�� XUQ                           T�ZUU��ZEUQ            �
             @UUUU��jUuUQ            ��             PU@UU�jUU]Q      �*   �Z��               PU��UU]Q    ����� ��UU�*                TU�UUTQU    ��U骪�UUU�               PUUUUPU   ��UUU��ZU  �
               @UUUUPU  ��ZUUUUUU                    UUUPUPU��jU UUU                       UPU@U��jUU   @U                       TPUAի�ZU                             PPUA��jU                   UU       @5TUE��UU         @       T  U      �?TUE�VUU                     @      ?TU�UU        @         @          TU�ZUU        P          P     P      TU�UU�         P                @      TU�U�
                              TUeU�                  @           TUUU�                   @            TTUU��         @         @            UTUU��                   @            UTUU��                  @             UUUU�/                                UUUU�/                  @       @     UUUU�>       UU                @     UUUU��      P                 U     UUUU��                       @U     UUUU��        @               T @    UUUU��     @                         UUUU��     T                         UUU���    @                          UUU���          T        P              UUU���        @U       P              TYU���         @Q       @             T�U���  @      @T                @U   �jU��� P      PP        T      P   �ZUU�� P      PT       P@U     P    �ZUU�� T      PT              P    �VUU�� T      PT             TT    �TUU��       PT      @  P    TT    �TUU��       TT      @   @    TT    �TUU��       UT      @        TT    �TUU��       T      @       @TQ    (UiU��      @T     PU       @ TQ    (U�U�� @   @UU     U        P TQ    (U�U��     @UU   @         TQ    *U�V��/     @UEU  P          TQ   *U�VU��    @E@UEU      P     TT  �*U�ZU��   @E@UEU       UU     UT  �*U�ZU��
   @E@AUU      PQU   PUPT  �
�ZU��+ P  @EPAUU      TUU   TUQQ ��B��VU��� @ @TDUU     @TUQ @UUUQ ��Z��VU���Z P PUTUU     TAUUEUUUUUUQ�����������  TUTUUU  UUUUAUUEUUUUUUU�������������fUUUTUUUQUU�(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         TU                                    P P                               U       AU                            @Q T  @@                          @ PU@U                              @          T                                                             @           @ P                                                                            P                                      TU                                                                          @UU                                   TU                                   TU                       @                                      T          T@                          U         @UU                          @     U  TUU                                PU@U                             P    UUUU                              @U  U UU                               @UUU @                                 TUU                                                                                                                                                                       U@                                    P T                                  P   T                                      P                              T     PUP@U                                   UTU                                     @U                                                               E           PUU                         T         P                           P                                     @U      @U                             @@UU @UU                              UUUQU TUU                               PU TUU                  @U                 T                 UUUT                                  TU  UUUU@UU                           @    PUUUU                           @      U   TU                                       UU                                      @                     @              PU                     @              UU                      @             TU                                    @U                                    U                          T         TU                           @UUU      UU                            PUU    @U                               TUU  PU                                 UU TU                                   UU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             PU                                @UU @U@U                              TU  P   P                               P                                @  T    TU                          P   @     TU                                     TU                                    @UUU                                   PUUU                                     @                                    T                      P              P                       @PU          TU                         UUU        @U                          @UU   PUU U                            @U PUUUUUU                               TUU  UU                                @U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               $UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUU��UUUUU��_UUUUUUU57WUUU�0 pUUUU�UU\UUU0 �UUUU�_U\UUU�? � WUUU?���\UUU��\3WUUU   \���\�_UUU    W?���<|�_UUU ����?<��=\UUU � ?0�0����\UUU= <<�0���<��UUU�?���?�� ��UUU� ?<�? ��UUU�U<0<�� WUUuU� <<    ��WUUUU�<<   \�WUU�U�<< 0< p�_UU5W ?<0  ��\UU5�  ��� � ?pUU�� ��� �  <pUU5�_?  � ���UU5pU�0��|�� ��UU�_������ pU� �WUUU�� �� pU�p\UUU� �� |� pUUpUUU�\��W� _UU=p��UU��WUU� �WUU?p��U���UUU� �UU�p��U pUUU�?pUU� \U��0  _UU�  _U�0 WUU5 �UUU WU5 WUU5 |UUU�UU5�UUU5 WUUU�UU5pUUU���UUUU���UU��_UUU$UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUU��W��UUUUUUUUUUU� �����WUUUUUUUU5    ��\UUUUUUUU�  ?��<�WUUUUUUUU��?0��|UUUUUUU�� ��0���UUUUUUU�  ?�� ��_}�WUUU�0<<�� �  ���?|UUU������ � ���?�WUUUW���� � �UUUUU?0��  0<<0��WUUUU<0�0 �0<��\UUUU00�0 �00�� |UUUU � �0   WUU]��<0�?0   W��UUs� �<�?0 � W��UU��W� ��0� \�WU= \U?� �  pUWU WU=�� �?  �W�_U�UU� < � � \�_U�UU������� p�sUUUU�  < �� �  ��pUUU�� ? pU� ��pUUU  �� \U����pUUU�  � WU� �  7|UU�0 � ��UUU� 7UU� ?  pUUU�_5 �UUU�5� \UUUU� �_UUU���WUUUU5  \UUUUUUU|UUUUU WUUUUUUU_UUUUU�  WUUUUUUU�UUUUUU� �UUUUUUUUUUUUUUU��UU$�UUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUU��WUU�UUUUUUUUUUUU� �_���}UUUUUUUUU  ����WUUUUUUUU � �?�\UUUUUUUU �?�����WUUUUUUU  ����|UUUUUUU� �?��?��_UUUUU�  ?0��?�����WUUU5 <�������?|UUU5��<�� ?���?�WUU5w���� 0�<��UU�UU�?�  <?<<��WUUUU�0 � 0<00��\UUUU�0 �? 0  �� |UUU��?0��    WUUW53<�  < \��U�\� <��? � p��U��3  �  � � ��W5   W�  �  _W����U�� �? � p�_U? _U��<��� ��_� �UU=� ����  �s� ���� p�� 0 �pUp  � \U�?  �pU�_   ?�WU�?� �_UU��    |UUU=��  WUU50   �WUUU��W \UU5   UUUUUUU5 pUU5 ��UUUUUUUU� �UU���_UUUUUUUUUU�UUUUUUUUUUUUUUU�0�UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU�;UU������������_UUUU�������������_UU�?��W���������sUU�? �WUU��������UU�?��UUUU����U���UU�?�UUUUU��U��U��?�_UUUUUUUUU��UU��?�_UUUUUUUUU�WU����WUUUUUUUUU�\U����UUUUUUUUUUs5\U����UUUUUUUUUU��_U����UUUUUUUUUUWUU���UUUUUUUUUU�UUU���UUUUUUUUUUUUUU���UUUUUUUUUUUUUU���WUUUUUUUUUUUUU���WUUUUUUUUUUUUU���WUUUUUUUUUUUUU��?�_UUUUUUUUUUUUU��?UUUUUUUUUUUUUU�� �UUUUUUUUUUUUUU���WUUUUUUUUUUUUU��<WU�WUUUUUUUUUU��<_U=|UUUUUUUUUU��?0U�UUUUUUUUUU���0��  WUUUUUUUU����  \��UUUUUU�����  ���WUUUUU����   ���WUUUUU����?0    ��_UUUUU�����    ���UUU������  �����sUUU������  ��W���UUU������  ��W���UUU���<�?  ����UUU�_��<�� �����UUUU�_��<���� ��WUUU�_U�< ��� �\UUU�_UU? ��? ��5\UU��_UU? ��? ���\UU��UU� �?�� �WWUU���WUW<<� ��UUUU��_UW<0<��UUUUU�sUW���3��UUUUU�5�pU]00��UUUUUU5�pU]��p�UUUUUU5W_U]00puUUUUUU�UUUu00puUUUUUUUUUUu0�p]UUUUUUUUUU�5�0p_UUUUUUUUUU����?\WUUUUUUUUUUU_�� �UUUUUUUUUUUU��� �UUUUUUUUUUUUU���uUUUUUUUUUUUUU5�\_UUUUUUUUUUUUU��WUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUU�_UUUUUUUUU�uU�u���}���]���]���_U�WU�_WUpWU��W���W�?�W�?�W���U�pUU_UU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �(          �P%T		   P@UUUUUUUUUU ��            �P%T
	   P@UUUUUUUUUU               �Q)T
	   P@UUUUUUUUUU               �Pi�
	   P@UUUUUUUUUU   ��          �Q*�	   P@UUUUUUUUUU               �Qj�
	   P@UUUUUUUUUU               �Qj�	   P@UUUUUUUUUU     �          �Qj�	   P@UUUUUUUUUU     V          �Qj�	 �* P@UUUUUUUUUU     V          �Qj�	   P@UUUUUUUUUU ����V          �Qj�	   P@UUUUUUUUUU     V          �Qj�	   P@UUUUUUUUUU     V          �Qj�	 �* P@UUUUUUUUUU     �          �Qj�	 V% P@UUUUUUUUUU                �Qj�	 V% P@UUUUUUUUUU                �Qj�
 V% P@UUUUUUUUUU                �Qj�� V% P@UUUUUUUUUU `UEU          �Qj��  V% P@UUUUUUUUUU               ����*  V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      V% P@UUUUUUUUUU                      �* P@UUUUUUUUUU `UTT                    P@UUUUUUUUUU    �                   P@UUUUUUUUUU     �                   P@UUUUUUUUUU   ��                   P@UUUUUUUUUU   ��                   P@UUUUUUUUUU `UT�*                   P@UUUUUUUUUU   �J                   P@UUUUUUUUUU    �J                   P@UUUUUUUUUU   �R                   P@UUUUUUUUUU   �V                   P@UUUUUUUUUU `UU�R                   P@UUUUUUUUUU  @ �V                   P@UUUUUUUUUU  @ �V                 �* P@UUUUUUUUUU  @ �R                   P@UUUUUUUUUU    �V                   P@UUUUUUUUUU `U�V                   P@UUUUUUUUUU    �R                 �* P@UUUUUUUUUU    �V                 V% P@UUUUUUUUUU    �V                 V% P@UUUUUUUUUU    �R                 V% P@UUUUUUUUUU `�V                 V% P@UUUUUUUUUU    �V                 V% P@UUUUUUUUUU    �R                 V% P@UUUUUUUUUU    �V                 V% P@UUUUUUUUUU    �V                 �* P@UUUUUUUUUU    ��                   P@UUUUUUUUUU ����B                   P@UUUUUUUUUU    �@                   P@UUUUUUUUUU     @                   P@UUUUUUUUUU     @                   P@UUUUUUUUUU     @                   P@UUUUUUUUUU     @                   P@UUUUUUUUUU     @                   P@UUUUUUUUUU     @                   P@UUUUUUUUUUTUUUUUU                   P@UUUUUUUUUUTUUUUUU                   P@UUUUUUUUUU                          P@UUUUUUUUUU                        �* P@UUUUUUUUUU       ��
  ����   ���
   P@UUUUUUUUUUUUUUUUUU
      �        P@UUUUUUUUUUUUUUUUUU       �        P@UUUUUUUUUUUUUUUUUU  ���*  ����  ���* P@UUUUUUUUUUUUUUUUUU  XUU%  �UUU  XUU% P@UUUUUUUUUUUUUUUUUU  XUU%  �UUU  XUU% P@UUUUUUUUUUUUUUUUUU��ZUU����UUU���ZUU% P@UUUUUUUUUUUUUUUUUU  XUU%  �UUU  XUU% P@UUUUUUUUUUUUUUUUUU  XUU%  �UUU  XUU% P@UUUUUUUUUUUUUUUUUU  ���*  ����  ���* P@UUUUUUUUUUUUUUUUUU                    P@UUUUUUUUUUUUUUUUUU                    P@UUUUUUUUUUUUUUUUUU                    P@UUUUUUUUUUUUUUUUUU QUE@           UU$ P@UUUUUUUUUUUUUUUUUU       ����       P@UUUUUUUUUUUUUUUUUU      ����*      P@UUUUUUUUUUUUUUUUUU      ������      P@UUUUUUUUUUUUUUUUUU     ��  �*     P@UUUUUUUUUUUUUUUUUU UUD  �*TeU���  UE$ P@UUUUUUUUUUUUUUUUUU    ��BUeU�*     P@UUUUUUUUUUUUUUUUUU    �*TUeUU��"     P@UUUUUUUUUUUUUUUUUU   ��BUUeUU��     P@UUUUUUUUUUUUUUUUUU   ��TUUeUU�*    P@UUUUUUUUUUUUUUUUUU UUP�*UUAeUU�*U% P@UUUUUUUUUUUUUUUUUU  �JUU eTU�� @  P@UUUUUUUUUUUUUUUUUU   �JUUAeUU��     P@UUUUUUUUUU          �RUUUeUUU� @  P@UUUUUUUUUU          �VUUUeUUU�  @  P@UUUUUUUUUU         UUU�RA e@�UU% P@UUUUUUUUUU@UUUUUUU  @ �V �*e�J�   P@UUUUUUUUUU@UUUUUUU  @ �VA�*e�J�   P@UUUUUUUUUU@        @ �RU�*e�JU�   P@UUUUUUUUUU@          �VUJe�RU�    P@UUUUUUUUUU@       EU�VUJe�RU�UU! P@UUUUUUUUUU@         �RU�*e�JU�    P@UUUUUUUUUU@  ����   �VU e@U�    P@UUUUUUUUUU@  �  �   �VAUUeUU�    P@UUUUUUUUUU@  �  �   �R UUeUU�    P@UUUUUUUUUU@ ��  � U�VAUUeUU�U  P@UUUUUUUUUU@ V�  �    �VUUPeTU�    P@UUUUUUUUUU@ V�  �    �RU@ePU�    P@UUUUUUUUUU@ V����    �VUUPeTU�    P@UUUUUUUUUU@ V�  �    �VUUUeUUU�     P@UUUUUUUUUU@ V�  �    �����������    P@UUUUUUUUUU@ V�  ������BUUUUU����* P@UUUUUUUUUU@ V%       �@UUUUU(     P@UUUUUUUUUU@ V�*��     @UUUUU      P@UUUUUUUUUU@ V%        @UUUUU      P@UUUUUUUUUU@ V%        @UUUUU      P@UUUUUUUUUU@ �*        @UUUUU      P@UUUUUUUUUU@          @UUUUU      P@UUUUUUUUUU@          @UUUUU      P@UUUUUUUUUU@     UUUUUUUUUUUUUUUUUUU@UUUUUUUUUU@     UUUUUUUUUUUUUUUUUUU@UUUUUUUUUU@            UUUUU        @UUUUUUUUUU@            UUUUU        @UUUUUUUUUU@            UUUUU        @UUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ �*   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ �*   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ V%   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ �*   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@                                     @                                     @                                     @     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU     UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU     �(                                                                                                                          ���*  ����  ���*  ����  ���*  ����        �          �          �           �          �          �    ��
  ����   ���
  ����   ���
  ����   ��UU	  `UU�   VUU	  `UU�   VUU	  `UU�   VUUU	  `UU�   VUU	  `UU�   VUU	  `UU�   VUUU���jUU����VUU���jUU����VUU���jUU����VUUU	  `UU�   VUU	  `UU�   VUU	  `UU�   VUUU	  `UU�   VUU	  `UU�   VUU	  `UU�   VU��
  ����   ���
  ����   ���
  ����   ��                                                                                                                               @QUTEDUUU       UTQUTUQQ   ��*            ����   @ @  @       ����
          ����*  @    @     �������        P   ������  @ @  @     ��� ��
       ��  �*   @  @    ���
UY��  TUEQTUE �*TeU��� TUEQUU �*�PUYU��
      ��BUeU�*       ��B
UUYU��         �*TUeUU��"     @ �*TRUUYUU��"       ��BUUeUU��    @��BUTUUYUU��      ��TUUeUU�*     ��TUUUPYAU�� TUPT�*UUAeUU�*EPUUT�*UUU@Y UU�*    @ �JUU eTU��  @  �JUUUUPYAUU�*       �JUUAeUU��    @   �JUUUUUYUUU�*     @ �RUUUeUUU�  @  �RUUUUUYUUU�*      @ �VUUUeUUU�   @  �VUUQ@Y PA�*AUUT�RA e@�TUUUU�RA@�JY�R �*     �V �*e�J�     �V �Q�JY�RA�*@    �VA�*e�J�    �VA�U�JY�RU�*@    �RU�*e�JU�    �RU�U�RY�TU�*@     �VUJe�RU�     �VUU�RY�TU�*EUUQU�VUJe�RU�UUUQU�VUU�JY�RU�*      �RU�*e�JU�  @   �RU�U@Y PU�*      �VU e@U�  @   �VUQUUYUUA�*      �VAUUeUU�  @   �VAU@UUYUU �*      �R UUeUU�  @   �R UQUUYUUA�*UU �VAUUeUU�TUUUUE �VAUUTYUU�*@      �VUUPeTU�     �VUUUPYTU�*@     �RU@ePU�     �RUUTYUU�*      �VUUPeTU�      �VUUUUUYUUU�*        �VUUUeUUU�        �VUU��������*       �����������       ����AUUUUU@�����������BUUUUU����������BUAUUUUU@
        �@UUUUU(        �@UAUUUUU@          @UUUUU          @UAUUUUU@          @UUUUU          @UAUUUUU@          @UUUUU          @UAUUUUU@          @UUUUU          @UAUUUUU@          @UUUUU          @UAUUUUU@          @UUUUU          @UAUUUUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUAUUUUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@UUUUU              UUUUU             U@UUUUU              UUUUU             U@UUUUU              UUUUU             UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                                                                                                                        UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                                                                                                                                                                  ����  ���*  ����  ���*  ����  ���*   �          �          �           �          �          �         ���   ���
  ����   ���
  ����   ���
  ��UU�   VUU	  `UU�   VUU	  `UU�   VUU	  `UUU�   VUU	  `UU�   VUU	  `UU�   VUU	  `UUU����VUU���jUU����VUU���jUU����VUU���jUUU�   VUU	  `UU�   VUU	  `UU�   VUU	  `UUU�   VUU	  `UU�   VUU	  `UU�   VUU	  `U���   ���
  ����   ���
  ����   ���
  ��                                        �����������������������������������*����                                                                                                                                                                                                                                                                                                                                                                                                     ����
                                  �   (                                  �U@P�                                   IUR��                                   	UB��                                  `	UB��                                  `�B��                                  `
�F��                                  `�B��                                  `�F��                                  `�F��                                  `�F��                                  `�F��                                  `�F��                                  `�F��                                  `�F��                                  `�F��                                  `�F��                                  `�F��                                  ��F��                                  ��F�)                                   �F�
                                   ����                                                                                                                                                                                                                                                      (
UU�UU�UUUUUUUUUuUuUUUUUWUUUUUUUUUUU�UUWUUUU]UUUUWUUUUUU�UUUU�UUWUUUUUUUUU_UUUUWUUW��WU]UUUUW� U��UUUU� pU�WUUUW5 ��wUUWU�  � |UUUu�    �UWWu5  �pUUU���pU]U5 ����UU]5 �� �UWu� ��p�UU� �? �UUU���3��U�<�? �U� �30 WU� �? 0 wUU�� 0 \UW �� \UU <?0 \U]= �  _U�� ���  WUU7 �  WUU ��  WWU �� TUU���� WU]=���UUU5����0UUU�<  3�UUU�����?pUUUU ���?pUUUU����?pUUUU= ���_UU*UUU�UU�UUUUUUWUWUUUUUUUUUUUUuUUUUUuU�UUUUUUUUuUUUU]UUUUUUU�UUUUUUUUUUUUUuU�UUUuUUUU}UUUUUUU]U��UuUUU��_U?�UuUUUU�pU�WUUUUU7��  WuUUUU� �UUuUu�    �UWUUUU    WWuU]U  ��UUUU��� WUUu� ��� W]U�U�� �WWUU� ���uUU�� �? �uUU�5��3 �UUU5�? �UUU7�30 �UUU�? 0 pUUU�� 0 puUW �� pUUU= <?  _]U]5 � ��UUU5 ���  wUU�5 �  |UU ����UU50 ���UU� ������]UU?�?�U]U����WUU< ��WUU���?��WUU= ��� �UUU5 �� �UUU5� ��� \�WU�� �� TUU�����*�����*(    ((    ((�?�?((�?�?((<<<<((<<<<((���?((���?(( <<  ( <<  (�����(�����(<<<  (<<<  (�?<  (�?<  (  <  (  <  ��*<  ��*<     <  ���*���*(�((�((��((��((�"((�"(���*���*        ��������   <  ��*<  ��*<  (  <  (  <  (�?<  (�?<  (<<<  (<<<  (�����(�����( <<  ( <<  (���?((���?((<<<<((<<<<((�?�?((�?�?((    ((    (�����*�����*   <��*<��*<( (<(((<(�*<(  <��*<��*<  (<�*(<(((<( (<��*<��*<   <��������        ���*���*(�"((�"((��((��((�((�(���*���*C      @�   �    �@��   �    @��� ��    @� �� �    @��" ���    Т� ���    Q��� �@��    �B�@!H �    9F��  ��$�    D� ��� �    @�� �  ��    @� �  E    @� � @F    @��"��&    AP������@�    � �  �                     �       .� �  0    B � ��   N� �!@ ��  (�L�@  (��D ��@ 0(p � @ �� 0(O� � @H�(A ����4�� (AR � H   (M� �PIB   (A� �PJ�    (A ��IB�@   �����"��    ��������    �                        �  ��@   �  � ���@!  � � �P��@�@�  ����P��B�@H�  �����D�Q�B*�� H �-���C@0� H �� �����10�( ����Q�@ȃ��Ȁ���F���r  ��������A�    �����B�A��  ! �@���B�@�  �q �����D��    ���zB�D��    ��(B����   � @ �@� �   @                    �         ���� ��        D@ ��!        �� ��!        F� ��        Mg  �00      �R��� `      O���� `      A @�!`      O� �$A0      A @$�        O� H $@        )  H@$�        $�D��        %��B(        ��  A        v                 ���      ����Q!@�!��    @  R!@L�""    O�  ��!B! ""    @  �@)�"""    �� ��P)B��""    @���B)B� ""    O�  �R)B�!""    @  �R)B��""    O�  �Q)B� !�    A  �A)B� �    ! ���      !��NԈA�0��    �  "%@@��        @�                       @    @     P  @@@     ��@ ���B     �@   �B     @�  �B   @� �0  ��B ��! 0����  -�  A@  !    G@  )�    A@  )�    A@  ��  @  a�@ �@��  ��  � �@��x�  @  �@@���(        @                     @ �     ���$@���  ��AD@ ����  �@���O���@   @��U@(@ �U�@��"0�@����t@ ����0@�� QDB��   @��QO� �� @ �@�� �D@������ @����D@����@ 	����D@����@  @�B@����@  �@��@���� @  �@������ P  @@���  ����     @0                 �  �@@   �  �@�  �@�  �  �@� �@��  � �@���O�  ���O��� HA�  �� HADH�hA	0DH�hAD��^��`D��^�D	 J@�`D	 J@D��JB�`D��JB$N��0$N�B
 HB��  B
 HB�	�HB�  �	�HB�D  �D�8DA�  ��8DAD C@��  D C@   @@�      @@                @  �  �   ���". �  �����B ��  �pAPB� B  @� *��!B@	�����b0��� r�1R0D��@N�!BD���B1�!B D�@BQ�aB ���b?rOQ��B D�B@I� B  @��@��$B  @�@@B�B  (�� ApQ��B�  �  �@�� B                      �  � �@ ��� �"�@$���O��@,�@B"�@ O�(O�J� �.�HA �@b"�����RhA ���^���R^� @@ �N�J@(�!O�L��` JB$��A@D�_�N�"�AO�Db�@ HB!@AL�B�DHB��!D�(EbD�`!�!D@"EEDA@A�L� AA�C@ �D ��H�@@                  �  �� @�@  �� �"����@�@  ���"��!)@�@  � ��!)@O���" "���)@HA0����"��0��hA0����� %@^��@ � #@J@ ��   �!!@JB � �� $A��N� �� b $�!@HB  � B $@!@HB  � � $�!@D�  �@ �!BDA  ���� A (-�C@  �   � � @@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �*                                      ��                                    Z�                                   �[Ze
                                   �Ve                        @U        �Ve                   PU @U P       ��UU=                    UU   U      ��UU9                  P   TA   P      ��UU9                           @      �UUU9                                  �UUU�                 @                ��UU�
                @                 �VUU�* PU                            P�VVU�UT@                    UE      @VU� U              T       TUU    T  UUe    @U          PU     @U           U      P           U @UUU           @    TU           @U UT                 @               U                   @U                            @        P�                                   @T�                            �      PWU�                            �oUm    �WV�                            �kWUU @�[U�                            �UUUU�VU�                           �VUU���VU�                           �jUUUU���UU�                           �jUUUU���UU�                           �[UUUUU�UU�>                           �[UUUUU�VU�:                           �ZUUUUU�VUZ9                           �VUUUU�Z�U)                           ��ZUUUU�Z�V)                           �ZUUUUU��Z�U�                           �ZUUUVUտZ�U�                           �VUUUZUկZ�U�                           �VUUUZUկV�U�                           �VUUUZU��YUU�                           �VUUUYU��VUU�                          �VUUUYUU�VUU�                          �VUUUYUկUUUZ                          �VUUU�UկUUUZ                          �VUUU�UկUUUZ
                          �VUUU�UկUUUZ
                          �UUUU�U��UUUZ
                         ��UUUUiU��UWUV	                         ��UUUUi���UWUV)                         ��UUUUU�V�V^UU)                         ��VUUUU�U�Z]UU)                         �VUUUU�UUZYUU%                         �VUUUU�UUZUUU%                         �VUUUUiUUZUUU�                         ��VUUUUYUUZUUU�                        T��VUUUUYUUZUUU�                        T��VUUUiUUUZeUU�                        P��VUUUzUUUjeUU�                         ԫVUUUzUUUi�UU�                         @�UUUU�UUUi�UU�                          �UUUU�UUUi�UU�                          UUUU�UUUe�UU�U                          TUUU�kUUe�UU�U                         @UUU�kUUU�UU�VU                         UUU�kUUU�UU�ZU                         UUUիUUU�UU�jU                         UUUիUUUUUUUjU                         UUUկUUUUUUUj                          UUUU�UUUUUUUj                         @UUUU�UUUUUUU                          PUUUU�UUUUUU                           PUUUU�VUUUUU                           @UUUU�VUUUUU                             TUUU�VUUUUU                              TUU�VUU                               PTU�VU                                  PU�VU                                  @U�ZU                                    @�ZU                                      U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ���                                 ����W���  ��  �?  �?  ��  ��  ��     ��_U �@_U�   �  �       �������+  �@ T?    �        @U��V��*  �   4  0  �    0  0   @��V�W�  �   �� ���00�0� �� �    ��QTU��  �   ���0�� 0000��0���0�    �k P�V � }  �0 �� � 0 0    �k   uE � }  ��0 �� � 0 0    �Z   �A � }  �� � �      �Z   �A � }  ��� � � � � � �    �   � � } ��                 �   �  � } ��                 �   �  � } ��>  0         0   0   �   �  �@}  �W>  � �� ��  �  �   �   �  P@i PV> � 0 0  0  � 0 �    �   �  `  � @�> 0    0  0 0 � 0    �   �
  `  � @�: 0 �  �  � 0  0    U   �  �  � @�: � < < � �   %   �*  � � @�: � �       �k  � �[ @�: 0 � � 0 00       �k    �oP�� 0 � � 0 00       ԫ     ��T�� �� 00 00 �� 0��  @@  ի     �����  ? � �  ? 0 ?  @    ժ     ��U���   0   0   0   �    @    @��    ��U���   0   0   0   �         @��
    ��U���   �   �   �    �(                          ��                                     ���                                    �Z�/                                    �Z��                                  ��Z��                                  ��VU�                                  ��VU�                                  ��VU�                                  �kUUz?                                  �kUUy?                                  �jUUi?                                  �jUUi�                                 @�jUUe�
                               @@jUUe�
                              @ @VUUe�*                                  PUe��                                   Ue��j                                  Ue�j�                            @      Pe�j�                            @       �j�                                    @j�                                    j�                            P P     Pi���*                           UUUPUUUj��U�                           �oUUUUU��ZU�%                           �oUUUUU��VU�%                           �VUUUU��VV��                           �UUUUU��VU��                           �kYUUUU��VZ�                          ���jUUUU��UY�                          ����VUUU��VY��                          ����ZUUU��ZU��                          ��[�ZUUU��VU��                          ��WUiUUU��UU��                          ��VUiUUU��U���    U                    ��VUiUUU��V���    @U                   ��VUeUUU��V���      U                   ��VUeUUU��VUU�    @U                   ��VU�UUU��VUU9    PUU                  ��ZU�UUU��VUU�    U                    ��ZU�UUU��UUU�                         ��ZU�UU���UUU�                          ��ZUUVU�Z�WUU�                         ��ZUUVU�ZYUU�                         ��ZUUVU�ZUyUU�                         ��ZUUVU�ZU�UUU                         ��jUUVU�jU�WUU                         ��jUUU��iU�WU�                         ��jUUU�[eU�WU�
                         �ZUUU�ZUU�WU�
                         ��ZUUU�ZUU�WU�
                         �VUUU�VUU�WU�
                         �UUUU�VUU�WU�&                         �UUUU�VUU�WU�%                         �UUUU�jUU�_Ui�                         ��UUU��jUU�^U��                          �UUU���jU�^U��                          �UUU�j�jU�nU��                          �UUU�jUVUU�U��                          �VUU��UVUU�U��                          �VUU�jUVUU�U��                          �VUU�jUUUUzV��                         �VUU�ZUUUUzVU�                        ��VUU�ZUUUU�VU�                        ��VUUUZUUUU�VU�
                     PUU��VUUUZUUUU�VU�
                    @  ��VUUUZUUUU�VU�                       �ZUUUZUUUU�VUU                  PU   �jZUUUZUUUU�VUU                 U    U�ZZUUUYUUU��VUU*                P     PU�ZZUUUUUUU��VUei                     PU�ZeUUUUUUU��ZUe*                     @U�ZeUUUYUUU��ZU�
               @       �Z�UUUYUUU��ZU�
               @         U�UUUUUUU�VZU�               @         T�UUUUUUU�VUU�V                        �VUUUUUU�FUU�V                        PUUUUUUU  PU�V                          TUUUUU  TUU @              P            UUU @UUU PU               @            U  PUU                                  P  @                 @                   P)                  T                  T�                   PUUU            PUU�                      �[    PUU     UUU�                      ��P�UUUU TUUUU�                      ��ZU�VUUUUU�_UUUU�                      ��ZU�VUUUUU�oUUUU�                      ��UU�VUUUUU��UUUU�                      ��UU�ZUUUUU��VVUU�                     ��UUUZUUUUUU�VZUU�                     ��UUUjUUUUuU�VZUU�                     ��UUUjUUUUuU�ZjUU�                     �jUUUjUUUUuU�ZjUUU                    ��jUUUjUUUU�U�jjUUU                    ��jUUUiUUUU�V��jUUU                    ��jUUUiUUUU�[��jUU�                    ��fUUUiUUUU�[��jUU�                    ��YUUUiUUUU�[��ZUUU                    ��YUUUiUUUU�[��ZUUU+                    ��YUUUieUUU����VU                      ��VUUUe�UUU����VU                       ��YUUUU�UUU����Z                       ��YUUUU�UUU����V                        ��iUUUU�VUUU���                       T��YUUUU�VUU���?                        U��UUUUU�VUUU��                       PU�jUUUUU�VUUUU)                        PUU@UUUU�ZU@U                         @  UUUU�V                                  UUU�                                   TUU�                                   PUUe                                   PUUU                                    PU                                                                                             �� �� �� �� �� ��  �  �  �  � 0  0  0  0  0  0  � 0 � 0 � 0 � 0  0  0  0  0  0  0 0 � 0 � 0 � 0 �  �  �  �  �  �  � 0  0  0  0  < < < < < < � � � � � � � � � � � � � � � � 0 00 00 00 0� � � � � � 0 00 00 00 000 00 00 00 00 00 �� 0�� 0�� 0�� 0� � � � � �  ? 0 ? 0 ? 0 ? 0   0   0   0   0   0   0   �   �   �   �   0   0   0   0   0   0   �   �   �   �   �   �   �   �   �   �               �?  �?  �?  �?  �?  �?  ��  ��  ��  �0  �  �  �  �  �  �        � �  �  �  �  �  �          �  �  �  �  �  �    0  0  0  0�00�00�00�00�00�0� �� �� �� 000000000000000000��0���0���0���0� �� �� �� �� �� � 0 0 0 0� �� �� �� �� �� � 0 0 0  0 � � � � � �     0 � � � � � � � � � � � � � � � � �                              �                                                    0   0   0 ,U�UUUUUUUUUUUUUUUUU�WUU�UUUUUUUUUUUU�?�_�WUUUUUUUUUUU� �? _UUUUUUUUUUU�    ��WUUUUUUUUUUU ���UUUUUUUUUUU= ?�?< UUUUUUUUUU�<��WUUUUUUUUU< �0�?0_UUUUUUUUU�������|UUUUUUUUUs������UUUUUUUUU]U �WUUUUUUUUUU�� �_UUUUUUUUUU�� �UUUUUUUUUU��  �WUUUUUUUUU 0�? �UUUUUUUuU �?  ��W�UUUUU������  ?�_UUUU?�_3 � 0<���UUUU� pU5����0��_UUU \U��0� �0<��UUU�WU�?? ����?_UU�WU��3��� � �pUUUUU���?�� � W�UUUU� �0 � 0 \�UUUU5   <� �  \5�WUUU ���0��\��WUUU�  ?� ��  pU?\UUU3 � � ?  �U\UUU= �  ��   _5UUU��U�p}<�p�UUUUUU=  _U� ���UUUUUU �UU��  W�UUUUUU5 _UUU < W�UUUUUU��UUUU� W�UUUUUUUUUUUU5� ��UUUUUUUUUUUU5�? ��UUUUUUUUUUUU�� ��UUUUUUUUUUUUUU? �UUUUUUUUUUUUU�  pUUUUUUUUUUUUUU5 \UUUUUUUUUUUUUU \UUUUUUUUUUUUUU WUUUUUUUUUUUUUU���UU0U�UUUUUUUUUUUUUUUUU�WUU�UUUUUUUUUUUU�?�_�WUUUUUUUUUUU� �? _UUUUUUUUUUU�    �_UUUUUUUUUUUU ���UUUUUUUUUUUU= ?�?UUUUUUUUUUU�<<�WUUUUUUUUUU< �0�UUUUUUUUUU�����?�UUUUUUUUUUs������WUUUUUUUUU]U��_UUUUUUUUUUU��  �UUUUUUUUUUU�� �UUUUUUUUUUU�� �WUUUUUUUUUU 0 �_UUUUUUUUuU �?UUUUUUUU�����? �UUUUUUUU?�_�  �WUUUUUUU� pU5< � �UUUUUUU \U� �� ��W�UUUUU�WU��0�  ?�_UUUU�WU���0<���UUUUUUU�0�?��0��_UUUUU���? �0<��UUUUU5   �?� ����?_UUUU   <�� � �pUUUU�  ��� � � W�UUUU3 �5�� �0 \�UUUU= W� � \5�WUUU��U ���\��WUUUUUU� ��  pU?\UUUUUU= ��?  �U\UUUUUU5  ��   _5UUUUUU��� <�p�UUUUUUU�_U� ���UUUUUUUUUU��  W�UUUUUUUUUU� < W�UUUUUUUUUUU� W�UUUUUUUUUUU�0� ��UUUUUUUUUUUU��? ��UUUUUUUUUUUU�� ��UUUUUUUUUUUU ? �UUUUUUUUUUU���  pUUUUUUUUUUUU�0 \UUUUUUUUUUUU� \UUUUUUUUUUUUU� WUUUUUUUUUUUUUU���UU)�UUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUU��WUU�UUUUUUUUUUUU� �_���UUUUUUUUUU  ���UUUUUUUUU � �?��UUUUUUUUU �?����WUUUUUUUU  ���\UUUUUUUU� �?��|UUUUUUUU�  ?0��?�UUUUUUUU5 <���?�WUUUUUUU5��<�� ?<�UUUUUUU5w���� 0���_UUUUU�UU�?� �����UUUUUUUU�0 �����WUUUUUU�0 �<��?|UUUUU��?0�?0?�WUUUW53<< <<<<��UU�\� <��<00��WU��3  � �0  ��\U5   W��?   �� |U����U��<  < WUU? _UUU=  � \��U� �UU��<� � p��U� �UU=� 0 � ��WUp�����?   _WU�_  �? ���� p�_UUU    ��� ��_UU��   ��W��  �sUU50   pUUU�? 0 �pUU5   _UUU�?  �pUU5 ��UUUUU=� �_UU���_UUUUUU���  WUUUUUUUUUUUUU�W \UUUUUUUUUUUUUUU5 pUUUUUUUUUUUUUUU� �UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUU�0�UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU�"�UUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUU��WUU�UUUUUUUUUUUU� �_���}UUUUUUUUU  ����WUUUUUUUU � �?�\UUUUUUU �?������_UUUUU  ��������WUUU� �?��?���?|UUU�  ?0��?���?�WUU5 <�����<��UU5��<�� ?�<<��WU5w���� 0�?00��\U�UU�?�  <3  �� |UUUU�0 � 0    WUUUU�0 �?   < \��UUU��?0�� � p��UUW53<� � ��W�\� <��? �  _W��3  �  ��? � p�_5   W� �� ��_����U�� ��  �sU? _U��< �� 0 �p� �UU=� ��U�?  �p� ���� pU�?� �_Up  � \UU=��  WU�_   ?�WUU��W \UU��    |UUUUUU5 pUU50   �WUUUUUU� �UU5   UUUUUUUU�UU5 ��UUUUUUUU�0�UU���_UUUUUUUUU��UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU�"UUUUUUUUUUU�UUUUUUUUUUUUUUU����WUUU�UUUUUUUU���?|UUU�_UUUUUU����?�WUU��WUU����<��UU� �_�����3<��WU  ��?���?0��\U � ���?� �� |U �?����?�  WU  ����? < \��U� �?���3� p��U�  ?0��< � ��W5 <�� ? 0 �  _W5��<�� 0   0 � p�_5w����� < � ��_�UU�? �� �  �sUU��0 ��?�� 0 �pUW5�0�����?  �p�\��?0<  ��?� �_��33�  U=��  W5  <  WU��W \��  ��?�UUUUU5 pU?   W���pUUUUU� �� ���U� \UUUUUU�� �_U��  WUUUUU�0�UpUU=��UUUUUU��U�_���pUUUUUU��UUU   ?\UUUUUUU�UUU    WUUUUUUUUUUU��   �UUUUUUUUUUUU50   UUUUUUUUUUUU5  �UUUUUUUUUUUUU5 �UUUUUUUUUUUUUU���_UUUUUUUUUUUU&UUUUUUUUUUUUU��WUUUUUUUUUUUUUUUU� �WUUUUUUUU]uUUUUU<  \UUUUUUUUs�UUUU���  pUUUU�WU��WUUU50  pUUUU�U5� WUUU� ��UUUU��W�? WUUU���0�UUUU= �   W�U�����WUUU    �����?����WUUU �?��0��� �WUUU ����0��� WUUU5 ��?������0��_UUU�   ?<��� \�_UUU5� <� � ? ? p�sUUU5\�� ?< � 0��pUUU5W5��<0���5�UUU�U��� < 0   �5�UUUUU� ?� ?< 00   ��UUUUW� <� ?< �� � ��WUU�\= 0��<�  0 0?WUU��  <�  ? �\UUU  ���� �  \UU�  ��00� �0 UU� �� � 0� < �UU��U�� ��U ��UUUU�� ����U� �WUUUU?�  ���UU? � \UUU� |? |� �UU� \UUU5? W��W� |UU�\��UUU��UUU�  _UU�\��U��? pUUU�  WUU�\��U= < \UUU�?�UU� WU�U ��WUUU�pUU5  WU}��  pUUU�  |UU�UUU50  _UUU _UU� �UUU5 �WUUU WUU3 pUUU5 |UUUU�WUU3 \UUU���WUUUU���UUU��WUUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �(          P@UUUUUUUUU                         P@UUUUUUUUU                         P@UUUUUUUUU ��             ���*     P@UUUUUUUUU `U                     P@UUUUUUUUU `U                     P@UUUUUUUUU `U            �
  ����  P@UUUUUUUUU `U            U	  `UUU  P@UUUUUUUUU `U            U	  `UUU  P@UUUUUUUUU `U            U���jUUU�* P@UUUUUUUUU `U            U	  `UUU  P@UUUUUUUUU `U            U	  `UUU  P@UUUUUUUUU ��            �
  ����  P@UUUUUUUUU                          P@UUUUUUUUU                          P@UUUUUUUUU                          P@UUUUUUUUU                     @U% P@UUUUUUUUU               ����      P@UUUUUUUUU               ���*      P@UUUUUUUUU               �����     P@UUUUUUUUU                 �*    P@UUUUUUUUU               TeU��� E! P@UUUUUUUUU               UeU�*   P@UUUUUUUUU               UeUU��"   P@UUUUUUUUU               UeUU��   P@UUUUUUUUU ��            UeUU�*  P@UUUUUUUUU               AeUU�*D% P@UUUUUUUUU                eTU��    P@UUUUUUUUU               AeUU��   P@UUUUUUUUU ��            UeUUU�    P@UUUUUUUUU `U            UeUUU�    P@UUUUUUUUU `U             e@� T% P@UUUUUUUUU `U            *e�J�   P@UUUUUUUUU `U            *e�J�   P@UUUUUUUUU `U            *e�JU�    P@UUUUUUUUU `U            Je�RU�   P@UUUUUUUUU `U            Je�RU� T! P@UUUUUUUUU ����   ���
  ��*e�JU�    P@UUUUUUUUU    �          e@U�    P@UUUUUUUUU    �         UeUU�    P@UUUUUUUUU    ����  ���* UeUU� @  P@UUUUUUUUU    �UUU  XUU% UeUU� T  P@UUUUUUUUU    �UUU  XUU% PeTU�    P@UUUUUUUUU ����UUU���ZUU��@ePU�    P@UUUUUUUUU    �UUU  XUU% PeTU�    P@UUUUUUUUU    �UUU  XUU%UeUUU�    P@UUUUUUUUU    ����  ���*�������    P@UUUUUUUUU               UUUU���* P@UUUUUUUUU               UUUU(    P@UUUUUUUUU                UUUU     P@UUUUUUUUU  QU      EU UUUU     P@UUUUUUUUU      ����  @  UUUU     P@UUUUUUUUU     ����* @  UUUU     P@UUUUUUUUU     ������ @ UUUU     P@UUUUUUUUU     ��  �*@  UUUU     P@UUUUUUUUU `T �*TeU��� EUUUUUUUUUUU@UUUUUUUUU    ��BUeU�*@UUUUUUUUUUU@UUUUUUUUU    �*TUeUU��"@ UUUU       @UUUUUUUUU   ��BUUeUU��@ UUUU       @UUUUUUUUU   ��TUUeUU�* UUUU       @UUUUUUUUU `P�*UUAeUU�*BUUUUUUUUUUUUUUUUUUUUUU   �JUU eTU��UUUUUUUUUUUUUUUUUUUUUU   �JUUAeUU�� UUUUUUUUUUUUUUUUUUUUUU   �RUUUeUUU� UUUUUUUUUUUUUUUUUUUUUU   �VUUUeUUU�  UUUUUUUUUUUUUUUUUUUUUU `U�RA e@�HUUUUUUUUUUUUUUUUUUUUUU  @�V �*e�J� UUUUUUUUUUUUUUUUUUUUUU   �VA�*e�J� UUUUUUUUUUUUUUUUUUUUUU  @�RU�*e�JU� UUUUUUUUUUUUUUUUUUUUUU   �VUJe�RU�UUUUUUUUUUUUUUUUUUUUUU `U�VUJe�RU�HUUUUUUUUUUUUUUUUUUUUUU   �RU�*e�JU�UUUUUUUUUUUUUUUUUUUUUU   �VU e@U�UUUUUUUUUUUUUUUUUUUUUU   �VAUUeUU�UUUUUUUUUUUUUUUUUUUUUU   �R UUeUU� UUUUUUUUUUUUUUUUUUUUUU  T�VAUUeUU�HUUUUUUUUUUUUUUUUUUUUUU   �VUUPeTU� UUUUUUUUUUUUUUUUUUUUUU   �RU@ePU� UUUUUUUUUUUUUUUUUUUUUU   �VUUPeTU� UUUUUUUUUUUUUUUUUUUUUU   �VUUUeUUU�  UUUUUUUUUUUUUUUUUUUUUU   ����������� UUUUUUUUUUUUUUUUUUUUUU ���BUUUUUUU���UUUUUUUUUUUUUUUUUUUUUU   �@UUUUUUU(  UUUUUUUUUUUUUUUUUUUUUU    @UUUUU   UUUUUUUUUUUUUUUUUUUUUU    @UUUUU   UUUUUUUUUUUUUUUUUUUUUU    @UUUUU           UUUUUUUUUUUUUU    @UUUUU           UUUUUUUUUUUUUU    @UUUUU           UUUUUUUUUUUUUU    @UUUUU   UUUUUUU UUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUU UUUUUUUUUUUUUUTUUUUUUUUUUUUUU      P UUUUUUUUUUUUUU       UUUUU          P UUUUUUUUUUUUUU       UUUUU          P UUUUUUUUUUUUUU       UUUUU          P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ���* P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU �    P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU �    P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��    P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�    P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�    P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��  P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�   P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�   P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��   P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   �* P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���  P UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU     P UUUUUUUUUUUUUUUU��VUUUUUUUUUUUUU     P UUUUUUUUUUUUUUUU�	VUUUUUUUUUUUUU   �* P UUUUUUUUUUUUUUUU��ZUUUUUUUUUUUU   V% P UUUUUUUUUUUUUUU�"�XUUUUUUUUUUUU   V% P UUUUUUUUUUUUUUU�*��UUUUUUUUUUUU   V% P UUUUUUUUUUUUUUUU���UUUUUUUUUUUU   V% P UUUUUUUUUUUUUUUU	��UUU             V% P UUUUUUUUUUUUUUUU���UUU             V% P UUUUUUUUUUUUUUUU� �UUU             V% P UUUUUUUUUUUUUUUU)(�UUU@UUUUUUUU   V% P UUUUUUUUUUUUUUUU�
jUUU@UUUUUUUU   �* P UUUUUUUUUUUUUUU���VUUU@             P UUUUUUUUUUUUUUU� ��VUU@             P UUUUUUUUUUUUUUU��� ZUU@             P UUUUUUUUUUUUUUU)��*XUU@             P UUUUUUUUUUUUUU���*��VU@ ��
  �*     P UUUUUUUUUUUUUU�)(��VU@           P UUUUUUUUUUUUUU�
 ���VU@           P UUUUUUUUUUUUUUb��UU@  ���*      P UUUUUUUUUUUUUUb��
��UU@  XUU%      P UUUUUUUUUUUUUUb��
��UU@  XUU%      P UUUUUUUUUUUUU�b
�Z�UU@ �ZUU%      P UUUUUUUUUUUUU�`
 �V�UU@ �XUU%    �* P UUUUUUUUUUUUU�h) �U�UU@ �XUU%      P UUUUUUUUUUUUU�X� hUbUU@ ����*      P UUUUUUUUUUUUU�X��ZUbUU@ �          P UUUUUUUUUUUUU�h��X��UU@ �����*   �* P UUUUUUUUUUUUU%`��Z��UU@ ��        V% P UUUUUUUUUUUUU�jUUU��UU@ �        V% P               �   �� @ �        V% P               �   �  @ �        V% P                       @ ��        V% PUUUUUUUUUUUUUUUUUUUUUUUU X�        V% PUUUUUUUUUUUUUUUUUUUUUUUU X�        V%                            X�        V%                            X�        ���*  ����  ���*  ����  ����X�             �          �       �X�     �(Uj����V�V�i��jUj�RUUUUUUUUPUUUUUUUUUUU�����Z��ZiZ�U��ZU��  TUUUUUPUUUUUUUUUUUj��e�V�UiUZi�U�Z��PUUPUUUUU @UUUUUUUUUU�UeU�Rj���ZieU�V��
TUU TUUUU  UUUUUUUU�UYV�BZi��iYe��U��BUUUUUPUUUUUEPUUUUUUU�V�ZU
ZYe����j��( PUUUUUAUUUUUTTUUUUUUUVfi�*i�Z���UUj�*UUUUUU UUUUUTUTUUUUUU@VYe�*dU�*�Vj�V�
UUUUUUUUPUUUUPUPUUUUUUHZ�Z���Zj �Z�V%�@UUUUUUUUUAUUUUAUAUUUUUUJ�V�B��Z�Z�*TUUUUUUUUUEUUUUTEUUUUUU
@���
U�Z�Ui�UUUUUUUUUUUUUUUPEUUUUUU(
 P *(`UeU���PUUUUUUUUUU TUUUQEUUUUUU�*��
��jJYeU�
TUUUU PUUUUTUUUQUUUUUUU ���*@��RIY�U�@UUUUU�BUUUU TUUQUUUUUUU��
U�P	e�U�PUUU  �
  TUUTUUQUUUUUUU �BUU�R)�j��BUUU�*����PUUPUUQUUUUUUUUU PUU�JTeJUU�
�*�RUUQUUUUUUUUUUUUTUUU*P���JUU�J!@U� RUUAUUUUUUUUUUUUTUUU�U��@UU�@ UU�TUU UUUUUUUUUUUTUUUU*  �*TUU�X�UU�V�UUEUTUUUUUUUUUUUUUUU���� UUU�X�UU V�TUEUUUUUUUUUUUUUUUT�
�*TUUU�X�ZU jRTUEUTUUUUUUUUUUUUUEU@
UUUU�XhU�RTUEUUPUUUUUUUUUUUUUAUUU@UUUU!X`UA�
RTUEUU@UUUUUUUUTUUUQUUUUUUUUU ZUhUQ�
RTUEUUUEUUUUUUUUUTUUUQUUUUUUUUU(VUhUQ�RTUUUUEUUUUUUUUU@UUUQUUUUUUUU(VU�UQ�RTUUUUUUUUUUUUUDUUUQUUUUUUUU�VU�UQ��RTUUUU TUUUUUUUUUU@UUUUUUU�UUhUU��BUUUUUUPUUUUUUUUUUEUUUUUUU��UUhUU��
UUTUUUQUUUUUUUTUUEUUUUUUU�jUUhUU��*TUUPUUUAUUUUUUUTTUUEUUUUUUU�ZUU�UU���TUUQUUUEUUUUUUUTTUUEPUUUUUU�ZUU�UU�PUUPUUPEUUUUUUTTUUEUAUUUUU�ZUU�UU�RUU@UUUQUUUUUUUUTUUEUEUUUUU�YUU�UU�VRUUUUUQUUUUUUUUTUUUEUUUUU�YUU�UU�jBUTUUQUUUUUUUTPUUTUUZiUU��YUU�VU`JUUPUUQUUUUUUUUTAUUUTUU�ZUU�UUV�VjUZa(UEUQUUQUUUUUUUUTEUUUPUU�UUU�UU�jU����`(UEUAUUQUUUUUUUUTUUUUQUUUUUhU��UeU����a UEUEUUUUUUUUUUPUUUUUUUUUZ��VU�UU�*�a!UEUEUUUUUUUUUUQUUUUTUUUU!V%ZU�VZU�"�a!UEUEUUEUUUUUUUQUUUUETUUZY�V�UUiU�UU��!UEUUUEUUUUUUUEAUUUUQTUU�Z�U�VUUQVUj��!UQUUUEUUUUUUPEUUUUPTUU��U�U�j��iUi��%UQUUUEUUUUUUAUEUUUUTTUUUjU�Uej��fUi��&UQUUUUUUUUUUQUEUUUTPUUUjU�VYVeU�Uj��&UQUUUUUUUUUUQUEUUUUQU �ZU�UVUUUUV�U�
UQUUUUUUUUUUUTUEUUUEUQU*�ZU�UZUQ�V�U�
UQUUUUUUUUUUUTUEUUUAUQU��VU��ij���Y�UU
UQUUUUUUUUUUTUEUUUQUAU���VUi��i��iZ�UU�TUUUUUUUUUUUUTUTUUQUEU� �VUj�QeQY�VU�TQUUUUUUUUUUUTUEPUUPUEU!D"VUj�UUUUUY�VU�PQUUUUUUUUUUTUEQUUTUEU E�UUb�UUUUUY%VU�RQUUUUUUUUUUUUEAUUTUE(U�VUY�QUeUY�UU�RUUUUUUUUUUUUUEEUUTUE
UYZU���i��iZ�U��RUUUUUUUUUUUUUEUUUTUE�B�U�U�Vfj��fVjU��PEUUUUUUUUUUUUEUUUPU�@�ViU�ZZUQ��ZU��TUUUUUUUUUUUUUEUUUQU�D�ViUejYUUU��fU��TUUZiUUUUUUUEUUEUUUAU�T�V�UU�ie�e��UUi�PUU�ZUUUUUUUEUUEUUUEU�T�V�YU��i��ijV�i�RUU�UUUUUUUUQUUEUUUEU�T�V�VU�ZEQ�ZUU�URUUUUUUUUUUUQUU@UUUEUU T�V�ZUUjjU��VU�ZURUUUUUUUUUUUUUUDUUUAUU T�ZU��Z���Zi��*VURi�UUUUUUUUUUUUTUUQUU U�ZU���ViU�U���UUR�jUUUUUUUUUEUUTTUUQUU(U�ZUUU�Z��i��VUUURUVUUUUUUUUUUUTTUUQU(U�ZUUUU�UFVYUUUUURUUUUUUUUUUUUUUTUUUU*U�ZUUUU�VUUZUUUUURUUUUUUUUUUUUUUTUUUU&U�ZU����QTY���VURUUUUUUUUUUUUUEUUUUUU&U�Ze������i���*fUBUUUUUUUUUUUUUEUUUUUU&U�Z�ZUUUjU�VUU�ZUJUU PUUUUUUUUEUUUUUUV��Z�ZUUi��Z�UU�ZUJZi��BUUUUUUUUEUUUUUUV��Z�VU�jiU���UUZ�J�Z� JUUUUUUUUEUUUUUUV��Z�V��VVUUV�ZUjUI�U!HUUUUUUUUEUUUUUU�V��Z�U&V�jU�ZUbViVIUUaTHUUUUUUUUEUUUUUU�T��Z�U�Ue�V
fU�U�UIUUaTUUUUUUUUE@UUUUU�T��ZiUiUe� fU�U�UJUU`�*UUUUUUUU@UUUUUaT��VbejUe	V�eU�f%VIUUh� UUUUUUUUUUUUU`TY�VZ�ZUe�U�eU�Z�VJUX� UUUUUUUUAUUUUUhTY��Z�fUeU�UeUeZ�Z*UZ� TUUUUUUUAUUUUhP���Z�UU�iU�iUUY�V*UZ��TUUUUUUUPTUUjP��Vi%VU�Z��ZUUb�U&U�j��TUUUUUUPTUU�VQ��Vi��UUYV�UU�j�U&UhZ��PUUUUUUTDPUU�PU��Uf���Ui��U��ZeV&UXZU�RUUUUUUT@@UU�TU��U�U��j��j��jUi�&�jU�PUUUUUPT P U�T��jY�UUUUUUUUUUUY�&�jU�RUUUUUP      �U��VZ�VUUUUUUUUUUZ���jUUUUUU@ @ T�U���VUVUUUUUUUUUUV���jU*PUUUU @UUUUU�U��fUUVUUUUUUUUUUV�U�jU�RUUUU  UUUUU�U��f�UU�UUUUUUUU�U�U
��URUUUUUUUUUUU�U��feUU�UU���V�U�U�U	��URUUUUUUUUUUU�U��feUU�UU���Z�UeU�U��URUUUUUUUUUUUVU��eUUU���Z����UaU�U(��URUUUUUUUUUUUV���iUUU�������jU`U�U���ERUUUUUUUUUUU�V��ZiUUU��Y����jUaU�U���URUUUUUUUUUUU�U���ZUUUU�������U`U�V����URUUUUUUUUU�U�V���YUUUU�����j�VeU�Va���URUUUUUUUUU�U`V���YUUUU���j���VUU�Ua���UUUUUUUUUU�VhV���YUUUUf��j���VVU�U����U*PUUUUUUUY�VXU�jYYUUUUf������ZVU�U����U�RUUUUUUUj�ZXU�jZUUUUUe����j�ZVU�Ua���URUUUUUU�j�ZXU��YUUUUUi��Z�Z��VU�Ua���ZUJBU�UUUU���*X���iUUUU�Z��jV��jUU�Ve��XUYBU�UUUU����Z���eUUUUU���jU��jUUUVeY�XUYB��UUU�����Z���eUVUU����jU��jUUVei�XUYJ��Z����UU�V�V�eUVUU�����Y���UUVee�XUY	��ZUUUUU��UU�jeUVUUU��������UUVUe�*VUU���jUUU����*aeUVUUU��������jUVUe�(VUY���� U  
    `�UVUUe��������UUUVU��(UUUY���i�UVUUe��������jUUVU�V�UUUY���          XUUVUUe��������eUUVU�U�UUY����ZUZUUe��������UUVU�T�VUU	             jU�UUe��������UU�VU�T��TUIUU�U�UUe��������UU�UU�Q�����JUU           ���UUe�"
  ���iU�UU�UaU��*@UU�ZU�  �ZU�UU�UiUUUUUU              ��*        �jUU���ZUUUUUUU   �jU�UUUUUUUUUU                          ����UUUUUUUUUU    QUUUUUUUUUUUU                           UQUUUUUUUUU      PUUUUUUUU                            UUUUUUUU       PUUUUUUU                            QUUUUUU         TUUUUU                            QUUUUU        UUUUU                              UUUU          QUUU                                UU           QU                                @U                             Q    @                            @                      @                                                                                                           @                                                                                                                                      @       (	UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUU\UUUUU�� pUUUUU=< pUUUUU� �U�U ���?�W ��U �_� ���?�p���� �U?��_ 0W �W50 W �U��0�U���U� �0 �}U�� ��U�� \�0p�UW\�U �U5 WuU�W��\]U5p}� ?pWU�_�70�UUUU�� 0WUUU3 WUUU �_UUU� ��?pUUUU <pUUUU���pUUUU UUUU�  0\UUUU� 0�WUUUU5 0 UUUU0� WUUUU \UUUU \UUUU����_&UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUUUUUUUU_UUUUUU_UUUUUU_UUUUUU_U���WU_U���_�_U���WU���s�WU�p�WU�����W�<  <�W�<<<<�W�<  <�U�<�<�U��0��UU����UU���UU���_�UU5  \}UU���}U����U�����U�����U����?pU3  0pU����\U<���_U���UU�p5 WUUp��UUUpUUUUU�_UUUU&UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUUUUUUUU_UUUUUU_UUUUUU_U���WU_U���_U_U���_U���s�WU�p�WU�����W�<  <�W�<<<<�W�<  <�W�<�<�U��0��UU����UU���UU���_�UU=  |�UU���}UU���}U�����U�����U����?pU3  0pU����\U����_U��=�WU��5�WUUp5�UUU�_5�UUUUU�UU&UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUUUUUUUU_UUUUUU_UUUUUU_U���WU_U���_U_U����_U��p�WU�  �WU�����W����?�W����?�W����?�W����?�U������UU�����UU����UU5��\�UU�  _�UU���}UU���}U�����U�����U����?pU3�0pU����\U���_U���UU� p5 WUUp��UUUpUUUUU�_UUUU&UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUU}UUUUUUUUUUUU_UUUUUU_UUUUUU_U���WU_U���_U_U����_U��p�WU�  �WU�����W����?�W����?�W����?�W����?�U������UU�����UU����UU5��\�UU�  _�UU���}UU����}U��<��U�����U����?pU3�0pU����\U����_U��=�UU��5 WUUp5�UUU�_5�UUUUU�UU2      @� �       �@�� �  �    @���� ��!@    @� �" !@    @��"�� !B    Т��.2)�    Q����"")B    �B�@�"")B    9F��  �"")B    D� ����"")B    @�� ��.2)B    @� �@"")B    @� �� ��    @����A    AP����� @@    � �  D   @                     ��  @!   ���,� ���  ���� @H�  �����@� B*� ���D���@@0 ��D"$( �10 ����%( ȃ!����$�r ��H����$�  �  @�@D�"b �� � ��F#t�!��  � B!��D� ��  � B!@ D ���  �"B! D ���  ������D� �0�  �     D                   D �@�@      .� D �@�B      B D�@��      N� ����@      �[B�@��      ��YB�@�@      p YB�B����  O� _r��� ��  A �B�`����  AR XB�����  M� IB�Ш�      A� �B�Q�      A uӋG��      ��"b�B�       �� "@�      �  �  @�      v         � �       �����"�  ` !����p   ��b@� @ @    A � @ "0 � ����n���0 �"���R"  �"@� B"  @�!��� B"� @�!p�N� @��b@��D"A�  ���@BO�H/�  ��d�@�@0�  @D�@@,�H��   ( ADF�     �H   A�                    �        @ ��� ���   � ���""��   B" �""��J� @�""0h!b"�������d0D&^�Ow�$D�$@ 8� 	� �!L� ��	@ @!D������P p�Db  ��@�   @@L�B�� �d0`P  @ D�	@� H�  @D@
 �� D  L L� A��p�� B  C D �   @p A                  �  ��    ����(��    @����@�P@P��  ���B @���@P@  @�B��"�  )�O�0@�B���!  �@`@�B���"���`DD�󀀌��H�@`�D���@�   O�0�B� ��(� �@  B� ���@�,�O�  A� �� @�PA  @����@���!  @�@pBEt!  @����.�" ,��  ��@ @  �                   �     �  �� �    ���Q ��    ��  R� B  �� B  ���!B"�!B  �@��b0"��b ��P�1R0"�1R���B�!B"�!B  �R�!B "�!B  �R�aB "�aB  �Q��B "���B  �A� B  �r� B ���$B  "�$B��NԄB   �B  "%��B�   ��B�  � B   � B                	@       � �@	@      ��@����    ���@	@ ��   ��@O�	@   � � HA��.2	 0�"�hA(""	 ��0����^�""�� ��RJ@��""��  ��RJB��""   ��RN���.2	   ��BHB��""	@   ���"HB�� ��   �P�"D���H�  � �DA@ *��  �`�AC@        �@@�@@                              �     �   !@�!��  �!  !@L�""   �!B! "" @ ` 0)�""" ��A 0)B��"" ?v��")B� ""   �� )B�!"" @ � )B��""� ` )B� !� @ H�  )B� � @ D  �  @@ N�  �A�0��@ D  @@�� @p @   @�    @                              .��            BH            BH            Oq            �H0          rD`          NBa`          B1AA`          BQ��0          OQD            I             ��            B��            Q��            ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �(UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                                        @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                            T                          P      @TP                      P Q@    A TPET                    U P@Q     T                       P P @  P   @                  P @   @@AU @U  T                  U U  @  E @UP                @   U@ TQDU                  T PEQTA@P  APP P@                A  AA@   P  T     @U           PT@  U  @P  QT   @D U P      T  AU   @     PQP     T@U UDU         @EA @U   @        P@@      UT      PA@U        @        @ U       UU          T T  @E      TU                     PP@ T                            TP@EDQPP P                                                            @Q@ PQ@                           P  UP E                                                                 TQ  @ T                                  T                                    PU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               P                                     @@                                   P                                     @@                                   D T                                   Q                                     @                                     @@PD                                 AE              �������������      T                             �    @UTPDP              �W@T@T�T@	X    P@E             �UUUUUUUUU�UUU	   T                �VUUUUUUUUUUUU	   @EQ   @              �Z��Z��Z��Z��Z	   @U                �j��j��j��j��j
   PE                 ��*��*��*��*�   U  P @               ��
����
���   @TU   U                `EEEUTTTEEEU$    U                     `UEUUUTUUEUU%  PU                      UUQPUUQ%  PPT @                   TT@ATT@%  P P                  T@Q@T@Q�������                  UQQQUQQ)      AU                  UUUQUUUUUQZ``}                  TEU@UTTEU@VUUUY�Ue                   `PPAPDZUUUUUUeAP                 `EPPEUj�Vj�Vj%T        @        `EEEUTTTEEEU�������)          P        `UEUUUTUUEUU�������Z            ������/UUQPUUQ�*�*�V         P �     �TT@ATT@ATT�UA          �PP�T@Q@T@Q@T@�UQ       DT@aUUUeUYUUQQQUQQQUQ�U       DPD@�UUUUUUUVUUQUUUUUQUUUUU�U       A�Vj�Vj�VVEU@UTTEU@UTTEU�E       @PT@��������RPAPPAP�������   P��������EPPEPPE�      <     EEj�Fj�ZjEEEUTTTEEEUTTTEEEiT�T��    PPQYAUUUTUUEUUUTUUEUUUTUUEUYU�UUeU�   @XUQQUUQQUUQQUUiUUUUUU�   D TUYT@ATT@ATT@ATT��Z��Z��   D UT@Q@T@Q@T@Q@T@��j��j��   TQU UQQQUQQQUQQQUQ�*��*��*   TXUUQUUUUUQUUUUUQUUUUU�
��
��
   D XEUDUTETEUDUTETEUDUTETEUUEUTEU   PQQ XPAPPAPPAPPP    UT  EPPEPPEPPEPPE	    P  HEEUTTTEEEUTTTEEEUTTTEEEUTTTEEE	    PU  XEUUUTUUEUUUTUUEUUUTUUEUUUTUUEU	VVRRVVRRVVRRVVRRVV
����������������������������������������aaaaaaaaeaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaiYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTUUUUUUUUUUUU�VUUUUUUUUUUUUUUUUUUU�UUUUU�ZQQQQQ��RQQQ�RQQQQQQQQQQQQQQQQQjQ�RQQQQ�ZTTTTT��jTTT�VTTTTTTTTTTTTTTT���Z�ZTTTT�ZUUUUUjU�ZU��UUUUUUUUUUUUUUUUeUUe�VUUUU�ZEEeE�JE�jE��EEEEEEEEEEEEEE�EIEE��EEEE��FQQ�Q�RQ��Q�jQQQQQQQQQQQQQQ�QQQQ�jQQQQ��QUU�U�UU��VU�jUUUUUUUUUUUUU�VUUUU�UUU��VU�)�������EE�FjEE�Ej�FEFEEEEEEEEEEE��FEEEEE���j�FEUU�VZUUjU��UUYUUUUUUUUUUU��VUUUUUU��jUZUTT��VTTZTTTTTTTTTTTTTTTTT�j��TTTTTT�jTZT�����UU��UUUVUUUUUUUUUUUUUUUUUU�UUiUUUUU�ZUZUQQ�jQQQQQQQQQQQQQQQQQQQQQ�jQQ�QQQQQ�RQjQTT�ZTTTTTTTTTTTTTTTTTTTTT�VTT�TTTTTTTTjTU��UUUUUUUUUUUUUUUUUUUUUU�UUU�VUUUUUUUiZ��JEEEEEEEEEEEEEEEEEEEEEEiEEEEFEEEEEEE���jQQQQQQQQQQQQQQQQQQQQQQQjQQQQ�RQQQQQQ��UUUUUUUUUUUUUUUUUUUUUUUUUZUU�U�ZUUUUUU�Z�����EEEEEEEEEEEEEEEEEEEEEEE��FEEE�EEEEEEEE�FUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUU�VTTTTTTTTTTTTTTTTTTTTTT��ZTTTTTTTTTTTTT�T��UUUUUUUUUUUUUUUUUUUUUUjUUUUUUUUUUUUUUU�U�(UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                                        @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                            T                          P      @TP                      P Q@    A TPET                    U P@Q     T                       P P @  P   @                  P @   @@AU @U  T                  U U  @  E @UP                @   U@ TQDU                  T PEQTA@P  APP P@                A  AA@   P  T     @U           PT@  U  @P  QT   @D U P      T  AU   @     PQP     T@U UDU         @EA @U   @        P@@      UT      PA@U        @        @ U       UU          T T  @E      TU                     PP@ T                            TP@EDQPP P                                                            @Q@ PQ@                           P  UP E                                                                 TQ  @ T                                  T                                    PU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ����������������������������������������aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTUUUUUUUUUUUU�VUUUUUUUUUUUUUUUUUUU�UUUUU�ZQQQQQ��RQQQ�RQQQQQQQQQQQQQQQQQjQ�RQQQQ�ZTTTTT��jTTT�VTTTTTTTTTTTTTTT���Z�ZTTTT�ZUUUUUjU�ZU��UUUUUUUUUUUUUUUUeUUe�VUUUU�ZEEeE�JE�jE��EEEEEEEEEEEEEE�EIEE��EEEE��FQQ�Q�RQ��Q�jQQQQQQQQQQQQQQ�QQQQ�jQQQQ��QUU�U�UU��VU�jUUUUUUUUUUUUU�VUUUU�UUU��VU�)�������EE�FjEE�Ej�FEFEEEEEEEEEEE��FEEEEE���j�FEUU�VZUUjU��UUYUUUUUUUUUUU��VUUUUUU��jUZUTT��VTTZTTTTTTTTTTTTTTTTT�j��TTTTTT�jTZT�����UU��UUUVUUUUUUUUUUUUUUUUUU�UUiUUUUU�ZUZUQQ�jQQQQQQQQQQQQQQQQQQQQQ�jQQ�QQQQQ�RQjQTT�ZTTTTTTTTTTTTTTTTTTTTT�VTT�TTTTTTTTjTU��UUUUUUUUUUUUUUUUUUUUUU�UUU�VUUUUUUUiZ��JEEEEEEEEEEEEEEEEEEEEEEiEEEEFEEEEEEE���jQQQQQQQQQQQQQQQQQQQQQQQjQQQQ�RQQQQQQ��UUUUUUUUUUUUUUUUUUUUUUUUUZUU�U�ZUUUUUU�Z�����EEEEEEEEEEEEEEEEEEEEEEE��FEEE�EEEEEEEE�FUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUU�VTTTTTTTTTTTTTTTTTTTTTT��ZTTTTTTTTTTTTT�T��UUUUUUUUUUUUUUUUUUUUUUjUUUUUUUUUUUUUUU�U U�UUUUU��UUUU��WUUU�\UUU=�|UUU���WUU 0 WUU � WUU   WUU  �UUU=  pU_U�  _�sU�?�W=�UU����UU����U����_U��?�WU���0 WU���� WU����U����W?��_���� �U��? �U�����U��W��UU W�pU� �U�_UU�UUUU� �UUUU��UUUUU�UUU UUUUUUUUUUUUUUU��UUUUU��WUUUU3?\UUU�30pUUU�0�UUU5 3�_UU � \UU 0\UU=   \UU5  �WUU�  �UUU� |UUUU _UUU���WUUU�?WUUU��<_UUU��3|UUU�?��UUU�?�WUU�??_UU�??\UU���\UU��_U����pU��?_U��? �pU�   0pU�  <pUU  pUU=  �_U$UUUUUUUUUWUUUUUU�uUUUUUUu]UUUUUU]�UUUUUU�u]�WUUU�]�_UUUU���pUUUU}���UUUU��<�WUUU� UUU5  pUUU5   pUUU�   pUUU�  �_UUU�  WUUUU ��WUUU= |�|UUU�?���UUU����UUU�����UUU�����UUU����UUU�����UUU��?sUUU���?UUU���?\UUU����UU������UUU���? WUU5 p�_UU5 p50pUU���UU� \��WUU��\U�UUU�_U}U$UUU��UUUUU�UUUUUU��UUUUU�UUUUUU��UUU���UUUU����UUU3?\WUU�30pWUU�0�UUU5 �_UU �\UU   \UU=   \UU5  �WUU�  �UUU� |WUUU _WUU���WWUU���_UU��?<\UU�?�3_UU���WUU���WUU����WUU��WUU���_UU�����UU�����UU���pUU�=<pUU��|UU���_UUpU�WUUsUUUUU�UUUU U��UUUUUU��WUUUUU3?\UUUU�30pUUUU�0�UU�W5 �_Uu] �\U�u   \U]�=   \U]5  �WU�u�  �U�_W� |U�u]U _U}�U���WU_UW��_�WUU��?|uUUU����UUU���pUUU���\UUU���pUUU�?��_UUU���\UUU����\UUU����_UUU����WUUU���UUUU ? _UUU�� |UUU�����UUU�U�UUUW�UUU��W�UUU$�UUUUUu]UUUU_�UUUU�uUUUU�]�_UU��?|UU�?��UUU?WUU� _UU00�U�  <�U�   �U�  �UU �UU  \UU= �WUU� �|UU�?<�UU����W��� �_�����������?������WU��?�\U����\U����sU����sU����_UU 0\UU�|UU��pUU<0\UU��WUU=3�UUU�?�UU UU�WUU�UU�_UUW_U��pU�UU���U��W��<�W�_U� u�U5  p�WU5   p]}U�   p]UU�  �__UU�  WWUUU �UWUUU= |�UUUU�?_�UUU��3|�UUU����uUUU���?wUUU�� �UUU�����UUU����sUUU�����UUU����UUU���WUUU����WUUU����WUUU���?\UUUU �|UUU���pUUU� <|UUU�3��_UUUU?0 _UUUU�?�WUUU U�UUUUUU��UUUUU��WUUUU�\UUUU=�|UUUU���WUUU � WU�U   WU�_   WU}}  �UU��=  pU�__�  _U�}u��WU��U���UU�WW���WU__U���W�WuU�� �UUU����}UUU���?_UUU���?\UUU���_UUU��0\UUU����_UUU���WUUU����_UUU���|UUU � pUUU���UUU��U��UUU\���WUUpU WUU�U��WUU UU�WU�WU�_U]UU��pU�WU���U]U��<�W�W� _U5  p�W5   pWU�   pWU�  �_WU�  �WUU ��UUU= |�UUU�?_�UU��3\�UU���p�UU�?��UU�����WU��?<WU��<�WU����UU���UU�?���UU�����UU�����UU� 0\UUU��pUU�� �pUU� 0\UU� �WUUU��UUUU���UUU UU��UU�_UU��WUuUUU3?\U�_U�30pU}UU�0�U�_U5 �_}UU �\�_U   \]UU=   \]UU5  �W]UU�  �U]UU� |�UUU _?pUU������U��??��U���0��U�����wU�����wU�?�?<�uU���0|uU�����puU}����puUU����|uUU����UUU�?��pUU� ��UU�  p�UU |�UU�_��WU�U�UU�WU�UU�UUU��WU UU��U�UU��W��UU3?\�U�30p��U�0��U5 ���U ��U   ��U=   �UU5  ��UU�  ��UU� |uUUU _uUU���WuUU��WuU���0�uU������W����<W������U�?���W�����W����uU���0�uU����|]UU��_]UU�p]UU 0�]UU� ��UUU� ��UUU���WUUU \UU����_U UU�WU��U�_U�UU��pU��U���U�U��<�W��� �U5  p��5   puU�   puU�  �_uU�  WuUU �UuUU= |UuUU�?_UuU��3�_uU������U��?��U�?���sU��3��U������U����uU��?�uU=��?suU���?uUU����uUU� �wUU� wUU?�=�_U��5�|U� p�pUUsUsUU�|U�\U U�UUUUU��UU�U��WUWW�\U�U=�|UWW�����U � �WW   ��U   ��W  ��UU=  p�UU�  _�UU��W�UU���UuUU�?_uUU��|uUU=�3�wUU����WU��<WU����UU���0WU?�0�WU� �0wUU�0�3wUU����wUU�  wUU�  �]UU�  �UUUU��|UUUU�pUUUU��UUUU���UUU U��UUUUU��WUUUU3?\UUU�30pU�U�0�U]W5 �_] �\�U   �_W=   �uU5  ���U�  ��]U� |uuUU _}UU���W]UU��__UU��?|WUU����UU��0pUU���\UU���pUU�?��UU���\UU����_UU����UUU����WUU5��_UU � |UU= � �UU��W�?WU5 W WU��\=�WU��_��UUU���WUU���_�U����U��p�U�  �U���������?�����?w����?w����?w�����wU����uU���uU5��\uU�  _]U���]U���]�����W�����_����?p3�0p����\����_��=�u��5 WUp5�UU�_5�UUUU�U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �(                                                                                                                      @                                      PU                                      U                                      PQ                                      PU                                      PU                                      TU                                      DU                                      TU                                      T                                      TU                                      TU                                      TU                                      UU                                      UU                                     @UU                                       P                                     PUA                                                                            T             @                                    P @                                    P @U                                    PPU                                    PE                                    PE                                   UPA                                  UTU                                  UTQEE                                 @UUTUUU                             U TUUUUUU                            UUUUUUUUUU                          @UUUUUUUUUUUUU                              TUUUUUUUUU                       @U   PUUUUUUUUU                         TU  TUUUUUUUU                                TUUU                               U  @EUUU                            U @U DUU@UU                           P  TT  T                                                                      T   P                               T @ U                                    UU                                                                                                                                                                                                    P                                       @U                                        UU         P                                       P                                      T                                     T                                     T                                     U                                   @Q U                                   @A U                                   PE@                                  PUAUP                                 PUAUT                                 TUEUUU                                @UUEUUUUU                              UUUUU PU                                PUUP                                PUUU U                               @@     PU                                                                                                         P       @UU                          @      P                               P     T                                     @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 T                                                                           @P                                   �PP                                  �
��                                 @�j�V�                                T������*                               @U�V�����                               PU�VU���V            U                 UU�VU��UU          @                PUU�UUUUUU)          P                 TUUiUUUUUU��        T T               PUUU�UUUUUUU��       de              PUUUU�VUUUUUU���      �Ui              �VUUUUUUU��UU�����    ����
             �ZUUUUUUUU�jUU������ ��j���     �
    ��jUUUUUUUU��UU��������������   ���*   UUUUUUUUUUUU��UU����Z�Z��j����jU�jU������(                                                                                                                                                                                                                                                 @                                  P P                                  T T                                  PP T                                   T                                  UU DU                                  UUU UU                                 UUUEQU                                 UUUUUU                                UUUUUUUT                                UUUUUUUU                               UUUUUUUUU                               UUUTUUUUU                              UUTU  TUUU                                TQUU                                 UUUP@UUUU                              @U                                     U@                                  @U  U                                   PUA                                      U                                      @                                                                                                                                                                                                                               @                                      @                                      P                                     P                                     P                                    T T                                    ET                                    TQ                                   @TP                                  @UUU@                                 @UUTQ                                 PUUUUU                                 UUUUUUU                              TUUUU@UU                                @UUU@                               @UTU TT                                     @U                 @                                    P @                                    P @U               UU                 PPU             @                     PE           PPU                      PE           U                       UPA                                  UTU                                  UTQEE                                 @UUTUUU                             U TUUUUUU                            UUUUUUUUUU                          @UUUUUUUUUUUUU                              TUUUUUUUUU                       @U   PUUUUUUUUU                         TU  TUUUUUUUU                                TUUU                               U  @EUUU                            U @U DUU@UU                           P  TT  T                                                                      T   P                               T @ U                                    UU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                P                                      P                                      @                                    @@                                    @P                                    @Z�                                TU P���Z                                UU���ZU                              @UU���jUU                              @UU���VUUU                              PUU���UUUU                            PUUUU��UUUU                          TUUUUUU�jUUUUU             U         UUUUUUUU�jUUUUU            @        TUUUUUUUU�jUUUUU�*           P        UUUUUUUUUUU�UUUUUU�          T T      TUUU�VUUUUUU�VUUUUU�
          de  
  TUUU��UUUUUUU�jUUUUU��j         �Ui���ZUUU�Z�ZUUUUUU����UUUUU��        �������ZUU���UUUUUUU�����VUUU���  TU  jUUUUUUU�Z����UUUUUUU������jUUU��VUUUUUU3UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�W�_UUUUUUU5���UUUUUU�   WUUUUUU0 0\UUUUUU��pUUUUUU5� sUUUUUU�<�pUUUUUUU �UUUUUU�  0�UUUUUU��� WUUUUUU�  WUUUUU�  \UUUU���  \UUUU�     \UUUU5  �? \UUUU5  �� WUUUU� � �UUUUU� �  pUUUUUU_ �WUUUUU��? �UUUUUU�����WUUUU������WUUUU�����_UUUU�0��0�_UUUU�0<���UUUU� � ?|UUUU�   ��UUUU5 �0 �UUUU� �UU��?0�  pU�  0?�?  _UU����� �WUUUU?�� �UUUUU5�< � WU���� ����5    ��   ����?3����UUU5����\UU��?��pU�  ������UU��? �5  �UUU5  �  �UUU  �  pUUU  � �_UUU�����UU3UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUU�W_UUUUUUU5��UUUUUUU� 0 _UUUUUUU� �UUUUUUU� WUUUUUU500\UUUUUU�0�pUUUUUUU� sUUUUUU�  pUUUUUU���UUUUUUU�0�UUUUU��� WUUUU5��  WUUUU5     WUUUU     WUUUU     WUUUU   � WUUUU5  ��UUUUU� �� pUUUUUU��? \UUUUUUU���UUUUUUU5 ��_UUUUU��?���UUUUU�?�?��UUUUU��0��WUUUU=��30�WUUUU53��_UUUU5 < _UUUU5   �pUUUU ? UUUU��� pU����?  \U5  �� �WU������ �UUUUU��?�UUUUU?�<�UU���� ���    33  ����������UUU���<WU������ \U5  0��5� pU��� p  pUUU  p  pUUU  p  \UUU  p �WUUU���_��_UU3UUUUU�UUUUUUUUU�_UUUUUUUUpUUUUUUUU0�WUUUUUUU5� \UUUUUUU� �UUUUUUU�  WUUUUUU�0\UUUU��U=�pUUUU5 W0 sUUUU � 0 pUUUU � � \UUUU \� sUUUU �3 �pUUUU  �  pUUUU   �UUUU�  0  �UUUUU    �UUUUU�    pUUUUUU?   pUUUUUU�  \UUUUUUU=  WUUUUUUU��UUUUUUUU� pUUUUUUU�? \UUUUUUU5 ��_UUUUU��?��UUUUU�?�?��UUUUU��0��WUUUU=��30�WUUUU53��_UUUU5 < _UUUU5   �pUUUU ? UUUU��� pU����?  \U5  �� �WU������ �UUUUU��?�UUUUU?�<�UU���� ���    33  ����������UUU���<WU������ \U5  0��5� pU��� p  pUUU  p  pUUU  p  \UUU  p �WUUU���_��_UU3UU�W_UUUUUUUU�|sUUUUUUUU���UUUUUUUUUWUUUUUUUU|UUUUUUUU0�WUUUUU�W50 \UUUUU\5� pUUUU� p��UUUU5 p5 WUUU5 �5 00WUUU5 �5 0 WUUU5  ?��UUUU�  �  sUUUUU � �UUUUU 0 �UUUUU� �   WUUUUU    WUUUUU=    WUUUUU�  �UUUUUUU  pUUUUUUU5  \UUUUUUU� \UUUUUU�?  WUUUUUU5  �UUUUUUU� �UUUUUU�����UUUUU������WUUUU��00�_UUUU�0����_UUUU�0<� �UUUU� � <|UUUU�   ��UUUU5 � �UUUU�? �UUU�?0�� �UUU= ?��� pUUU�����? pUUU3  ��? \UUU����  \UUU0����?WUUU���UUUU���� ���    33  ����������U ���UUU����5  �UUU5  �  �UUU����  pUUU  � �_UUU�����UUUU��VUUUUUUUU��jUUUUUUUU���VUUUUUUU
���VUUUUUU诪��UUUUU謪���ZUUU��������j
��������UU����jUUUUUU���ZUUUUUUU���UUUUUUUUU�VUUUUUUUU��VUUUUUUUUUUU��jUUUUUUUUUUU���VUUUUUUUUUU
���VUUUUUUUUU诪��UUUUUUUU謪���������������������V
�����������VU����ZUUUUUUUUU���ZUUUUUUUUUU���UUUUUUUUUUU��VUUUU���VUUU����ZUU�����������VU����ZUU����UUU���VUUU��jUUUU��ZUUUU��UUUUU6UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��WUUUUUUUUU��\UUUUUUUUUU�UUUUUUUUUU0 WUUUUUUUUU5� |UUUUUUUUU5� �UUUUUUUUU�� WUUUUUUUUU0\UUUUUUUU� �\UUUUUUUU5  \UUUUUUU5 0 WUUUUUU��5���\UUUUUU5 �0 <\UUUUUU5 <�  \UUUUUU5     \UUUUUU5     \UUUUUU�    WUUUUUUU=    WUUUUUUU��  �UUUUUUUUU�? pUUUUUUUUU��\UUUUUUUUU5  �UUUUU���W���_UUUU5  �����UUUU��������UUUUUUU������WUUUUUU?0��\UUU���� ����UU   ���   �UU���<3����UUUUU��  pUUU����   pUUU5  0��� pUUU����0��3 \UUUUUU�����WUUUUUU�����UUUUUUU�?��UUUUUUUU����UUUUUUUUU?���WUUUUUUU�����_UUUUUUU�?3��pUUUUUUU5���?�UUUUUUU5<�=� WUUUUUU���? \UUUUU�  �  \UUUUU  0   \UUUUU  0   WUUUUU  �  �UUUUUU�����WUU.UUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_�UUUUUUUUU����WUUUUUUUU0  \UUUUUUUU� �pUUUUUUUU5  �UUUUUUUU� 3 �UUUUUUUUU���UUUUUUUUU 00WUUUUUUUU �WUUUUUUUU WUUUUUUUU�   \UUUUUUU��  \UUUUUUU?   \UUUUUUU�   \UUUUUU�   � \UUUUUU�  �WUUUUUUU ?  WUUUUUUU� �UUUUUUUU| p_UUUUUUU�W� ��UUUUUUUU����WUUUUUUU���?�_UUUUUUU=��UUUUUUU�<<��UUUUUUU3���UUUUUUU�   WUUUUU�0 �� �WUUUUU5< <  WUUU��?��� �UUUU ��3�  |UUUU����? �_UUUUUU5����WUUUUUU��� �\UUUU��?�? ����WU�    033   \UU��?�������WUUUU�0??��sUUUU��?���0�UUUU  ?_� WUUU���  �   WUUUU5   7   WUUUU5   7  �UUUUU5   7  UUUUU�������UUU.UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUUUUUUU �WUUUUUUU��   \UUUUUUU�� �pUUUUUUU�  �UUUUUUUU= 3 �UUUUUUUU����UUUUUUUUU 00WUUUUUUUU �WUUUUUUUU  WUUUUUUUU3  \UUUUUUU�5  \UUUUUUU3  \UUUUUUU    \UUUUUU�   � \UUUUUU�  �WUUUUUUU ?  WUUUUUUU� �UUUUUUUU| p�UUUUUUU��? ��WUUUUUUU���?�_UUUUUUU=��UUUUUUU�<<��UUUUUUU3���WUUUUU� �� �WUUUUU50 <  WUUU������ �UUUU  �3�  |UUUU�����? �_UUUUUU� ��UUUUUU� 0 0�WUUUU�� 0 ����_U� 0  �   pUU�?  �����_UUU5  0�WUUUUU5  �WUUUU�?   � WUUUU0    WUUUU�� 0  �UUUUUUU�����_UUU ��? ��?�����?��3?����� ��? ��? <3 <3 ��                                                                                                                                                                                                                                                                                                 �(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �*�*                                   �
�   ��         T                     P!@�����         U                     T U� � V�     @ U                     T�U�@j     @ U                    T�UVHP`     @@U                    T�ZVhh     P@                    ThV`�J     P@                   T`�Vah�     TQ@    @U            Th�V�Ua�     TUPUT    @T            TUh�V�U`�      TUPE   @E            TUh�V�U`�      UUQUUU   @U           TUh�V�Ua�     PUUQUUUUU  @U@ @U       TUh�VUUa�    @UUUU TU  PUPU PU       T��UUU`�      TUUT     U@APQ       T��UUh�    TU@UU@UA  PUPT PQ       T��UUZ�     P         PQTQTU      TU��UUZ�      UP      PUUUUTUU      TU��UUZ�               PUUUUEUT     TU��UUZ                 PUUUTUUUU     TU��ZUUZ!                TUUUUUUUUQ    TU�XUUZ                 TUUUUUUUUU    TU�JU(                UUUUUUUUUUU   TU�HU(                 @UUUQUUUUU   TU�U(Q
               @UUUQU  PUUU TU�UU                    PEUU     TU�U�TU�                 PUUUTA UUUU TU�U�TU�                    UTP       TUU
VU�                      T      TUUBUU�                     UU  T     T�UJTU�                      @U      T�UFUE)                        T      T�VVUE	                               TEYVU
                                TYVU�                                TZRU                                TV�BU                                TV�PU                                T�V�TU�                                T�V�TU�             
                   T�U�UU!           ���         ����
     T�U�UQ            hUU�*       `UU�
    TEU�UQ��*       �VUTT�       �UUTU�
   T�U�U(  �*   ���jUUUU�*      ��UUUU��
 T�UUU�*   �����jUYUAFUV�*     jU�UV  ��T�UVU�� �UU�UU@�P������VTU�  TaUUU�"@ DYVA   @    PA@   T`�VU�
   PD  @@       @�D    Td�UUa�    $         @   @ ` @ X�UUa�                 � �   �@TZ�UUa�                  @         @   TV�UUa�                                TV�UUU�                                 TU�UUU�                                 TUaUUU�                                 TUaUUU�                               ��TU`UUU�                  
  ��*      ��UTUhUUU�            �  �������j    �VeETUXUYUU��         ��� �VU�UU�U���
�VQUZTUTUXUUfU����
    �Z���VUETUUUUVUe�ZUUUUTUYUTUUVUUUfY��@��ZUUUfUEUUUUTUEUVUUYUUTUaUTU�UdYUU�j�U�QUUUUYTVYU�UTUHQUUUURTUePUUUUU%UUYUUUUUUUUUUUUUPRUUUUUTUUYU��@�UU�VUUUjUUU TUPPU@PUEUUTUUUU�  @ TeUeT%@ @@% T	 DA  PeA�TUUTU�    @  @UUE@ @(    �   U  TUVXU�        @         @ D  TUUUXU�
         P              TUVUhU�)                                TVh�!                               T�ZU`U�%              ��               T�TUaU`!             �jU�*       ���    T�UUeUa!            ��UYU��    �ZU��  T�UUha!         ��FTVUUQQ�� ��VUUUQ�
 T�UU�Ua��
     ���jEVUUUTUEUZ��UUUUU��T�UUhU`��* �����UUUUTUVQUUTEEQeUUUQUVQeQT�UEXUae���j�jUUUUUeUUUUTUUUUUUTYUUT�UUXUaeUUV�UUUUUTU`PU@PUEUUUTAT�UXUa� TT�UT@  @@ T DA@ PUA@DDQT�UUXUa� @UUF@ @        U  P T�UXU��    @          @D      TUUZU��@   @                 TUUZUa�                               TUUZUa�                               TUUjUa�                                TUUUZUa�                                TUUUjUa�                                TUUZXU��                                TUUYXU��                                TUUYXU��                                TUUYXU��                                TUUYXU��                                TUUYXU��                                TUUYXU��                                TUUYXU��                                �(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   T                                     @U                                    PU                                    TU                                   UU            @                      TU@          @U                    @U UU@          @e                  @UUP          @e                 @AUUP          @e  T     T         PAUUP          @e T     E        PUAUUTU          @E UU             TUAUUTU         @U @UT    @        TUAUUTQ  P     @U @UT    @U        TUQUUTU  PU     P PU �   @U        TUQUUTU  TU     PjTU T  PU      @UUUQUUUU @UU    Pe!TU P	  UU     UUUUUUUUUUUU PUU    Te%TU P	 TUUU   @UUUUUUUUUUUTUTUU    TUUUUUZ  @UU    @UUUUEUUUUUUUUUUU    UUUUUU�PAUTU      UUUUUUUUUUUUUUUUU@UUUUUUA              @UUUUQUUUUUUE  PA TUP   PU       PDUUUUU UUUU   TTPA@           @UU @UU   UUU    TQA                   T   P  U @EU PPUQ TU                        U  TU     E                            PU      D                                      P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            
                         ����         ���                      �VUE�       ��ZU�          ��         �VUQU%       �UQQU)        ��*"*��   �*VUUUe�      �jUUUU����  ��   �Z��*�� PYEeY�
    ��UYTUV������     �UU	  � dUUAU������EU !@PEEUeYU%    T     @AP    @ @�@@TY@ �@ @      !@          AU @  @ @     �  � @       �  �H          @                                      �j�                                   �ZUe�
     ��j   
                  �  ��U�U�
   ��ee����
  (              j�jUTVZUT) ���VeUU�UU�
���         ���U���UUUUUUU��UUYUUUUUU���Y�    ���jZ�UUU�EUUEUUUVUUYUUQUUUU�YUUU����U�YUUUYQTUTUUXUUUURUQeUUVYQVUUUUdUe�jUUUF�QEUU	UUUeQUUUUUXPUUUEUUUUUUEEUUUUVU�UEUUAPVDeQE@E QUUU YUPPU@TUU�ZUUUiUU%@ ��U%�U  � V� �U�U�EV @   P@��@ P  @ @    �  UU              @@     H       D@       @                   R                   �         �                                          @                                                                                                                                                                                                             ��              �*                    �jU�*       ��  ��V��                  ��UYU��    �ZU �jYUU���*            ��FTVUUQQ�� ��VUU�jUeQEUYU�����
     ���jEVUUUTUEUZ��UUUUEUTVUTV���* �����UUUUTUVQUUTEEQeUUUQQUUETeUUU�V���j�jUUUUUeUUUUTUUUUUUDP �A@EYUUUV�UUUUUTU`PU@PUEUU  @ @  @ TT�UT@  @@ T DA@ PUA@ @      @ @UUF@ @        U               @          @D               @   @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      UUU��UUU�UU��WUU�_U3?\UUw��30pUUw��0�UUuw7 �_UUw �\UUu   \UUU=   \UUU5  �WUUU�  �UUUU� <WUUUU �]UUU��0sUUU�?0pUU��<���UU�����UU�����_UU5�?�_UU5��<�UUU=���pUUU=���pUUU� ��pUUU�0��|UUU����_UUU� \UUUU _UUUU WUUUU���WUUUU� WUUUU5 \UUUU���_U UUUUUUUUUUU��UUU�UU��WUU�_U3?\UUw��30pUUw��0�UUuw7 ��_UUw �\UUu   \UUU=   \UUU5  �WUUU�  �UUUU� <WUUUU �]UUU��0sUUU�?0pUU��<���UU�����UU�����_UU5�?�_UU5��<�UUU=���pUUU=���pUUU� ��pUUU�0��|UUU����_UUU� \UUUU _UUUU���WUUUU� WUUUU� WUUUU���_U2UUUUUUUUUUUU���_UUUUUUUUUUUUUUUU�   �UUUUUUUUUUUUUUUUU� WUUUUUUUUUUU���U �\UUUUUUUUUU�����W5 �?pUUUUUUUUUU������  ��UUUUUUUUUU�����U �WUUUUUUUU��0 �� ��WUUUUUUUU���� �U �_UUUUUUUU����? �_���UUUUUUUU��������UU��UUUUUUUU������? �WU��UUUUUU�U�?�_����U5�WUUUUU�_�?�W���?�U5�_UUUU����? W���� �W��_UUUU����� W5 ���_��UUUU����� W �?����UUUU������  ����?�UU�W�����<   ��?�0�UU������   ��?��UU���U���?   �����]UU��U����    ������WUU�_U���?<   ��?�_UUU�UU��?�  �?|��?��_���UU���  �?|��?���s5p�WU��� �?p]�����5\WUU�� �?���_U���5WWUU�<? <���pU�����UUU��< �����U��UUUUUU��� ���_�U�WUUUUUU��� ���\�U�\UUUUUUu0��?�=puUs5\UUUUUUu50��p�_UU��_UUUUUUu5���\]UUUWUUUUUUUu5��<?\]UUU�UUUUUUUU��� � \]UUUUUUUUUUUU�� � � W]UUUUUUUUUUUU��� � WWUUUUUUUUUUUUU��� WWUUUUUUUUUUUUU� 3 � �UUUUUUUUUUUUUU]�0 wUUUUUUUUUUUUUU]��3�uUUUUUUUUUUUUUU�5���]UUUUUUUUUUUUUUU��<p]UUUUUUUUUUUUUUU�<�_WUUUUUUUUUUUUUUUU� ��UUUUUUUUUUUUUUUUU�pUUUUUUUUUUUUUUUUUU5 \UUUUUUUUUUUUUUUUUU� WUUUUUUUUUUUUUUUUUUU�UUUUUUUUUU:UUUUUUUUUU����WUUUUUUUUUUUUUUUU5   |UUUUUUUUUUUUUUUU� ��UUUUUUUUUUUU���_U � WUUUUUUUUUU�����U �\UUUUUUUUUU��?��_5  ?pUUUUUUUUU���<�� ��UUUUUUUUU��� ��_= ��UUUUUUUUU�� � 0 ���WUUUUUUUU�������W�?�_UUUUUUUU�?������_U��_UUUUUUU��?���� �UU�UUUUUU���W�����WU��UUUUUU����U����_U��W�UUUUU��WU��� U����?WUUU��?�_U����W����?\UU���� |UU��? ?����\UU���� �UU� ���W�W_UU������WU������_U�_�����|���� ����pU5�����?< ���������U������  ��?���5W�U��U���   ������_5\�U��U��?   ������_�pUUU��U��   �_���UU_UUU��W��    _���WUUUUU���_U��   <\�?�\UUUUU�p5\U��  �p���pUUUUU�\\U5�  ��U��pUUUUUUWWU� ���u�_UUUUUUU�Uu�3 0� w�UUUUUUUUUUu�� �< ���UUUUUUUUUUu�� 0? �_WUUUUUUUUUu �� �WUUUUUUUUUu �� �s5WUUUUUUUUUu5���0 ���UUUUUUUUUUu�� 0�uUUUUUUUUUUUu� puUUUUUUUUUUUUu� ���puUUUUUUUUUUUU�UpuUUUUUUUUUUUU�U��\uUUUUUUUUUUUU�U\uUUUUUUUUUUUU�U\]UUUUUUUUUUUUUW� 0\]UUUUUUUUUUUUUW0� \]UUUUUUUUUUUUUW0�� W]UUUUUUUUUUUUU]5��? WWUUUUUUUUUUUUU]���<�UWUUUUUUUUUUUUUuU3��pUWUUUUUUUUUUUUU�U� �_�UUUUUUUUUUUUUUU�����uUUUUUUUUUUUUUUU}5��U_UUUUUUUUUUUUUUUU��pUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUU� pUUUUUUUUUUUUUUUUUUU\UUUUUUUUUUUUUUUUUUUWUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUDUUUUUUUUUU����WUUUUUUUUUUUUUUUU5   |UUUUUUUUUUUUUUUU� ��UUUUUUUUUUUU���_U � WUUUUUUUUUU�����U �\UUUUUUUUUU��?��_5  ?pUUUUUUUUU���<�� ��UUUUUUUUU��� ��_= ��UUUUUUUUU�� � 0 ���WUUUUUUUU�������W�?�_UUUUUUUU�?������_U��_UUUUUUU��?���� �UU�UUUUUU���������WU��UUUUUU���W����_U��W�UUUU���UU��� U����?WUUU��sUU����W����?\UUU��?�UUU��? ?����\UUU����WUU�����W�W_UUU����_UUU������_UUUU����UUU��� ����pUUUU�����UUU�������UUUUU���UUUU����5W�UUUUU��?�WUUU����_5\�UUUUU����_UUUU���W�pUUUUU����UUUU���UU_UUUUU�����UU�_U�UUUUUUUU����?�WU�UUUUUUUUUUU����?�_��UUUUUUUUUUU���������UUUUUUUUUUU�����  ���WUUUUUUUUUU����  ���WUUUUUUUUUU����  ���_UUUUUUUUU��_�?   ���_UUUUUUUUU��W�    |��_UUUUU�_��UU�  �p���sUUUUU5��UU�  ��U���UUUUU��_U��  ��W���UUUUU��WU5�?  ����UUUUU���U�5�� �����UUUUUUU��U�5���� ��WUUUUUU��W�5 ��� �\UUUUU���_�5 ��? ��5\UUUUU�p5\�5 ��? ���\UUUUU�\\�� �?�� �WWUUUUUUWW�U<<� ��UUUUUUUUU�U�U<0<��UUUUUUUUUUUU�U���3��UUUUUUUUUUUUUW00��UUUUUUUUUUUUUW��p�UUUUUUUUUUUUUW00p�UUUUUUUUUUUUUW00puUUUUUUUUUUUUU]0�?puUUUUUUUUUUUUU]5���puUUUUUUUUUUUUU]5 �� \uUUUUUUUUUUUUUu���3\]UUUUUUUUUUUUUuU��W]UUUUUUUUUUUUU�U��?�U]UUUUUUUUUUUUUUW�  UWUUUUUUUUUUUUUU]�����UUUUUUUUUUUUUUU����W}UUUUUUUUUUUUUUUU��?WUUUUUUUUUUUUUUUUU��WUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUUU5\UUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUU��  ��  �� �0 �p�������������������� ��� ��� �� �� �� ��  �� �� �� �� �� ����_x�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      @                                      PU                                      U                                      PQ                                      PU                                      PU                                      TU                                      DU                                      TU                                      T                                      TU                                      TU                                      TU                                      UU                                      UU                                     @UU                                       P                                     PUA                                                                            T             @                                    P @                                    P @U                                    PPU                                    PE                                    PE                                   UPA                                  UTU                                  UTQEE                                 @UUTUUU                             U TUUUUUU                 �
@U      UUUUUUUUUU                 dT    @UUUUUUUUUUUUU                �AQUUQ        TUUUUUUUUU               `TUUUE  @U   PUUUUUUUUU              dUUUZU    TU  TUUUUUUUU              YU�UU�U           TUUU                V�UUUU        U  @EUUU               �U�AUEUU     U @U DUU@UU             �U�T�PU�      P  TT  T              jT)UePd                             UU�YU           T   P              �UUUZVU        T @ U               �UjTU�U            UU                 �T�QVUUE                               �T�QYUUU                               �jP�F%UQU                               �j@UV� h                              ��UU��Z�           P                   ��PUU�U�           @U                   ��BUUUU�             UU         P      ��
UUUUU                         P     ��PUUU                         T      �j@�UUQ                        T      ����V`                        T      ����� Z                        U      ������V                      @Q U      ������Z                      @A U       ������                      PE@      ������                      PUAUP       P���                      PUAUT       P�*                       TUEUUU      P�                       @UUEUUUUU     P�                       UUUUU PU  @ |�                       PUUP    @ ���                     PUUU U    D��j�                     @@     PU ��o��>                                  ��~��                                 �����*                  P       @UU   *����                 @      P      ������                 P     T       ����>�                       @        ��
�  j                               ����
   Z           PUUU               � �j��
T                                 �V��*W                                �V����W                                 �U����U                                 ��ZUjU                              @  j�VU�U                               @�Z��UU�V                                �Z�jUU�V                               �V�ZUUUV                               �V�VUUUY                               �U�UUUUU                                �U�UUUUU                            � �jUjUUUUU                               �jUjUUUUU                               �ZUjUUUUU                               �VUjUUUUU                            @�UU�UUUUU                              jUU�UUUUU                              �VUU�UUUUU                              �UUU�UUUUU   UUUUUUU                    jUUU�VUUUU                             �VUUUUVUUU�                             �UUUUUZUUU�                            �ZUUUUUYUUUj                           @�UUUUUUiUUUV                          PUUUUUUUUeUUUU            TUUUU       UUUUUUUUUUUUUUU                       PUUUUUUUUUUUUUUUU                        TUUUUUUUUUUUUUUU                         UUUUUUUUUUUUUUU                          TUUUUUUUUUUUUU                           UUUU�ZUUUUUUU                            @UUU�UUUUUUU                             @UU�VUUUUUU                              TU�jUUUUUU                    TUU       @UU�ZUUUUU                       T       UU��VUUUU                               PU���UUUU                        @      UU�jUUUU                         @U     PUUUUUUU                           U     PUUUU        �                         TUU         �
                          TU         @ji                                    T�ZU                                  @U�VUUUU                               PU�VUUUUU                               UU�VUUUUU                             PUU�UUUUUU)                             TUUiUUUUUU��                          PUUU�UUUUUUU��                        PUUUU�VUUUUUU���                       �VUUUUUUU��UU�����                      �ZUUUUUUUU�jUU������                   ��jUUUUUUUU��UU������
                 �UUUUUUUUUUUU��UU����Z�Z��UUUUUUUUUU�ZU���(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 @                                  P P                                  T T                                  PP T                                   T                                  UU DU                                  UUU UU                                 UUUEQU                                 UUUUUU                                UUUUUUUT                                UUUUUUUU                               UUUUUUUUU                               UUUTUUUUU                              UUTU  TUUU                                TQUU                                 UUUP@UUUU                              @U                                     U@                                  @U  U                                   PUA                                      U                                      @                                                                                                                                                                                                                               @                                      @                                      P         �                          P         A                          P                                  T T         h                         ET         UT                         TQ         UUT                       @TP        VU�                      @UUU@       XUB
                      @UUTQ       X�	                      PUUUUU       V�U(                      UUUUUUU     XU(                     TUUUU@UU      EV)                      @UUU@        �V*                    @UTU TT      �V�*                            @U   ���
                                    jU�
                                    VU�                           UU     UU�                         @         U�                       PPU          U�                         U           ��*                                     �                                     *                                     �                                     �             @                        *           P @                        
           P @U                                    PPU                                    PE                                    PE                                   UPA                                  UTU                                 UTQEE                                 @UUTUUU                     @      U TUUUUUU                           UUUUUUUUUU                         @UUUUUUUUUUUUU @U                         TUUUUUUUUU                      @U   PUUUUUUUUU                    j   TU  TUUUUUUUU                    j           TUUU                      i�       U  @EUUU   UUUU              �    U @U DUU@UU                    �    P  TT  T                     U                                 U         T   P                      U      T @ U                       U          UU                         U                                      UU@                       TUUUU       UU   �                                 UU P                                 UU
  P      P                           AU	   (     @U                          U)�         UU                       )T*                                    ��*                                     ���                                     U��@ @                                 U��*                                    U���                                    UկV
                                  ZU�U%                                   jU�U%                                   �UiU� @                                 �VeU�                                  �ZeUU
                                  �j�UUU                                  Uj�VUe                                 U�UVU�V                   TU  TUUUUU  U�VUU�Z                TU              U�VUUUUUU                              U�ZUUUUUQU                             UUZUUUUU PU                            UUiUUUUU @U                          UU�UUUUUUUU @U TUU                     UU�jUUUUUUUUU@UU                       UUU�VUUUUUUUUUU                        UUUUUUUUUU���                          UUUUUUUUU�
                               PUUUU�*     @UUU                        TUU��                   @UU              ���
 PUU           U ��ZU                               @U�A��UUU                               PU���ZUUU                   @UU      PUU��VUUU          @ @U              TUU��UUUUU          PU               TUUU��UUUUU                          UUUUUU��VUUUUU                       @UUUUUUU��ZUUUUU                       UUUUUUUUU�ZUUUUU�
                    @UUUUUUUUUU�jUUUUU��                    UUUU�UUUUUUU�UUUUUU�              �  UUUU�jUUUUUUU�ZUUUUU��  *         ���VUUU���VUUUUUU���jUUUUU��  �     ��������VUU��jUUUUUUU�����UUUU��* UUU���VUUUUUUU�V���jUUUUUUU������ZUU���U.
�_�UUUUUUU���_UUUUUU �_UUWUU�  pUU_UU5 ? �UWs]U� � ��\ssUU� ��\ssUU= 00�\ssUU ��\ssUU� �\ssUu�  �\ssU��  �\ssU�  �\ssU    �\ssU    �\ss�  �� �p�pU ? �U�0\U�  �_ \U5�? ��� WU�����_WU�?���5W��������5W�?<30�7W�����=_5< �  �p       <s       �p0�  �0s�  �<�p �3 <��?s �� ��5_��?���_5W50�� ��_5W�� � W5WU�� ��W5WU�?���W5WU��<?W5WU��3���U5WU� <�?W5WU��< \5WU p� p5W�  p} �7W  pU  W  \U  0W  \U5  W���WU����U.
�_�UUUUUUU���_UUUUUU �_UUWUU�  pUU_UU5 ? �UWs]U� � ��\ssUU� ��\ssUU= 00�\ssUU��\ssUU �\ssUu�  �\ssU��   �\ssU  �\ssU    �\ssU    �\ss�  � �p�pU ?��U�0\U�  �_ \U5�? ��� WU�����_WU�?���5W��������5W�?<30�7W�����=_5< �  �p       <s       �p0�  �0s�  �<�p �3 <��?s �� ��5_��?���_5W50�� ��_5W�� � W5WU�� ��W5WU�?���W5WU��<?W5WU��3���U5WU� <�?W5WU��< \5WU p� p5W�  p} �7W  pU  W  \U  0W  \U5  W���WU����U.
UUUUU��WUUUUU���WUUUU� 0�UWUUU  pU_UUU� � \Ws]UU3 � �\ssUU� ��\ssU� |�\ssU�0 ��\ssU�� ���\ssU�  0s�\ssU5  0_3\ssU5  ���\ssU5    �\ssU5    �\ssU� � �p�pUU� p�0\UU  p \U�� �?�� WU������_WU�?? ��5W��������5W�?<30�7W�����=_5< �  �p       <s       �p0�  �0s�  �<�p �3 <��?s �� ��5_��?���_5W50�� ��W5W�� ��U5WU�� ��U5WU�?���W5WU��<?W5WU��3���U5WU� <�?W5WU��< \5WU p� p5W�  p} �7W  pU  W  \U  0W  \U5  W���WU����U.
UUUUU��WUUUUU���WUUUU� 0�UWUUU  pU_UUU� � \Ws]UU3 � �\ssUU� ��\ssU� |�\ssU�00��\ssU�� ���\ssU�  �s�\ssU5   _3\ssU5  ���\ssU5    0\ssU5    �\ssU� �  s�pUU� ��0\UU  p \U�� �?�� WU������_WU�?? ��5W��������5W�?<30�7W�����=_5< �  �p       <s       �p0�  �0s�  �<�p �3 <��?s �� ��5_��?���_5W50�� ��_5W�� � W5WU�� ��W5WU�?���W5WU��<?W5WU��3���U5WU� <�?W5WU��< \5WU p� p5W�  p} �7W  pU  W  \U  0W  \U5  W���WU����U.
U�WUUU�UUUU=\U]U_UUU\uwWp_UU����ps]U �� \ssU5 ��  WssU�< �\ssUU� ��\ssUU 3 �\ssUU�� �\ssUU<�\ssUU�< ��\ssUU�����\ssUU? ?�\ssUU   �p�pUU�� \�pUU5< W \UU5 0W5 WU��  ���WU������_5WU�? 0�5W��������5W�?<?�7W��0 ��=_=<���  �p   � <s�00    �p00  �0s 00  <�p �0 ���?s �� �5_ �?���W5W5��� ��U5W��  ��U5WU��� ��U5WU�����W5WU���<?W5WU��<���U5WU� ?�?W5WU��< \5WU  �  p5W�  �} �7W  pU  W  \U  0W  \U5  W���WU����W.
U�WUUU�U_UU=\U]UWs]U\uwW�\ssU�����\ssU ���\ssU �� �\ssU� ���\ssUU?3�\ssUU���\ssUU  �\ssUU??�pssUU�����pssUU? ?p��pUU�� p\UU< \ \UU 0\5 WUU�  �W�WUU����UU=WU�� ��U5WU�� ��_5WU������5_����3���p�?<����p��0 ��<s< ��  �p     � �p�?     0s��  �0\?  <0W�0 ���?W�� �5W5�?���W5W��� ��U5WU< ��U5WU��� ��U5WU�����W5WU���<?W5WU�?<���U5WU�?�?W5WU��< \5WU  �  p5W�  �} �7W  pU  <W  \U  �W  \U5  \U���WU���WU.UUU�W�_UUUUUUUUU5���UUUUUUUU�   WUUUUUUUU0 0\UUUUUUUU��pUUUUUUUU5� sUUUUUUUU�<�pUUUUUUUUU �UUUUUUUU�  0�UUUUUUUU�� ��UUUUUUUUU3  WUUUUUUU=  WUUUUUU���   WUUUUUU�     WUUUUUU5     WUUUUUU5  <�UUUUUUU� ���UUUUUUU� <  pUUUUUUUU� �_UUUUUUU��� ��UUUUUUUU�����WUUUU����?���_UUUU5  ���0�UUUU���0<<��UUUUUUU� �?�pUUUUUUU� _UUUU��������UU    33  �UU���������UUUUU�?  WUUU���� �� �UUUU5  ����UUUU���??���UUUUUUU�����_UUUUUUUU3  WUUUUUUUU����_UUUUUUUU�3��UUUUUUUU�����UUUUUUU�?�<WUUUUUU���� \UUUUUU= ?7� pUUUUU�    pUUUUU5  �   pUUUUU5  �   \UUUUU5    �WUUUUU������_UUU.UUU�_�UUUUUUUUU����WUUUUUUUU0  \UUUUUUUU� �pUUUUUUUU5  �UUUUUUUU� 3 �UUUUUUUUU���UUUUUUUUU 00WUUUUUUUU �WUUUUUUUU WUUUUUUUU�   \UUUUUUU��  \UUUUUUU?   \UUUUUUU�   \UUUUUU�   � \UUUUUU�  �? WUUUUUUU � WUUUUUUU�� �UUUUUUUU| p_UUUUUUU�W� ��UUUUUUUU����WUUUUUUU���?�_UUUUUUU=��UUUUUUU�<<��UUUUUUU3���UUUUUUU�   WUUU���     WUUU5      WUUU���0   WUUUUUU��?�UUUUUUU� pUUUU���� ���UU    33  �UU���������UUUUU�  �UUUUU�������WUUUU5  p����UUUU����3��pUUUUUUU=���?�UUUUUUU��?� WUUUUU� �|�? \UUUUU  \  \UUUU�   �   \UUUU�   �   WUUUU�   �  �UUUUUU���W��WUU.UUUUU���WUUUUUUUUU� �UUUUUUUU5  �UUUUUUUU�  WUUUUUUUU� 0\UUUUUUUU0�\UUUUUUUU5� \UUUUUUUU�  sUUUUUUUU5  �pUUUUUUUU5< 0pUUUUUUUU��  �UUUUUUU�_�  �UUUUUUU5�<  �UUUUUUU5    �UUUUUUU    �UUUUUUU  �pUUUUUUU5 �? pUUUUUUU5 � \UUUUUUU��?  �WUUUUUUU�?��UUUUUUUU�����UU��UU�����WU �UU5��0�_U��WU53��sUUU5\U��?< ?\UUU�p� �  �WU��?�? ���� \�    033   pU��?������� pUUU�pU5 � pU��?\U��? \U  WU<0���WU���U�<����UUUUUU5�<�?�UUUUUUU5 ���WUUUUUU� ?���_UUUUUUU�����UUUUUUU�?3���UUUUUUU5���<WUUUUUU5<�� \UUUUUU��5� pUUUUU�  p  pUUUUU  p  pUUUUU  p  \UUUUU  p �WUUUUU���_��_UU���U���U����U����U �����������w����w����w����uU���uU��_uU p]U��]U���]���]����W����_� ��p����s�����WWUW�UU�UUU                                                                                                                                                                      �(                                                                                                                                                                                                                                                                                                                                                                                                                                           ?                                      ��                                       ?                                       7                                      ��                                      ��3                                     _?<                                    ����                                     ��                                     ��?                                    �ww�                                    ����3                                    0?                                  @p�0C                                  Pq�S                                  p�                                   p�                                   ����            ���                   |www            ��U<                  0\www           p�U1                  �_���           ��W�                 7��1           �_U=                 7���1           �|U5                  7��1            �Utq5                  W}U<0            _U}p5                 �UqU�            OU}p5                 �wU|�            OU}|5                 ������0          �OU}|5                ��������          �_Uqp�                �|�����         �WU�q�               �W����u�          �WU�q5               \w��uw        ��WU�q5               T��}w��C        ��WU��u               0pU           p�UU��U                p}           p�_U��U<                p�  3         P�WU��U<                p�� 7         \�]U��U1               p���7         \�]U��U5T              |��7         |�UUU�U5U              \}}<         |uUUW�U5U              \UqU          \uUUW�U5T              ��}U|w         \uUWEUuE             ������?�        \uUU\EU�              ���uw���C       \uUU\@U�              ��uw��7�        \uUU\pU              �uw���        _}U_qU              �u]w��u        WuUWqU�              w�]�uw�        W}UWqU�             @�w�}��?@       W}UUq�              @_U    �@      �W}UWu�               WW   ��       �U}UWU�                �_ � ��        �U}U�WU�               7p���        �UU��U               �����        �U_U��U              7s|<��        �UWUu�UW              �7s\W0��       �UWUU�U             ��_�U��       �UWUU�UUW              �UW�U1�        p�WUU�UU              �UU�U�         p�WUU�UUG              pUU�U�         p�UUU�UU              |}�U�<�<       |�UUU�UU ��           ��������       \�UUU}�UU 0�         �u]w��u�      _�UUUU�UU p        �|u]w��u<p     U�UUU�WU p        � _u]w��u]�      _UuUUU�WU |        ��W]�u�]�u��     UuUUUEW \         �U�u]�u]��      WUuUUUEW \         ��uu�5�]]�      WUuUUU�U�_         ��}�}���      WUuUUU�U�]         \U     0T     @WUuUUU�W�]         \u�� 0T     WU5UTUW��]U<         \�0  ?00     QWU5UUUW�=�UU0          \����0      TWU5UUU_��pUU�          � ���3     @UWU�UU�U��pUUq         ������3      �WU�UU�U��pUUA         \7< <��0      �UU�UU�U��pUUA         _7__����      �WU�UU�U��UuA         W��U� ?�      �UU�UU�U��_UuA         Wu�wU��      �WU�UUU�U�W_UuU         WUwU�  �     ��UU�UU�U�UWUuU         WU�wU� �     p�UU�UU�U�UWUu        ����wU�?��    p�UU�UU�W�UWUq�W UUU  �u]�wU��u]    |UUUUUUU�W�TWU�LSUUUUU ��}�wU��}�    �UUUUUUU�U�TWU�UOUU    ����������    �UUUUUUU�UUTWUU|UUA  ��q��q��   �UUUUUUU�UT�uU|UU  �<�q��q<p  �UUUUUUU�UUT��UU1     ���q��qW�  �WUUUUUU�UUT��TUU1      �@u����q\�  \WUUUuUU�UUT�WTUU5      �Tu���q\�   \UUUUuUU�UUTUW\UT5      �T]��q�q�   _UWUUuUWUUTUW\UT5      ����qq=\��@   WU}UUuUWUUUUW���?     @�}������}?P  ��UUuUWUUUUW��      @�uU 0� P    �WUuUWUUU��        P�U]    0 T  �� ���U����U   @@      ����� ��    �?  �U�  ��TA@TD      �5 ���      ������    PUU UUU      �}�|Q��<          <DUQUUUTU     ���=��?    UA �?  � TUUUUUEQEA    �}?�WQ���<    UU@  ��� @UEUTUUU    �u���u<    UU      QUUUUUTUUU  pu=�UQ���   @UUT   UUQUUUUUEUU   p�����   UUUUAUE@@PUTUTUUUUUUUUA  pU]�Us� 0  DPUUUUUE@UUUUUUUUUUUU  pUU�3�   @PUUUEUUUQUUTUUUUTUUUUEE]|UU�Us�   <0DUUUUUUTUUUUUUUUUUUU]UUUU�������������QQQUUUEUUUUUUEUUUuUWWUU|p�UQ�|��UUUUUUUUQQUUUUUUUUUUuU]UU]]]�ps��7�\3uEAUUUUUUUUQUUUUUUUU]�UU]]]�ps�UQ�7�\34UUUUUUUUUUUUUUUUUuUU�UuWU������������UUUUUUUUUUUUUUU]UUUUUw�]UUUUU�W���WUUUUUUUUUUUUUUUUUUU�UUUU]UuUUUUUUu�   WWTUTUUUUUUUUUUUUUUUWUUU��]�UuUU]�   �uUUUUUUUUU�UUUUUUUUUWUUUU]WwUUU�U��    WUUUTUUUUuU]UUUUUUuUuUUUUuW�UuUuWU    \UUQUUUTuUU�UU�UUWUUU]WUUU]_}UWUU��   \VUUUUUUU�UU�U]�U]Uu}U�UU�_�����     _UTUUUQU_]UU����������w]�U��  �WU    �UUUUUU�����        �����?            \UUUQUUU��?  T        �_U          _w�UUQUU    T                         |UUUUUUU                          P    p�UUUUE                         @    pUUUUUUU             UU       TUU      |WUUUTUU           PUUUU@             _UUUUUUU                              WUUUUUUU                              WUUUUUEU                              WUuUQUUU    UU E                      �W�UUUUUETTUU                          �]UWUUUUU                              qUwUeUUUU                              qUUUUUTUU                             P}WUuUUUEU�(TETETE @P @   *@@@@@P P     �P PTETE @��������*������������������������TE @���UUUU !jUUUUUUUUUUUUUU%  �VUUU @���UU  @���*�              �����   ���ZUU    @���**              �����   �UU       @���*�              �����   U         @���**              �����              @ !�              $  �          ��������**�����������������������     ���VUUU P!�VUUU     XUUU)  �hUUU   ���  V @ D * @T     X  ) @�b  D ��
    VUTA P!�UTU     XUQ)  �hPEU�VU	    �Z D D!*F ��     �j) @�b@�UEU	    �ZD P!�FP��     �jU)  �hU� TU	     �ZD D!*F��        �j) @�bD�
T��
      XD P �F�          `)  �hD	 T��
      X@ D!*�          `) @�b@	 ��    
   XE P!�F�          `)  �hT	 %        �U D!*V�          �V) @�b�
 %    �   �E P!�F)          �)  �h� *         �U D!*V)          �V) @�b�     �   �U P!�V)�����������V)  �h�        �� D!*�
PUUUUUUU�* @���     �       P!� ���������j
 (  �(               D!* ��        `)   @�  �      �     P!� ��TUUUUUUU��    �  �     ��
    D!*  (TUUUUUUU��   @�      �����
    P � (
UUUUUUUU�   �      ���
     D!* 
BUUUUUUUUX
  @�      �  @    P!���RUUUUUUUUUh�   �      �TUU    D!*`�PUUUUUUUUU��  @�      �TUU    P!�`*TUUUUUUUUU��   �      �TUU    D!*`UUUUUUUUUU�  @�      �TT    P!�`RUUUUUUUUUUU�   �      �TE    D!*`RUUUUUUUUUUU�  @�      �T     P �`RUUUUUUUUUUU�   �      �T@    D!*`RUUUUUUUUUUU�  @�      �TUP    P!�`RUUUUUUUUUUU�   �      �TD    D!*`RUUUUUUUUUUU�  @�      �T    P!�`RUUUUUUUUUUU�   �      �T    D!*`RUUUUUUUUUUU�  @�      �T    P!�`RUUUUUUUUUUU�   �      �TE@    D!*`RUUUUUUUUUUU�  @�      �TEP    P!�`RUUUUUUUUUUU�   �      �TT    D *`RUUUUUUUUUUU�  @�      �TUT    P!�`RUUUUUUUUUUU�   �      �TUT    D!*`RUUUUUUUUUUU�  @�      �TUU    P!�`RUUUUUUUUUUU�   �      �T@    D!*`RUUUUUUUUUUU�  @�      �TEE    P!�`RUUUUUUUUUUU�   �      �TUD    D!*`RUUUUUUUUUUU�  @�      �T@    P!�`RUUUUUUUUUUU�   �      �T@A    D!*`RUUUUUUUUUUU�  @�      �T D    P!�`RUUUUUUUUUUU�   �      �T    D *`RUUUUUUUUUUU�  @�      �TUE    P!�`RUUUUUUUUUUU�   �      �TA    D!*`RUUUUUUUUUUU�  @�      �TP    P!�`UUUUUUUUUU�   �      �TUQ    D!*`*TUUUUUUUUU��  @�      �TUP    P!�`�PUUUUUUUUU��   �      �TUU    D!*��RUUUUUUUUUh�  @�      �TUU    P!� ZBUUUUUUUUX
   �      �TUU    D * h
UUUUUUUU�  @�      �T     P!� `)TUUUUUUU��    �      �T @    P!* ��TUUUUUUU��    �      �dP    D � ��        `)   @�      �TP     P!*  ���������j
    �      �d T    D!�  XUUUUUUUUU   @�      �TUT    P!*  ����������    �      �dU     D!�                @�      �d    P *                 �      �T    D!�                @�      ��UU    P!*                 �      ��UU    D!�                @�  �   �T      P!*                 �  �   �  ��
    D!�               �B�      �����
    P!*               h
�      ���ZU    D!�               J)�      TUU     ���*(              J)�              �@���             �B� �              �P����"             �j�
�               TU���
            �Z����              (UU���"            ��j��
               UU���
           �Z�Z���               HUU���"           ����j��
              HUU���
          �Z���j���              HUU���"          ���j�����          ����HUU���������* �� ���Z�����*       ���   HUU���"      �  �������������   ���  ���HUU�����������


�  PTUU�
  ��*  �����HU���������*��*�
���������V� �  �������UU��������*����� (  PTUU��� ����������(T���������*���`�������������������������TU��������*��b�����������������������������������*�(b������������"��������
              �
b������������"������
  UUUUUUTUUUQUU��b������������"���
  @EUUUEUUDUUU���������������"�� @UUUE@TUQUUUDUUUUUU��VYe�UVYe�U�   TQUUUETUUQUUUDUUUUUU�
��VZi��VZi(UUUUUETUUUUUUTUUUQUUU��f�e�Yf�e�Y�QUUUUEUUUUUUUTUUUQUUU�Z����j����j���JQUUUUUEUUUUUUUTUUUQUUU�jX�VYe�UVYe�U�JQUUQUUUEUUUUUUUTUUUQUUU�jY������������ZUUUQUUUEUUUUUUUTUUUQUUU��Y�ZYe�UVYe����UUUQUUUEUUUUUUUTUUUQUUU��Y���f�i��f����UUUQUUUEUUUUUUUTUUUQUUU��Y�������������UUUQUUUEUUUUUUUTUUUQUUU��Y�������������UUUQUUUEUUUUUUUTUUUQUUU��Y�������������UUUQUUUEUUUUUUUTUUUQUUUY�Y�������������                        h�Y�������������UUUQUUUEUUUUUUUTUUUQUUU��Y�������������QUUUE@TUQUUDUUUU��Y�������������QUUUUUETUUQUUUDUUUUUUQ�Y�������������QUUUUUETUUQUUUDUUUUUUQ�i�������������UUUQUUUEUUUUUUUTUUUQUUUQ�e�������������UUUQUUUEUUUUUUUTUUUQUUUQ���������������UUUQUUUEUUUUUUUTUUUQUUU�Z�����jUU������UUUQUUUEUUUUUUUTUUUQUUU������Z�j������UUUQUUUEUUUUUUUTUUUQUUUiZ�����������j�UUUQUUUEUUUUUUUTUUUQUUUY�j�����������j�UUUQUUUEUUUUUUUTUUUQUUU�j�����������Z�UUUQUUUEUUUUUUUTUUUQUUU�����*���Z�����UUUQUUUEUUUUUUUTUUUQUUU�����*���j�����UUUQUUUEUUUUUUUTUUUQUUU�����*���j�����UUUQUUUEUUUUUUUTUUUQUUU��Z��*���j��j��UUUQUUUEUUUUUUUTUUUQUUU��j��*���j��Z��UUUQUUUEUUUUUUUTUUUQUUUY�����*���j��j��                        h���R�*���j��b��UUUQUUUEUUUUUUUTUUUQUUU����V�*���Z�je��QUUUE@TUQUUDUUUU����VT������Ve��QUUUUUETUUQUUUDUUUUUUE���VU����jUe��QUUUUUETUUQUUUDUUUUUUE��VDU�U�VUUe�
UUUQUUUEUUUUUUUTUUUQUUU����VTUI��UU���UUUQUUUEUUUUUUUTUUUQUUU����UTU���VUU���UUUQUUUEUUUUUUUTUUUQUUU�)��UTU���VUU��
UUUQUUUEUUUUUUUTUUUQUUU���jUTU���VUUU��UUUQUUUEUUUUUUUTUUUQUUU���ZUTU���UUUU��UUUQUUUEUUUUUUUTUUUQUUUE��VUTU��jUUUU��UUUQUUUEUUUUUUUTUUUQUUUE��UUTU��jUUUU��UUUQUUUEUUUUUUUTUUUQUUUEUUUUTUU�jUUUUTUUUUQUUUEUUUUUUUTUUUQUUUEUUUUTUUUEUUUUTUUUUQUUUEUUUUUUUTUUUQUUUEUUUUTUUUEUUUUTUUUUQUUUEUUUUUUUTUUUQUUUEUUUUTUUUEUUUUTU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUU��_�UUUUUUUUUUUUUU��� UUUUUUUUUUUUU�� �WUUUUUUUUUUUU��   \UUUUUUUUUUUU}?   pUUUUUUUUUUUU�?   pUUUUUUUUUUUU�   �W��UUUU�UUU�   |�pUUUU�UUU�  � ��W�WU5UUU?0     ��?\U5UUU�0�    ��� �UUU��    �������U?�0   ������< ����  �   ���������<  ?�   ��������� �    ���������U�    0 �������U�?  �   �������U ? <   � <�����U���  ��?� ����U5|UU  �\�?  ����U�|UU  _W��� ����UUUU� �U��_U���?UUUUUU|U5�_UUU���UUUUUU�WU�UUU��_UUUUUUUUU�UUU��UUUUUUUUUU�5pUUU��UUUUUUUUUUU5\UU�UUUUUUUUUUU�W����_UUUUUUUUUUUUU5���UUUUUUUUUUUUUU5��_UUUUUUUUUUUUUU5��WUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUU��WUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUU���_UUUUUUUUUUUUUUU\UUUUUUUUUUUUUUUUWUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU}U�UUUUUUUUUUUUUU_U5\UUUUUUUUUUUUU��_=�WUUUUUUUUUUUU� ��U_UUUUUUUUUU5�����_UUUUUUUUU����   pUUUUUUUU��������\UUUUU_U?��������p��UUUUp�����������? WUUU�������������\UUU ������������pUUU�����  ��������UUU����  � ����_UU����   �  �����p����<     ��������� 0���  ������� �UU��  ����� |UUUU��  ������ �WUUUUUU�? �����? UUUUUUUU� ����?�WUUUUUUUUU�����3|UUUUUUUUUU�� ���WUUUUUUUUUUU5   ��UUUUUUUUUUUU��  �_UUUUUUUUUUUUUU? �WUUUUUUUUUUUUUU� UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUU5|UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUu�UUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU5pUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUU���WUUUUUUUUUUUUU���|UUUUUUUUUUUUU�� �WUUUUUUUUUUUU��   |UUUUUUUUUUUU��   pU��UUUU�UUUU�?   ��pUUUU�UUU�<  �5�W�WU5UUU5�3  �  ��?\U5UUU��     �� �U�_U��     ���������?0    �����< �5?��   ���������5 �  0   <���������    0   ��������U? ��  ����������U��U?   ���������U�U�   < �?�����U�U�       ����U�U�   ��?   ����UUU?��  p��� ����UUU|  _��U���?UU��W� �UU��UUU���U��pUU�WUU��WUU��_U�0pUUUUU���_UU��UU�\UUUUU�p5\UU��UU� \UUUUU�\\UU�UUU_UUUUUUWWUU�_UUU�_UUUUUUU�UU��WUUUUUUUUUUUUU�_�UUUUUUUUUUUUUU5��_UUUUUUUUUUUUUU��WUUUUUUUUUUUUUU��UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU��WUUUUUUUUUUUUUU���_UUUUUUUUUUUUUU�p5\UUUUUUUUUUUUUU�\\UUUUUUUUUUUUUUUWWUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU}UUUUUUUUUUUUUUUUU_U�UUUUUUUUUUUUU��_5\UUUUUUUUUUUUU� �7�WUUUUUUUUUUU�7�<�UU_UUUUUUU_U?�����p�WUUUUUp������� �sUUUUUU����������pUUUUUU ���������\U_UUUU�����������p��WUUU�����������? \UUU����� �������pUUU���  ��������UU��� �   ������WU�� 0   �  �����\U� 0��  ������� � ��U�  ������  ? UUUU� ������??�WUUUUU��?  �����3|UUUUUUUU  ������WUUUUUUUU� ������UUUUUUUUUU� �����_UUUUUUUUUUU ���WUUUUUUUUUUU��  ��UUUUUUUUUUUUU}  �UUUUUUUUUUUUUU� �UUUUUUUUUUUUUUU� �UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUU5�UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU�pUUUUUUUUUUUUUUUU�\UUUUUUUUUUUUUUUUUWUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU>UUUUUUUUUUUUU��UUUUUUUUUUUUUUUUU�  �_UUUUUUUUUUU��_UU � pUUUUUUUUUU����_U5 �?�UUUUUUUUUU����U�  �WUUUUUUUU���?�_U �?\UUUUUUUU������U=  �sUUUUUUUU�?<  ��W� �UUUUUUUU� �� �_U= ��UUUUUUUU������U���WUUUUUUU�������WUU��WUUUUUUU����� UU��_UUUUUU���������WUU�UUUUUU����_����_UU�UUUUUU����WU��? �UU�UUUUUU����WU����_U�UUUUUU���_UU��? ���_UUUUUU���_UU����?�_UUUUU�_��UUU��?�?�UUUUU��?0�UUU��� ��UUUU���� _UUU������UUU���� �UUU��������U�U����  _UUU�������U������   �UUU���_��u�����?    WUUU��_��W���_��?    \UUUU�U�?\�_�W��    pUUUUUU��pU��_U�   ��UUUUUU=WsU5�U�   �?_UUUUU5\}U\�U�� ���UUUUU�pUUW�UU�� ��_UUUUU_UU���U� ���<�UUUUUUUUu5pU� ������UUUUUUUUU�_UU���� �WUUUUUUUUUUUU������_UUUUUUUUUUUU� ��?�UUUUUUUUUUUU � � �UUUUUUUUUUUU  �3��UUUUUUUUUUUU5  3�� ��UUUUUUUUUUU�5  �03��UUUUUUUUUUU�� �03  ��WUUUUUUUUUU�U�  ���WUUUUUUUUUUUW�  ��_UUUUUUUUUUUW5  ��U�UUUUUUUUUUUW5 � �U��WUUUUUUUUUW� ��\U����UUUUUUUUU]U�0�U]=�WUUUUUUUU]U30? �U]5�?WUUUUUUUU]U0<�\WW���WUUUUUUUU]U�0<�W]W��WUUUUUUUUUuUW���U�U��\UUUUUUUUUu�U��_UUU�7pUUUUUUUUU�uU��UUU��pUUUUUUUUUU_UU�UUUWUUUUUUUUUUUUU3�UUU5\UUUUUUUUUUUUUU��WUU�WUUUUUUUUUUUUUUWUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUU5 WUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUUU�pUUUUUUUUUUUUUUUUUUUU_UUUUUUUUU1U� ���><N�O OUL  �(                                                                              UU                                    @UUU                                   @UU                                   UUU                                   PU    TUUUUUUU                        UUI                                 PU`@��                                 TUTU�                                @UDY���                                PU�Ei*��                               UiY��*�                              @UTiAe��                              PUU�T
��            @                  TUAP�U���@UUUUUU   @                  UEEU���         T  @                 @UV�QV	TQR         @ @                 PU��AUPTZ                            TUTj�                             UeY��FUU%           @                @���AVZ��V                            @UUUUZPT                            PUUA�VUTUQ                            Td��PAUUe                            �Vei*�UUU                             UU�T�R�U                           @UZZ��Z�U�UU                           @���jUU�V                           P�UU���VUPUU           @                PU���>@UiTU            UUUUA@UUU       T��i��YT�YU                      @U   Ti����UUUUUU                            UU�Y��U�UZUU                            UUU�P�e�V�V                           U�V��`UUUUUU                           @��f_*ifUUUUQ                           @UUe�YjUUUUU          @               @AYUZY�VUUT                          @U���U�UQT           PU@UUUU        PU��XUUU�UAU                           P��U%UYVU�e�                           PY�VU��VUe%X                           PU��jU�V�U���                           PUUUYVU��U��                           Ti���%TUUU`�                           T�ViUejUUU*��                           T�WUUeU�VU嗯                           T�ij�Ye��U�*�                           TEe�jZYiUY���                           T���V�YeUU���                           ���ji��VVU���                           T囪iVU�����                           TQ�jU�UZ[���V                           T���ZUUUWeU��                           T��ZUUfU�UU�                           TU�����Z����V  TUU                     �ǚ�o�U��VUUi                           Tۛ������jYeU        TU                 T���i���VUUU                          P�gZj���iiVU                           Pʩ��Z����jU�                           P���V���UUU�                           P���������UUU                           @����oVUeU                           @}��i��ZYjUUU                           @U�����Uf�U                           @V�j����eVZUZ                  TU       �eUFi�jUYVU                            
��f��UZ��V                            Yw��^je�VUUU  @                        T�[X�jUUZUUU  PU                        �V��j�ZZ�
iU  U                       P�ֺ��ZjU�U  PQ                       PU�Z�ji���e  PU   @                  @e��jՐV�~�Z  PUP P                  @|�V�������  TUT T                   �ǧ�����V�j  DUPP T                   ����R����j[  TU T                   T�᪺�jV���  TUU DU                  P����UVj���  TUUUU UU          T      @UZ��e�kjj�  TUUUUEQU           @U     @U����V��  TUUUUUUU                  U��
Qii�  UUUUUUUUUT                  T����Z��Z�  UUUUUUUUUU                 Pe������V� @UUUUUUUUUUU                 @U�\��V���   PUUUTUUUUU                 U��Z�fU TUAUUTU  TUUU                Tee���ZZ�P    TQUU     T             P���z�U   TUUUP@UUUU                 UUb��ڥZ    @U                      TE��~)�k  @    U@                     PU�jV���  @ @U  U     @UU            U������   T  PUA     PU               T�k���         U                      PU����        @                        UU e�W     P    @UU                   PU�<��      P                           UUUe�       P                          @UU        U                          @UUU         PU               P          UU                           P                                      T                                     T                                     T                                     U                                   @Q U                                   @A U                                   PE@                                  PUAUP                                 PUAUT                                 TUEUUU                                @UUEUUUUU                              UUUUU PU                                PUUP                                PUUU U                               @@                                                                                                                        @UU                                  P                                     T                                     @                                                                                                                                                                                                                                                                               U                                     PUU                                    TVUU                                   UjUU                                  @�YU                                  P�UU�Y                           UU    ��VUPe                        UUUUU   �iUUUU                      @UUUUUUU  �eUUUUUU                     PUUU�jUU�ZUUUU�U             @U     TUUUUU��jU�UUUUUU�U            PU    @UUUU�����jEjVUUUUUUYUUU          TU  TUUU��������ZQ�UUUUUUUUTUUU       @UU PUU����������dUUUUUUUUUUe�jU      @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUU�(                                        U                                      AU                                     UU                                     @UU                                   DEUU                                    @U                                  �e PAU                                  ke T                                 �ZETA                                 �j(@UU                                 �VJFP                                ���HPU                                
 eV T                                VYEPQU                               @Y T P                               EY �F@      U                       TTD)�T         UUUUU  U             V �P HT                             T@U D�PP                @             UP �AA                             @P��                              APU-�U                              UQAI��
DT        PUUUUU              TQP���PU              T             UEI���j� P                            �UeZ�)�                            U�*���D               @            �Ua��
IPU              @             UZh�j T                            UU�ZU��~QU                           UUUIUR�6 @            @               UUEUU��_D                           UJU�                             UTTUU���WT                            TUAդ�                        PU P@�VUUUTT                             UEU�U����                            DUU��YUY�            @      PUU     E UUUUUe@PFT                           )@UUUZUYjZU                           V TU�UAA�EU            @UUUU         EUUUVU(AU                           �(P�UPUi�T                          �AUU�VPE`                          oTPU�U�VEU                          �QUUUUUe T                          j&�UUT�UaE                 @U      �&�QU�WUU�@T                          ZZ�UUUUZUiP            PU             7YZ�VUU��VU              T           �"�RUUU|Z�BP                           *ZUAUUUUVeZU                           �jZPUPUTU                           j�ZQUUUAUy�P                           kjUUU�UUUkUQ                           iUeUTUZI�VU                           eUEUUUU՗Q                           �UZUQUU�fT                            UUU_QyUUe�VU                            UYUUU��UVPUU                            UUUU�Z�U�UjU                            UU��UUUZZ�VU                            UU5UU`j�Z                            iUUUV�VekP                            TZ�WUUUPiAZ                            UUUhu���UU                            ZEe�eZUU�^                            �VUe�eVV�V                     @     UeU�ZX��kVU     T              @     �eUeUV��iVZ      PUU           P     i}VBd��gU                     P     UZUi�V�U�WU                      T     �������՗iU             PUU    P T     �VUY��UZ�U                    DAU     �VZiVjZiZY                    QUQ     �QZ���&��U                   @UUP    ZV����VfUZ                   PUUUUA   ժ�����֔U                  @UUUUTU   fze麯U�ZU                   PUUUUUUU   ef��XV�[�                  @UUUUUUUUU �ei��F�gZ                 TUUUUUUUAUU  Ze�_]���V             PU UUUUUUUUU    ��UV�f�_V                   UUUU TT  �k�����ZU                     UUU    @ �
��j�T`                 PU  @U      U��o��{U                   T         ���f*�U                    @U    UU �^��V}UU                      P @     ����a�V                       PPU      j���fUU                        U       �W�ZjVU                                 ���`UU                                 ��_�AU       P          PA            ��UU        P                        J�rWU        T           T           uUPU        T            T     P    TTU        T             U        UUU         U                T     UU        @Q U                        U         @A U                                   PE@                                  PUAUP                                 PUAUT                                 TUEUUU                             PU@UUUUUUU                            PUUUUUUUUPUU                          TUUUUUUUUUUUU                             @UUUUUUUUUP                            UUUUUUUUUU                         @UU  @UUUUUUUU                                @UQUUU   T@                         P  TTUU                            PU  TU @TUU TU                             @@U @                             @      P                                 @   U                               @   P                                    PU                                                                                                                                                            @                                              PU                             T     TUQU                              PU   UU@T                                  PU  P                                 PUPUT   UUU                          PU TUT @UUU                        PUTUUUTUUUUUU          @       PUUUU @UUUUPTU PU          UU      UUUUUUUUUUTUUPUU UU         PUUU    UUUUAUUUUUUUPUU�VUU AU        T@UUPETUUUUUUUUUUUUAUUjUUUET        UU QUUEUZUUPUUUUUUUUTU�jUUUEU       PUUU P�PUU% TUUUUUUUUUPUU���YUUU      TUU U�AUUUUUUUUUUUUUUUTU��ZUUUUU     UUU�Z*TYUUUUVUUUUUUUUU@U���ZUUUU    UUUE��JZUie�UYUUUUUUUUU PU��j�UUUUU   UUU����V�UUUe�VUUUUUU   @UE���jUUUUU  UUU����UVjZV�VUiUUUUUUU    ��ZZjUUTU  UUj��VY����jUUUUe�UUUUUUUUUU�������UPU U���VZ���������UUUUUUUUUUUU����jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU.
U�WUUU�UUUU=\U]U_UUU\uwWpUUU����p_UU �� ps]U ��  \ssU� �� �WssUU< �\ssUU� ��\ssUU   �\ssUU 3 �\ssUU�� �\ssUU<�\ssUU�< ��\ssUU�����pssUU? ?\�ssUU5   W�pUU����U5 \U��< ��� WU� p�_WU�� ��5W����3��5W�?� ��7W�� ��=_=< �� �p     � <s�?     �p0�  �0s0?  <�p��0 ���?s �� �5_��?���W5W50�� ��U5W�� ��U5WU�� ��U5WU����W5WU��<?W5WU�?<���U5WU��?�?W5WU��< \5WU  �  p5W�  �} �7W  pU  W  \U  0W  \U5  W���WU����W.UUUUUUUUUUUUUUUUUUUUU���_UUUUUUUU��?\UUUUUUU�  0 WUUUUUUU5 �UUUUUUUU�pUUUUUUUU� 0\UUUUUUUU�<WUUUUUUUU30 �UUUUUUUUU�  WUUUUUUU�  WUUUUUUU�   �UUUUUUUU5  ��UUUUUUU5   �WUUUUUU5    WUUUUUU5 �  \UUUUUU� ?  \UUUUUUU � WUUUUUUU   WUUUUUU�? ���UUUUUUU�� �_UUUUUUU�����UUUUUUU���?��WUUUUUU�?���_UUUUUUU?��UUUUUU� �0��UUUUUU�  ���UUUUUU50    WUUUUU50 �� �WUUUUU0 <  WUUU��?<�� �UUUU ��0�  |UUUU����? �_UUUUUU5����WUUUUUU��� �\UUUU��?�? ����WU�    033   \UU��?�������WUUUU�0??��sUUUU��?���0�UUUU  ?_� WUUU���  �   WUUUU�   7   WUUUU5   7  �UUUUU5   7  UUUUU�������UUU.UUUUUUUUUUUUUUUUUUUUU���_UUUUUUUU��?\UUUUUUU�  0 WUUUUUUU5 �UUUUUUUU�pUUUUUUUU� 0\UUUUUUUU�<WUUUUUUUU30 �UUUUUUUUU�  WUUUUUUU� WUUUUUUU0  �UUUUUUU��� ��UUUUUU��  �WUUUU�  �   WUUUU  <�  \UUUU �?  \UUU�  p � WUUU�  �   WUUU� ��? ���UUUU�  �� �_UUUUU �����UUUUUU ��?��WUUUUU5  ���_UUUUU�  ?��UUUUUU �0��UUUUUU=  ���UUUUUU�     WUUUUUU �� �WUUUUUU <  WUUU���� �UUUU ��0�  |UUUU����? �_UUUUUU5����WUUUUUU��� �\UUUU��?�? ����WU�    033   \UU��?�������WUUUU�0??��sUUUU��?���0�UUUU  ?_� WUUU���  �   WUUUU�   7   WUUUU5   7  �UUUUU5   7  UUUUU�������UUU0UUUUUUUUUUUUUUUU��UUUUUUUUU�7 WUUUUUUUU5 WUUUUUUUU0�\UUUUUUUU�0\UUUUUUUU� \UUUUUUUU� \UUUUUUUU5WUUUUUUUU5 �\UUUUUUUU� pUUUUUUUUUpUUUUUUUU�<\UUUUUUUU� 0sUUUUUUUUU0�UUUUUUUUU30�UUUUUUUUU��pUUUUUUUUU�\�UUUUUUUU5�� �WUUUUUU�_W��_UUUUUUU�� �_UUUUUUU5\��sUUUUUUU5\�?|_UUUUUU�s��uUUUUUUU�0��UUUUUU� �0��UUUUUU� 0|�UUUUUU� 00uUUUUUUU��_]UUUUUUU ��WUUUUUUU <wUUUUUUUU  \UUUUUUUU  pUUUUUUUU  pUUUUUUUU  \UUUUUUUU5  _UUUUUUUU5 �WUUUUUUUU���_UUUUUUUUU? pUUUUUUUUU �UUUUUUUU�   WUUUUUUU� 0 WUUUUUUU� 0 \UUUUUUU� 0 pUUUUUUU5 � �UUUUUUU50� �UUUUUUU5 �UUUUUUU����0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUWUUUUUUUU�� \UUUUUUUU=< \UUUUUUUU� sUUUUUUUU �pUUUUUUUU pUUUUUUUU� pUUUUUUUU\UUUUUUUU sUUUUUUUU 0�UUUUUUUU50�UUUUUUUU��0pUUUUUUUU� ��UUUUUUUUU� W�UUUUUUU�� � �WUUUUU�U��_UUUUU s� �_UUUUU�_U��sUUUUU5p_U�?|UUUUU�_�U��UUUUUUUW0�_UUUUUUW�0�uUUUUUU�\0|�UUUUUU�� 0�UUUUUU5 ��_uUUUUUU5 <��_UUUUUU5 �0wUUUUUUU�  \UUUUUUU�   pUUUUUUU�   pUUUUUUU�   pUUUUUUUU  \UUUUUUUU �WUUUUUUUU �WUUUUUUUU=��_UUUUUUUU� pUUUUUUUU�  �UUUUUUUU� 0�UUUUUUUU5 0 WUUUUUUU5 0 \UUUUUUU � \UUUUUUU0� pUUUUUUU pUUUUUUU����0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUU|UUUUUUUUUU�UUUUUUUUUU _UUU�UUUUU�pUU� �WUUU0�UUU��_UUU0 WU� �_UUU3 �\UU��sUU��0pUU�?|UU5 < �UU��UU5 ��WU0�UU5 <0\U�0�_U�� �\U0|uUU? <W� 0�UU�� ��U��_�UUU?� W=�W�UUU�?�W0WuUUUU��|��_UUUUUU�� pUUUUUUU5   pUUUUUUU5   pUUUUUUU5   \UUUUUUU�   WUUUUUUU�  �WUUUUUUU�  �_UUUUUUUU� pUUUUUUUU= �UUUUUUUU� �UUUUUUUU�  WUUUUUUU5  \UUUUUUU5 � \UUUUUUU5 � pUUUUUUU50 pUUUUUUU����0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUU5��UUUUUUUUU�0�WUUUUUUUU5��WUUUUUUUU���\UUUUUUUUU�_UUUUUUUU� �UUUUUUUU� ��UUUUUUUU�<_UUUUUUU� _uUUUUUUU5 �_�UUUUUUU�<�W�UUUUUUU�<�U�UUUU�UUU�UuUUU� WUU�W_UU� \}� �UUU��   pUU� �p�   pUU p=   \U� ��p5   WU�   _�  �WU� �  W�  �_UU��UU� pUU�  sUU= �UU5� \UU� �UU5� WUU�  WU �UUU5  \U |UUU5 � \U5 WUUU5 � pU5�UUUU50 pU�_UUUU����U���W�U���_�U����U��p�U�  �U���������?�����?w����?w����?w�����wU����uU���uU5��\uU�  _]U���]U���]�����W�����_����?p3�0p����\���_���u� p5 WUp��UUpUUUU�_UUUU���WUU���_�U����U��p�U�  �U���������?�����?w����?w����?w�����wU����uU���uU5��\uU�  _]U���]U���]�����W�����_����?p3�0p����\����_��=�u��5 WUp5�UU�_5�UUUU�UU�uU�u���}���]���]���_U�WU�_WUpWU��W���W�?�W�?�W���U�pUU_UU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �(  DUDUD
 �QUUU P  �   �
P P P P *   D� Q
QUU P ��������������������*  �  T U P ��jUUU�  D�ZUUUUUUUUTU����*�  Q  P ��jUU   �����"          TUUU���  T�
@���VUU     �����
              TU�   ���jUU       �����"                �����ZUU          �����
                �  D�"            �  D�"        *       �����
        ��������������������*     �����"      ���UUU�  T��UUU�    % ����* �����
    ��* � �  �� �    %   `U�������" ���   �UU�  T��AU�    *   `UUU�  D����UU   �� �  Q�� ��    *   `U  ������UUQU   ��V�  T��T��        `UE�  T�� UU     ��  Q���*      � ��@�  ��U��      �  ��%         ��UA�  T��U��      �  Q��%       �  ��E�  Q���*   �   V�  T��Q%            �E�  T��Q	    �    j�  Q��U*       �   ��  Q��Q	        h�  T��Q
          �U�  ���
       h�  Q��U
      �    �Z�  Q���         h�  T��U
������       Z�  T���    � �   ��  Q���TUUU  �   Z�  Q���          �  T�� ���������   Z�  T���         �  Q�
 �      ����*  ��  Q��          �  T�" ((UUUUU���j   �  T��*   � ���  �  Q�
 
UUUUUR  X   �  Q��    �����  �  �" �BUUUUURUUU   �  �
    ����   �  Q�
��PUUUUURUUi   �  Q�"    %  P�   �  T�"��TUUUUURUUi   �  T�
    $UUU�   �  Q�
)TUUUUURUUU   �  Q�"    $UUU�   �  T�"�
UUUUUURUUe   �  �
    $UUU�   �  Q�
�@UUUUUURUUe   �  Q�"    $UU�   �  T�"�TUUUUUURUUU   �  T�
    $UA�   �  Q�
�TUUUUUURUUe   �  Q�"    $U@�   �  �"�TUUUUUURUUU   �  T�
    $UP�   �  Q�
�TUUUUUURUUe   �  Q�"    $UT�   �  T�"�TUUUUUURUUU   �  T�
    $UQ�   �  Q�
�TUUUUUUPQU   �  Q�"    $UA@�   �  T�"�TUUUUUU PU   �  �
    $U �   �  Q�
�TUUUUUUR@UU   �  Q�"    $UD�   �  T�"�TUUUUUURUUU   �  T�
    $UP�   �  Q�
�TUUUUUURUP   �  Q�"    $UT�   �  T�"�TUUUUUURU@   �  T�
    $UU�   �  �
�TUUUUUURU @   �  Q�"    $UU�   �  T�"�TUUUUUURUT   �  T�
    $UU�   �  Q�
�TUUUUUURUUU   �  Q�"    $UUU�   �  T�"�TUUUUUURUUU   �  T�
    $UP�   �  Q�
�TUUUUUURUUU   �  �"    $UQQ�   �  T�"�TUUUUUURUUU   �  T�
    $UQ�   �  Q�
�TUUUUUURAUU   �  Q�"    $UP�   �  T�"�TUUUUUURUU   �  T�
    $PP�   �  Q�
�TUUUUUURUU   �  Q�"    $ Q�   �  T�"�TUUUUUURUU   �  T�
    $UEA�   �  �
�TUUUUUURUT   �  Q�"    $UUQ�   �  T�"�TUUUUUUR UP   �  T�
    $UAP�   �  Q�
�TUUUUUUR TP   �  Q�"    $UT�   �  T�"�@UUUUUURA@P   �  T�
    $UUT�   �  Q�
�
UUUUUUD P   �  �"    $UT�   �  T�"X)TUUUUU@   �  T�
    $UUU�   �  Q�
��TUUUUUU@   �  Q�"    $UUU�   �  T�"��PUUUUU  @   �  T�
    $UUU�   �  �
 �BUUUUURU    �  Q�"    $U �   �  T�" X
UUUUUPUU   �  T�
    $ �   �  T�
 h)UUUUURQP   �  Q�"    $�   �  �" �%     RUUU   �  T�
    $@�   �  T�
 �������RUUU   �  �"    $ U�   �  Q�"  VUUUUURUT   �  T�
    $UU�   �  T�
  ������RUT   �  �"    $Y@�   �  Q�"        RUU   �  T�
    $YD�   �  �
        RUUU   �  Q�"    $UA�   �  Q�"         PU   �  T�
    $iUU�   �  T�
        ��    �  Q�"    $iUU�   �  Q�"        ����*   �  �
    $U �   �  T�
        U���j   �  Q�"    $ ���  �  Q�"         PUUU   �  T�
    �����  �  T�
                �  Q�"    ���VU   �  Q�"                �  T�
    UUU    ����
�                �  Q�"            � ��*(               �  T�
            (Te���               �  Q�"            U����               �  �            JUU���               ����*(           BU����               � ����           RUU���               (Te���           RU����               U����           RUU���               JUU���       ���*RU�������������*��
   BU����     ��*   RUU���       �� ���RUU���   ��*  ��*RU��������������
�   *RU�������
  ����*RUe�������������*���* RUU�����  �������*BU��������������*����*RU����( ���������*
Ue�����������)�*����*RUe���������������(U������������)�*����*BU��������������������*���������)�*����*
Ue������������                ��
 ����(U����������� @UUEUUUUUUUTUUUQ��BU   �����������  PQUUUE@QUQUUDUU�*PUUU      ���* PUUUUUETUUQUUUDUUU�jUUQUUUEUUU!  UTUUUUUUETUUQUUUDUUU�jUUUUUE@TUQUUUDUUUUUEUUUUUUUTUUUQ�jUUUUUUETUUQ@TUDUUUQUUUEUUUUUUUTUUUQ�jQUUUUUUETUUQTUUDUUUQUUUEUUUUUUUTUUUQ�jQUUUQUUUEUUUQTUUTUUUQUUUEUUUUUUUTUUUQ�jQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�jQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�jQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�jQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�jQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�
                                      �VQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�UUUUUE@TUQ@TUDUUUUE@TUQUUDUUjUUUUUUUETUUQTUUDUUUUUUETUUQUUUDUUUVUUUUUUUETUUQTUUDUUUUUUETUUQUUUDUUUUUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQZUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�UQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�VQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�ZQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�                                      �VQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�UUUUUE@TUQ@TUDUUUUE@TUQUUDUUZUUUUUUUETUUQTUUDUUUUUUETUUQUUUDUUUdUUUUUUUETUUQTUUDUUUUUUETUUQUUUDUUU�UQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�UQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�UQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�UQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�UQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQjUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQUUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQUUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQUUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQUUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQUUQUUUQUUUEUUUQUUUTUUUQUUUEUUUUUUUTUUUQ�(                        @ UU P                                @ U  @                               PE    PU                             P  PUTUA                            @@E   UU                             @ AUU PE                              PAUU P                    @UUU      PU@ PT                    T         @U   PU                    T   PU      T  PU                     TU @     @UPUUU                     T         UU@U                    @  P  @U    @U                       T@  @TQU                             U   TU                              UU @U                              @TUT@                               @U U @Q                                U   @U                                P  @U                                  UAUUU                                  TUU                                    U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      T                                     @U                                    PU                                    TU                                    UU                                    TU@                                 @U UU@                                 @UUP                                 @AUUP                                 PAUUP                                 PAUUT                                 TUAUUT                                 TUAUUT                                 TUQUUT                                 TUQUUT                               @UUUQUUU                              UUUUUUUUUU�                           @UUUUUUUUUUU�  ��                      @UUUUEUUUUU�*�
                         UUUUUUUUi��%��A                         @UUUU)�j%��                        TPDUQUUh�%��U PUUUUUUAU          @UU    	�Z%��                      UUTUUUUUUUUU AUeUUUUUUUUUUUUUUUUQTUUUUUUUUT        `JUUUUUU PTUUUUUUUU   @TUUUUUUUU  DaFUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUUEA`VUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUFDDhVUUUUUUUUUUUUU@UUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUDUUUUUUUQUUUUUUUUUUUUE�hUUUUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUTV�`UTUUUUUUUUUUUUUUUPUUUUUUTUUUUUUUUUU�`UUUUUUUUUUUUUUUUQUUUUUUUUUUUUUUUYE�hUUUUUUUUUUUUUUUUUUPUUUUUUUUUUUUUUUUU�VXUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUZU�XQQQQQQQQQQQQQQQQQQQQUUUUVU�ZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUVU�UQQQQQQQQQQUUUUVU�VDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUQQQVU�DDDDVEURUUUUUUUUUUUUUQUUUUUUUUUUTUUUUUUUUUVUUVUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQVTTTTTTTTTTDEEEEEEEEEETTTTTTTTTEEEEUUUVUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUFEEEEEEEEEEUTTTTTTTTTTEEEEEEEEEETTTTUUU�UeUUFDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDUaUUUQUUF@@@@@@@@@  DD @  @@  UQUU                     �       (   U@UU    @@@@@    A  @ A     UdU                     �  �Q�  (  UTUV                     � jUU�P
    UPUV                      ZUUUUUU�    U`U                      ��������     UaU�                      �eYf�$I    U�U�                      �e�f�$I    U�U��                      �i�eX��)    U�U��                    ��fY�aX�%	   U�U��                     �iY�aX�� P U�U��                    ��Y��aX�� U�U��                    ��Z��aX��
P UaV��                     ����������    U�U��                      PEQEQ     aU��                    ��ZU�jU�Z)    UaU��                      �iU*�V�i   U`U��                     i��V Zi�   UaU�U                     %`�U�%`   U`U�                    �h��
��h�   UhU�                   ��ZY����Z�   UhU�                   ����ZU���J	   UhU�                    ���X�����X   U�U�                    ����������PUUhU�                   �������j  T�U�                   h����VXXXX� UUh`U�                   Z����Vhhhh�V ``UU                  �VhaaaVaaa�Z  ``U                  �ZhhaVa���V(  ``U                  `�VXXhV���Z!  `aU      T           h�ZXV���VX�  `aU      D         ��Z��VXV�Zh�
�`aUA      T         ��U`��Z�Z�Zha�`aUA                
�jh�V�iVX��V��haU@               * 
� h� (���XUU �   U           �����������������*XUU��  @U           �����������������
XUU�%    U            bff""""""""""ff&XEU�%  @              ���B�VPPU�!��� XE�%                  HUUQ�U AU�UU� XUT�                  ���T�UUAT�U��� XUT�                �b�U�VUPEQZU)f�XUT�      U        �@�UZUUUU�VT
XUT�  @ @U         �P�V������  
�*XU��  PU  U         "T�V�     
 Be*TU��  @            "U�V�������* R�*TU��         @      b�j�������
�V`*TU��           U     b���   � ��*TU h�          @U     b��(���*� d*TU X�          U     b@��h  �� �*UU Y�                "P���ZUUU�Be*UU Y�     @          "T����UUUU	�R�*UU X�     PU          "U���UTU)
�V`*UU Z�     @          b���fUPU%�*YU V�                 b��fUPU
d*
UU�V� P               b���fU@U�*
ZU�V�             T �b@���fU�JU
(Be*
VU�U� P       @@UUA�"P�j�fU��U
 �*JVU�U�                U�"T�V�fU��U
 `*XV�U�               EA�"�V�f    
 � V�U$              PUU�b�V�f    
TUUUU4UUUUUUUUUUUU���UUUUUUUUUUUUUUUUU  �WUUUUUUUUUUUUUUUU ? \UUUUUUUUUUU����U5 �pUUUUUUUUUUU����_�  ��UUUUUUUUUU������U �WUUUUUUUUU�??��W= �?\UUUUUUUUU�?� �_� �_UUUUUUUU��  �U= �UUUUUUUU����� �W����UUUUUUUU������UU�WUUUUUUU������� �UU��WUUUUU�W�������?�_U��_UUUUU��� �������U��UUUU������_����WU�UUUU������WU������UUUU����� �U���  ��UUUU�����  U�����UU�W�����  �W��?���UU������    |�����sUU���U���    ��?� �OUU��U��?    ���?���_�_U��? ��? ��������sU�UU�? ��? ������������UU� ��� ��W������5p�WU� ��� ��_=���5\WUU ��� ���__��U5WWUU <? �W��sU�W���UUU �<� �W��U�\UUUUU5 ���3 W��Us5\UUUUUU5  ��� W5p�U��_UUUUUU5 �����W��UUWUUUUUU�� 0��3���?WU�UUUUUUU�� � �<���\UUUUUUUUU��  �����s5\UUUUUUUUU�� ��0����_UUUUUUUUU�U0���WUUUUUUUUUU�U0 <���UUUUUUUUUUUUW5�0 �p�UUUUUUUUUUUUUW5 � �p�UUUUUUUUUUUUUW5����s�UUUUUUUUUUUUUW�0��<suUUUUUUUUUUUUUW����\uUUUUUUUUUUUUU]U��?_uUUUUUUUUUUUUU]�=��u]UUUUUUUUUUUUUuu����WUUUUUUUUUUUUU�_U5<�UUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUUU\UUUUUUUUUUUUUUUUUUU�WUUUUUUUUU<UUUUUUUUUUUU��UUUUUUUUUUUUUUUUU�  �_UUUUUUUUUUUU��WU � 0UUUUUUUUUUU����W5 �?�UUUUUUUUUU�����  �WUUUUUUUUU�����W �?\UUUUUUUUU�?<� �=  �sUUUUUUUUU�  ?�� �UUUUUUUUU� �? �W= ��UUUUUUUU���������WUUUUUUU�� ���?��UU��WUUUUUUU��������_U��_UUUUUUU�?�����?��UU��UUUUUUU�?��W�����WU��WUUUUUU�?��U��� U��_UUUUUU�?<�UU�����W=�_UUUUUU�?0�WUU�� |��_UUUU�?0�WUU��� ����sUUUU�� �_UUU������pUUUU���UUU��?����sUUU�_���UUU�����]UUU���?��WUUU��?�_��UUUU����� |UUU����W�WUUU����� �WUUU���W�5\UU�����3  |UU���U��\UU�����?  �W��U�UW_�_�����  |��WUUU5\U5��_�����?���WUUU�WU��W�����? ��_UUUUUU��U������ ��UUUUUU��UU����� ���UUUUUUU��UU�?��� ���W�UUUUU��WUU? <? ���?WUUU���_UU= �<� �_��?\UUU�p5\UU5 ���3�W���\UUU�\\UU5  ����UUW_UUUUWWUU5 �����U�_UUUUUU�UUU5 0��3 W��sUUUUUUUUUu5 � �< W���UUUUUUUUUu�  ��� W7W�UUUUUUUUU�� ��0 W7\�UUUUUUUUU�� 0� W�pUUUUUUUUUU�U0 ���U_UUUUUUUUUU�U �  ��UUUUUUUUUUUUUW�  �p�UUUUUUUUUUUUUW5 ?��_�UUUUUUUUUUUUUW5���<W�UUUUUUUUUUUUUW�0���_�UUUUUUUUUUUUUW�� w�UUUUUUUUUUUUU]U�?�uUUUUUUUUUUUUU]�=��U_UUUUUUUUUUUUUu}�7��UUUUUUUUUUUUUUU�WU5�?WUUUUUUUUUUUUUUUUU5��UUUUUUUUUUUUUUUUUU�<�UUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUUU\UUUUUUUUUUUUUUUUUUUWUUUUUUUUUUUUUUUUUUU�UUUUUUUUUU?UUUUUUUUUUUU��UUUUUUUUUUUUUUUUU�  �_UUUUUUUUUUUU��WU � 0UUUUUUUUUUU����W5 �?�UUUUUUUUUU�����  �WUUUUUUUUU�����W �?\UUUUUUUUU�?<� �=  �sUUUUUUUUU�  ?�� �UUUUUUUUU� �? �W= ��UUUUUUUU���������WUUUUUUU�� ���?��UU��WUUUUUUU�� �����_U��_UUUUUUU�������?��UU�UUUUUUU����W�����WU�UUUUUUU����U��� U�UUUUUUU��0�UU�����W=UUUUUUU�� �WU��� |�UUUUUUU�� �WUU��� ��UUUUUUU���_UU������WUUUUUU��UUU��?���WUUUUU�_�?�WUU�����_UUUUU���? |UUU��?��_UUUU�����  �WUUU����_�WUU�����   |UUU�����\�_�����   �UUUU����?\5��_��?   WUUU��W��\��W��? ��?\UUUU�U�_W��U��? ��?pUUUUUU�U��UU� ����WUUUUU��UU��UU� ��� UUUU�WU��WU� ��� �WUUU�s5W���_UU <? �_UUUU��W�p5\UU �<� �UUUUWU�\\UU ���3��UUUU�UUUWWUU  �����WUUUUUUUU�UUU ������_UUUUUUUUUUUU 0��3��_UUUUUUUUUUUU5 � �< �sUUUUUUUUUUUU5  ��� �sUUUUUUUUUUUu� ��0 �sUUUUUUUUUUUuU0� ��UUUUUUUUUUUuU0 � ��UUUUUUUUUUU�U �  ���WUUUUUUUUUU�U�  �p��WUUUUUUUUUU�U5 ?��_U�_UUUUUUUUUU�U5���<WU���_UUUUUUUUUW�0���_U���sUUUUUUUUUW�� wUW��UUUUUUUUUWU�?��U��UUUUUUUUUW�=��U�U5p�UUUUUUUUU]��7�U}U��UUUUUUUUUU]uU5�_UUU�?WUUUUUUUUUu]U5�_UUU�\UUUUUUUUU�WU5�_UUUs5\UUUUUUUUUUUU��UUU��_UUUUUUUUUUUU���UUUWUUUUUUUUUUUUU�?WUU�UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUU5pUUUUUUUUUUUUUUUUUUU5\UUUUUUUUUUUUUUUUUUU�WUUUUUUUUU7UUUUUUUUUUUU��UUUUUUUUUUUUUUUU�? UUUUUUUUUUUUUUU�  �UUUUUUUUUUU���UU< WUUUUUUUUUU���_U�?\UUUUUUUUU����U5 �pUUUUUUUUU��< �W� ��UUUUUUUUU�? U �UUUUUUUU�� < �U� �WUUUUUUU�����_U��WUUUUUUU���� �UU�WUUUUUUU������ �W��WUUUUUUU������5�UUUUUUUU��������_UUUUUU����_U��<���_UUU�����\U�������sUUU����0|UU�� �����UUU����|UU����_���UUU����|UUU���_��UUU�����UUU���W��UUUU�����WUUU�_U�WUUU����?�_UUUUUU�\UUU����� UUUUUUs5\UU����� UUU�UU��_UU��W����UUU�WUWUUU��U����_���UU�UUUU�_UU��?���UUUUUUU�WUU���  ��UUUUUU��UUU�� ����UUUUUU�UUU�� ����WUUUU��_UUU� �?��_U�_U���UU�0<� �_U�_U����UU� �� � |��sU����UU�     0�p pU���UU5     0� \U�\�UU5     �� �WU�5\sUU��     �WUu5\]UUU   0  _�UUU5WUUUU50    �U}UUU�UUUUU5�   �pUUUUUUUUUUU   � �_UUUUUUUUUUU   0 �_UUUUUUUUUUU   0 �UUUUUUUUUUU�  �  �UUUUUUUUUUUU�   � �WUUUUUUUUUUUU?  ��_UUUUUUUUUUUU� ��UUUUUUUUUUUUU��U5 �UUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUU|UUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUU_UUUUUUUUUUUUUUUUU�UUUUU���U���U����U����U �����������w����w����w����uU���uU��_uU p]U��]U���]���]����W����_� ��p����s�����WWUW�UU�UUU          �(Z)YU� �jd�Re���V�� @VjEA�ZP�������Z)YU� hj��Re���V�� P�jU�����������ViYU� hjj�Re`�jZ�� @V�Z����U������UiYU��hjEZ�Reh�Zj�� Pf��VY���������U�UU��jjEZ�Re!h�ZjZ�
 T�U����V�������U�UU��j�UV�Re Y�V�V�F�d��U���Vi�V���*�U�UU`�j�V�bU`Z�V�V�V� ��jU�ZVUi����Z�U�UU`�j�V�bU`V�Z�V�V� ��jUUjZUi����V�U�UU`���%V�*�V�Z�V�V��d�ZUUjVUe�Zf�V�U�TU ����V�*`U�Z�V�Z��d�ZUUjVUUUZj�V`U�TU h���U�*`U�Z�V�Z�f�ZUU�VUUUZV�V`U�TU*X��fU�*`U�Z�VUZ� j�VUU�VUUUj	��V`U�PUX��jU�*aU�ZUUUi�VUVUU�UUUUjI��Z`U�XUXi�fUU*aU�VUUU��VUUUU�UUUUjiV�Z`U�XU
Xe�jUU
VaU�UUUU�VUUUU�UUUUjaV�ZhU�XUXU�jUU�FbU�UUUU��VUUUUUUUUUj�V�ZXU�ZUXU�ZUU�FbU�UUUU��UUUUUUUUUU�eUUjXU�ZUXU�ZUU�JjUUUUUU�FdUUUUUUUUUU�eUUjZU�ZUXU�VUU��VUUUUUU�FdUUUUUUUUUU�fUU�ZU�JU�XUUUUU��VUUUUUU�VhUUUUUUUUUU�jUU�&VU�JU�XUUUUU��VUUUUUU�VXUUUUUUUUUU�jUU�&VUUJU�ZUUUUU��UUUUUUU�ZXUUUUUUUUUU�jUU�&VUU�U�UUUUUU��UUUUUUU�ZXUUUUUUUUUU�jUU�&VUU�U�UUUUUU��UUUUUUU�jXUUUUUUUUUU�ZUU�&VUU�T�UUUUUU��UUUUUUU�jYUUUUUUUUUU�ZUU�&VUU�T�UUUUUUUjUUUUUUU�jYUUUUUUUUUUUVUU�*VUU�T�UUUUUUUjUUUUUUU�jXUUUUUUUUUUUUUU��VUU�U�UUUUUUUiUUUUUUU�jYUUUUUUUUUUUUUU�fUUU�U�UUUUUUUYUUUUUUU�jYUUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUUjYUUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUZUUU�TYUUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUZUUU�TZUUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUZUUU�XVUUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUU�VUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUU�VUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��FUUUTUUUTUUUTUUUTUUUTUUUTUUUTUUUTUUUQT��VTUTUTUTUTUTUTUTUTUTUTUTUTUTUTUTUTUTEEE�EEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEETTT�TTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTT*DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                                   ���                                   �Z *                                  �V  �
                                 X    �                                �     �
                               �     T�
                              �     U �                             �     U  
                            ��A   PU  (                           ���UU  TU  �                           jU��UUUUUU  �                         �V  �ZUUUU�  @
                        �j  �ZUUUU�U@)                        �U   �jUUU�ZU �                        Z   TjUU�VUU �                      �    P�UUUUUU T
                      �    P�ZUUU�UU P)                      `    P�jUUU�UUP�                      h     PP�ZU��UUP�                     X     P�����UUTU                          T����jUUUUT
                          T����ZUUUU@)                         @UV���VUUU �                        TU@UVU��VUUUU �                       PUUTUVUUUUUUUU�                      T UUZUUUUUUUUT                      UUUUZUUUUUUUUU                   � @UTUU�VUUUUUUUUU                   � @UUUU�VUUUUUUUUU�              ��� h @EUUUZUUUUUUUUUU�               Z���Z @QUi�VUUUUUUUUUU�              �  ��UU PUUU�UUUUUUeVUU��              �  P�ZUPUUVjUUUUUEU�UU��              h   U�UUUUUVZUUUUUZ�UUi%              X    U��UUUU�ZUUUUU�UVUZ*                  T��ZUU��ZUUUUU�V���
                  P�VjUUi�ZUUUPUU�Z���
                  P�V���V�ZAYUPUU�j�Z�                  T�Z��j��V�U@UU��UU�      ��*         U�ZZ�j��V�VPUA��j��       �Z�       PEUUZ�VU��U�VPU ����*       ZU�*   � @UUUUZU�V�jU�V@U ����*      �TU�   � @UUU�VU���ZU�@ ����*      j@U�*  �V PUUU�VUU��UUA�P ����
     �V  UT� �UUUUU�VUU�jUUE�TP����     h  T �* �UUUUUU�VUUUUUUE�TT����     Z   T��*��UUUUU�UUUUUUPE�TTP����*   �   P�����jUUU��UUUUU @�VQP ��jU�  �   PP���U��UU�jUUP @�VEUU @UU@�
  h   @P��jU���Z�jUU    P�jTU     �*  Z    @UP��jUUU���ZU    P��U@U    @�� �    @UQ��ZTU���UU    T��ZU    PU�
�    PU��V PU��ZUU    T��jU    T��*�    PU��  UU�VU     TUP��VU   PU����    TU��  TUUUU     TUQ��ZU   TU���Z     TU��  PUUU      TUU���Z  UY��Z    @UU��  @UUU      TUE����U  UY��V     UUU�j  @UUU      PUE����U@UU�j    @UUUE�j   @UVU       PUE��Z�UUUU��V    @UUUE�j   PUZU       PUE��j�UUUU��     PUUUE�j   PUjU       PUU��jUUUU���     TUUUE�j   PUiU       TUU��ZUUUU��j     TUUUU�j   TUiU     @UU���VUUU��j     TUUUU�j   TUiU     PUU��� UUUe�j      TUUU�j   TUiU     TUU��j UUUe�Z      TUUU�j  UU�U     UUU��Z UUUi�Z      TUUUU��  UU�U     @UUU��VUUUU��Z   @ UUUUU��  UU�U     PUUU��V UUU���Z   @U@UUUUU��  UU�U  UU UUUU��@UUU���Z   PUUUUUUU��  UU�UPUUUUUUU��PU�����Z  TUUUUUUU��V@UU�UTUUUUUU��jPU�j���ZP UUUUUUUUU�VUUU��UUUUUUUUU��jPUUiU��ZUUUUUUUUUUUU�ZUUU��UUUUUUUU��ZPUjU���ZUUUUUUUUUUUUjZUUU��TUUUUUUU��ZTU�V���ZUUUUUUUUUUUU�jUUU��TUU�ZUU���VTU�����ZUUUUUUUUUUUU����U�jTUU�jUU���VUU�����ZUUUUUUUUUUUUi�����ZQU����VU���UUU�����ZUUUUiUUUUUUUi�U���Ve�����jU���UAUU�����ZUUU�UYUUUUUU��Z�����ZUU�����jUPUU�����ZUUUiUUUUUU��j��U��V�ZUP�����VTUU�����ZVU�Z�ZUUUU��j��UUjUUUUUQ����jU@UUU�����VVUi���VUU���V��UUUUUUUU����UUUUUU��������Z���jUU��U���VUUUUUUUT��ZUAUUUi��������V����V��j����ZUUUUUUUU@�VUUUUUU�����V�������Z�������jUUUUUUUUTUUU��UUU�����ZUU��������������UUUU    UUUUU����������jU���������
   ��ZU�UU @TUUUU������ �   ��������� �����* @   ����*      ���
 ��������  ��
�                    ��*  ������*      �                          U����                                 TQ                                    @UU                     @U             @��                     @@ PU    U  @�V        UTU        @TV@  @�   U   PUUUUU            @�T@  @d                           TA�P �(i� ��ZU�iZ)YU� �jd�Re���V�� @VjEA�Zi� ��ZU��Z)YU� hj��Re���V�� P�jU���i� ����j�ViYU� hjj�Re`�jZ�� @V�Z����� �Y��UUUiYU��hjEZ�Reh�Zj�� Pf��VY��� �i�jUUU�UU��jjEZ�Re!h�ZjZ�
 T�U�����U� ��jUUUU�UU��j�UV�Re Y�V�V�F�d��U����U! ��ZUUUU�UU`�j�V�bU`Z�V�V�V� ��jU�ZV�U! i�ZUUUU�UU`�j�V�bU`V�Z�V�V� ��jUUjZ�U! Y�VUUUU�UU`���%V�*�V�Z�V�V��d�ZUUjV�V% Y�VUUUU�TU ����V�*`U�Z�V�Z��d�ZUUjV�V�Y�VUUUU�TU h���U�*`U�Z�V�Z�f�ZUU�V�V%�Z�UUUUU�TU*X��fU�*`U�Z�VUZ� j�VUU�VUZ$�U�UUUUU�PUX��jU�*aU�ZUUUi�VUVUU�UUj$�UUUUUUU�XUXi�fUU*aU�VUUU��VUUUU�UU��UUUUUUU�XU
Xe�jUU
VaU�UUUU�VUUUU�UU��UUUUUUU�XUXU�jUU�FbU�UUUU��VUUUUUUU�iUUUUUUU�ZUXU�ZUU�FbU�UUUU��UUUUUUUU�YUUUUUUU�ZUXU�ZUU�JjUUUUUU�FdUUUUUUUU�TYUUUUUUU�ZUXU�VUU��VUUUUUU�FdUUUUUUUU�TZUUUUUUU�JU�XUUUUU��VUUUUUU�VhUUUUUUUU�TVUUUUUUU�JU�XUUUUU��VUUUUUU�VXUUUUUUUU�VVUUUUUUUUJU�ZUUUUU��UUUUUUU�ZXUUUUUUUU��VUUUUUUUU�U�UUUUUU��UUUUUUU�ZXUUUUUUUU��VUUUUUUUU�U�UUUUUU��UUUUUUU�jXUUUUUUUU��VUUUUUUUU�T�UUUUUU��UUUUUUU�jYUUUUUUUU��VUUUUUUUU�T�UUUUUUUjUUUUUUU�jYUUUUUUUU��VUUUUUUUU�T�UUUUUUUjUUUUUUU�jXUUUUUUUU��VUUUUUUUU�U�UUUUUUUiUUUUUUU�jYUUUUUUUU�jVUUUUUUUU�U�UUUUUUUYUUUUUUU�jYUUUUUUUU�jVUUUUUUUU�T�UUUUUUUUUUUUUUUUjYUUUUUUUU�jVUUUUUUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUUjVUUUUUUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUU�VUUUUUUUU�T�UUUUUUUUUUUUUUUU�ZUUUUUUUUU�VUUUUUUUU�TYUUUUUUUUUUUUUUUU�ZUUUUUUUUU�VUUUUUUUU�TZUUUUUUUUUUUUUUUU�ZUUUUUUUUU�VUUUUUUUU�XVUUUUUUUUUUUUUUUU�ZUUUUUUUUU�UUUUUUUUU��VUUUUUUUUUUUUUUUU�VUUUUUUUUU�UUUUUUUUU��VUUUUUUUUUUUUUUUU�VUUUUUUUUU�UUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUTUU��FUUUTUUUTUUUTUUUTUUUTUUUTUUTUTUTUTUTQT��VTUTUTUTUTUTUTUTUTUTUTUTUTEEEEEEEEEEEEE�EEEEEEEEEEEEEEEEEEEEEEEEEETTTTTTTTTTTTT�TTTTTTTTTTTTTTTTTTTTTTTTTT*DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                                                                                                                                                                
                                       �         
                             �
       ��
                            �	      � �                           �	     �   
                           Z�*    
    (                           ZY�*  �    �                           �ZU�� �     �                         ��UUU�
h  @  @
                        �j�UU���  @U@)                        �U�UUU�V TUU �                        ZjUUU�j UUU �                      � jUUU�j@UUU T
                      � ZUUU�j@UUUU P)                      ` VUUU�j PUUUUP�                      h  UUUU�j TUUUUP�                     X  UUUU�Z TUUUUTU                       UUUU�ZUUUUUUUT
                       UUUU�ZUUUUUUUU@)                       UUUU�ZUUUUUUU �                       UUUQ�ZETUUUUUU �                       UUUU�V@UUUUUUU�                      UUUQ�V@UUUUUUUT                      UUUQ�PUUUUUUUU                   � @UUUT�TUUUUUUUU                   � @UUT�UUUUUUUUU�              ��� h @UU�jUUUUUUUUU�               Z���Z @UU�jEUUUUUUUUU�              �  ��UU PAA�ZAUUUUeVUU��              �  P�ZUP  P�VQUUU�U�UU��              h   U�UUU D��UAUUU�Z�UUi%              X    U��UUPU�jUQUUU��UVUZ*                  T��ZUUU�ZYQUU���V���
                  P�VjU��jUiUUU���Z���
                  P�V��UUUU�UUU���j�Z�                  T�Z��UUUU�UU�����UU�      ��*         U�ZZ�@UUU�ZU�����j��       �Z�       PEUUZ�V UUUU���������*       ZU�*   � @UUUUZU�UUUU��j������*      �TU�   � @UUU�VU�UUUUU���������*      j@U�*  �V PUUU�VUUUUUUUj���*����
     �V  UT� �UUUUU�VUUUUUUU�U������     h  T �* �UUUUUU�VUUUUUUU�Z������     Z   T��*��UUUUU�UUUUUUUU���jP����*   �   P�����jUUU��UUUUUUU����Z  ��jU�  �   PP���U��UU�jUUUUUUU��j  @UU@�
  h   @P��jU���Z�jUU UUU�PU       �*  Z    @UP��jUUU���ZU UUUi         @�� �    @UQ��ZTU���UU PUUj         PU�
�    PU��V PU��ZUU UT�ZU         T��*�    PU��  UU�VU  U��jU       PU����    TU��  TUUUU  U���VU   @   TU���Z     TU��  PUUU   ����ZU  P  UY��Z    @UU��  @UUU   ����ZP  UU  UY��V     UUU�j  @UUU   ����ZQ PUU@UU�j    @UUUE�j   @UVU    �Z��ZQ TUUUUU��V    @UUUE�j   PUZU    UUU�jAUUUUUUUU��     PUUUE�j   PUjU    UUU�jAUUUUUUU���     TUUUE�j   PUiU    U T�jUUUUUUU��j     TUUUU�j   TUiU    TU�jTUUUUUU��j     TUUUU�j   TUiU   TUU�jTUUUUUUe�j      TUUU�j   TUiU   QUU��TUUUUUUe�Z      TUUU�j  UU�U   UUU��VPUUUUUUi�Z      TUUUU��  UU�U    UUUU�ZAUUUUUU��Z   @ UUUUU��  UU�U    UUUU�jEUUUUU���Z   @U@UUUUU��  UU�U  UUUUUUZ�UUUUU���Z   PUUUUUUU��  UU�UPUUUUUV��PUU�����Z  TUUUUUUU��V@UU�UTUUUUUVj�UUUU�j���ZP UUUUUUUUU�VUUU��UUUUUUUUV��VUUUUiU��ZUUUUUUUUUUUU�ZUUU��UUUUUUUZ��ZUUUjU���ZUUUUUUUUUUUUjZUUU��TUUUUU�V���V���V���ZUUUUUUUUUUUU�jUUU��TUU�UU�V�����������ZUUUUUUUUUUUU����U�jTUU�UU�Z�j���������ZUUUUUUUUUUUUi�����ZQU���UU�Z�jU��������ZUUUUiUUUUUUUi�U���Ve����UUUV��U��������ZUUU�UYUUUUUU��Z�����ZUUUU�V���V�������ZUUUiUUUUUU��j��U��V�ZUPU��V�����������ZVU�Z�ZUUUU��j��UUjUUUUUQ���������������VVUi���VUU���V��UUUUUUUUjUU���������������Z���jUU��U���VUUUUUUUUUU���������������V����V��j����ZUUUUUUUUU��������*�����V�������Z�������jUUUUUUUU��������* �����ZUU��������������UUUU    ������*  �����jU���������
   ��ZU�UU @T  �����   � �   ��������� �����* @              ���
 ��������  ��
�                    ��*  ������*      �              @U         U����               PUUUUUU         TQ                                    @UU                                    @��                                U  @�V        UTU           T     @�   U   PUUUUU               d     @d                        .UUU�W�_UUUUUUUUU5���UUUUUUUU�   WUUUUUUUU0 0\UUUUUUUU��pUUUUUUUU5� sUUUUUUUU�<�pUUUUUUUUU �UUUUUUUU�  0�UUUUUUUU�� ��UUUUUUUUU3  WUUUUUUU=  WUUUUUU���   WUUUUUU�     WUUUUUU5 �  WUUUUUU5 0��UUUUUUU� �0 �UUUUUUU� � pUUUUUUUU�0�_UUUUUUU��0��UUUUUUUs�0��WUUUUUU�5����_UUUUUU���0�_UUUUUU5����UUUUUU�0� �pUUUUUUU�0�  _UUUUUUU�  pUUUUUU�0 �� pUUUUUU5��� pUUUUUU? << \UUUUU��� �� \UUUUU� ��� WUUUUU� <?� �UUUUUUU���pUUUUUUU3 pUUUUUUU����?�UUUUUUUU�3��WUUUUUUU���?\UUUUUUU?���pUUUUUUU���UUUUUU� ?p�WUUUU�  �  0\UUUU5     �pUUUU5     p�UUUU5   0  _WUUU�������U�U.UUUU�W�_UUUUUUUUU5���UUUUUUUU�   WUUUUUUUU0 0\UUUUUUUU��pUUUUUUUU5� sUUUUUUUU�<�pUUUUUUUUU �UUUUUUUU�  0�UUUUUUUU�� ��UUUUUUUUU3  WUUUUUUU=  WUUUUUU���   WUUUUUU�     WUUUUUU5     WUUUUUU5  ��UUUUUUU� � �UUUUUUU� <  pUUUUUUUU� �_UUUUUUU��� ��UUUUUUUU�����WUUU��_U�?���_UU�  p����0�UUU����0<���UUUUU���� �pUUUUU5\3   _UU���� ���UU5    ��  �UU����33���UUUUU5\3 � �UUU���0 �� pUU�  �5����_UUU����?���UUUUUUU��� WUUUUUUU3 �_UUUUUUU����_UUUUUUU��3��sUUUUUUUU�����UUUUUUU�??WUUUUUU����� \UUUUUU= ?7? \UUUUU�    \UUUUU5  �   WUUUUU5  �  �UUUUUU5    pUUUUUU������_UU.UUUUU�W�_UUUUUUUUU5���UUUUUUUU�   WUUUUUUUU0 0\UUUUUUUU��pUUUUUUUU5� sUUUUUUUU�<�pUUUUUUUUU �UUUUUUUU�  0�UUUUUUUU�� ��UUUUUUUUU3  WUUUUUUU=  WUUUUUU���   WUUU�UU�     WUUUWU5     WUU}5\U5  ��UUU��pU� �� �UUUW�U� � pUUU5\WU��?pUUU�p5\U�U���UU�W��pUU���3WU5\WsUU���3WU�p5\sUU���3WUU��psUU���3\UUW�pUU��\UU5\pUU�?\UU��pUU0� \UUU pU� �? \UUU���U=    |UUUUU�  ���UUUUU�0  � WUUUU5�  0��\UUUU5 ���\UUUU�����WUUUUU3������UUUUUUs�� |UUUUUU��� �_UUUUUUU����UUUUUU�0�����UUUUUU�0<�?WUUUUU ��� \UUUUU ?� \UUUUU5 0  \UUUUU� �0 �WUUUUUU �  |UUUUUUU��|��WU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUWUUUUUUUUU� \_UUUUUUUU� ��UUUUUUUU5 WUUUUUUU5 WUUUUUUU5  WUUUUUUU5� �UUUUUUUU���WUUUUUUU5�  WUUUUUUU0 �UUUUUUUU0��_UUUUUUU50<pUUUUUUU� <\UUUUUUU pUUUUUUU<�_UUUUUUU���WUUUUUUU5�\UUUUUUU��\UUUUUUUU7��\UUUUUUUU�� \UUUUUUU�0�pUUUUUUU�0�\UUUUUUU5� _UUUUUUU�  pUUUUUUU  �UUUUUUU  �UUUUUUU5  �UUUUUUU5  �UUUUUUU� 3 pUUUUUUUU� pUUUUUUUU?\UUUUUUUU� \UUUUUUUU��3WUUUUUUU� �WUUUUUUU�  \UUUUUUU5  \UUUUUUU5  pUUUUUUU  pUUUUUUU pUUUUUUU� 0pUUUUUUU�?�?_UU0U�_UUUUUUUUUU=pUUUUUUUUUU�UUUUUUUUUU�UUUUUUUUUU�_UUUUUUUU�00pUUUUUUUU��UUUUUUUU �UUUUUUUU �0_UUUUUUU� pUUUUUUU �UUUUUUU�  �0WUUUUUU� < \UUUUUUU <\UUUUUUU� �\UUUUUUUU WUUUUUUUU��WUUUUUUUUU|]UUUUUUUUU�WuUUUUUUUUUUU�WUUUUUUUUUUUUU�UUUUUUUUUU� �WUUUUUUUUU��_UUUUUUUU� �_UUUUUUUUU��sUUUUUUUUU�?|UUUUUUUUU��UUUUUUUUU33�UUUUUUUUU�0�_UUUUUUUU33|uUUUUUUU� 0�UUUUUUUU�_�UUUUUUUU��W�UUUUUUUU0WuUUUUUU�U��_UUUUUUW pUUUUUUU�  pUUUUUUU�   pUUUUUUU�   \UUUUUUU�   WUUUUUUU�  �WUUUUUUUU �WUUUUUUUU WUUUUUUU�� \UUUUUUU \UUUUUUU� 0\UUUUUUU  \UUUUUUU=� WU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU]UwUUUUUUUUU���UU��UU�_� ��UU �� p�0��U�   ? �����U�  3  0�sU�3  3    �\U�� �3�3��U�� ��0��UU�? ���UU <   _�?_UU 0   w��UUU<0  �u�_U$]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]]UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUP�  �C����O����O�  OTUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUU UUU<TUU�TUU�PUU�CUUU�UUU?TUU�PUUU�CUUU�TUU�TUU�TUUU�TUUU0TUUUUUUUUUUUTUU�TUU�TUU?UUUU<UUUU<UUUU<UUUU<UUUU<UUUU<UUUU<UUUU<UUUU<UUUU<UUUU�TUU�TUU?TUU UU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �(UUUUUUUUUUU	  Q!�                       UUUUUUUUUUU	  T!*                       UUUUUUUUUUU	   ���                     �EEEEQQQQ����* ������������������������DDDDDDD  D!                        DDD����*�
    ��������������    	FDDDDjD����*
(    ��������������    ��$����*
(                �    @@@   �� ����*�
    ��������������         �   �   D!                               J�����������������������������     B  
 �D)     ���������������         B   (�R"�����(           ���
�     �   �$
"�! �� ��            �(��*         �$���D)�
   �(           �        �* $(�"(��
��            �(��
       �� (�"�!"� �(           �  �       ��"	��F)��(����            ���
�        
*��
 �"   �(           �           (����� ��
���            ��*��        � )*$ 
   (            �*   *      �
		( 
!�������              �����     � H	��@! �  �               ���    � H@
  T������                 �   � (�
  Q   �                        � 	 �  T!��*                    ��    	 )  T �          ���          *   ( 	 	  Q!*         �jUU�@            ��	 	  T!�         hUUUU
            �@J $  Q!*        �V���U�P            
@�$  T!�        `U*  jUE            (� �$  Q!*        Z�   �V)        *    $ �$  T!�       �U
    h�P       �   �� �$  Q!*       `�     �UB       B  �� ��  T!�       X)      Z	       
	 ����  Q!*       V      `%U       ($ B���
  T �       �  �
   �%       ��  
T�   Q!*      ��       ��P      �� (	(@*�
  T!�      `%   $    VR        J
� �  Q!*      `	   $    XB       	� � )  T!�      X	  �
    XI        ��   	  Q!*      X        `I       �P$   
	  T%�      V    �  `%       �    %  Q*      �        �%       � (   ($  T�      �        �%E      �* $   ��  Qa*      �     � ��%    *   �� ���  T!�     �%        �T    �  ��@ * �
  Q *     �%       �B��     �* 
 � B	  T!�     ��
      ���T    (   
	��  Q!*     �%�      $P�    �   ($ )  T!�     �e(     	��T    �    � $   Q!*     ��Z�   � HB
�    (     )�$�  T!�     �%� � *B�@�T          ��$�  Q!*     �%��� T�    �   �*����  T!�     �e`  P���*�T    � �* 	
��*  Q!*      ���!�  *��        �
(�    T!�      � ��J	`� �%E    �
 ���  @@  Q *      �� �i�	��%          � 	E  T!�      V
PUh�B)`%           
T  Q!*      XB��Z� ��eI    �
      ( P	  T!�      X� �Z $PjI           �P	  Q!*      `)PU`		�XB    �       D	  T!�      `%����IB
VR      ����������
  Q!*      ��
 �B���P                T!�       �@U ���%                Q *       Z��h �$d%     ��������  T!�       X) h�� $Z	      ��������
  Q!*       h���$�UB     !�      (  T!�       �UZ�$i�P     !�       $  Q!*        Z���V)      !�       %  T!�        `Uj� jU      !     �@	  Q!*        �V���U�P      !��������  T!�         XUUUU       !           Q!*         �jUU�@       !           T!�          ���         !����������
  Q *                       !"���������  T!�                       !           Q!*                       !           @!�                       !          �
 *                       ! ������ �� �                       !        �"*                       !       (*((�                       !�      � �� � *                       !       � ��*�                       !   ��  � ��"� *                       !�
 ( 
 � 
�(�                       !  �� � ( ��"*                       !`�"Pj� ��( �                       !�
���� X	
�**                       ! P�	X � X%�`%�                       !`�Bj`	� ����*(                      !����J� 
 ����XUUUUUUUUUUUUUUUUUUUUUU! X��
���BUe���"                      !``` *@��PT����ZUUUUUUUUUUUUUUUUUUUUUU! ����Z��UU���fUUUUUUUUUUUUUUUUUUUUUU!���@
�� U����ZUUUUUUUUUUUUUUUUUUUUUU! ��@
 UUU���fUUUUUUUUUUUUUUUUUUUUUU  "$� UU����ZUUUUUUUUUUUUUUUUUUUUUU ������ UUU���fUUUUUUUUUUUUUUUUUUUUUU         TU����ZUUUUUUUUUUUUUUUUUUUUUU         �TUU���fUUUUUUUUUUUUUUUUUUUUUU         �PU����ZUUUUUUUUUUUUUUUUUUUUUU ����������RUe���������������������������         ZU����                       TUUUUUUUU����*(RUUUUUUUUUUUUUUUUUUUUUUU        T      P                       P P P @UUUUUUUP P P P P P P T@T@T@       T@T@T@T@T@T@T@EPEPEPT P P EPEPEPEPEPEPEP@ @ @ E@T@T@@ @ @ @ @ @ @ TUUUUUUUU@PEPEPTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU @ @ TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                      UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                     UUUUUUUUUUUUUUUUUQQUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEQUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEQUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQETUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�(   @T�"                          Q!*      U�
                          T!�  ��   ��*                     ��
    *    ����
 ���������������������� ����*�      Q                           D!*  �
����
�   ��������������
   �*����*�  
(�����
   ��������������   (�����**  
(�����
   �                (�����*�  �
����
�   ��������������
   �*����**      Q                           D!�  ������������������������������������**    "Q
      *������������
      �D)�  �
����� �� �            �� �*(�R"*   ��j�� �"*            �� 
"�!�  �** (Q�� "�            �   �����D)*  
 
��� 
���"*            ��
�(�(�"�   "��h� � �            �� ��"�!*  � (�Q��*
�� *            �������F)�    � ��     �             �  ��
 �"*  
 "(�$� ����**            ����*����� �  ( ��
	�� �  �            �� ��*$ *  �*
�B�������*              ����( 
!�    �*P    �                �� ��@!*  ��  U��*��*                 ��
  T!�  �� @  *                    ��
  Q *      U����                        T!�      �"          ��P            T �     @T�
         �UU�           Q!*      U�"        �UUUU)P           T!�     @T�
        ZU��V�B          Q!*      U�"       �U� (�U	         T!�     @T�
       h� � Z�P          Q!*      U�"       V)  � �UB         T!�     @T�
      �U  (  V	         Q!*      U�"      `�      h%         T!�     @T�
      X	      ��T        Q!*      �"      X       �P         T �     @T�
      V       VB        Q!*      U�"     ��        XI        T!�     @T�
     �%        `	        Q!*      U�"     `% �     `%        T!�     @T�
     `	      �%        Q!*      U�"     X	 	 �
  ��T        T!�     @T�
     X 	      �        Q!*      U�"     X �  $  ��       T!�     @T�
     X       �
�P        Q!*      U�"     �     �
  PXR       T!�     @�
     �        
�ZR        Q *      U�"     �*       B
XR       T!�     @T�
     ��
     ��@YR        Q!*      U�"     ��      $�ZR       T!�     @T�
     �j  � 	)XR        Q!*      U�"     �� ��IYR       T!�     @T�
     �h  
P J�PYR        Q!*      U�"     �i���@�`��XR       T!�     @T�
     X����h�� VR        Q!*      U�"     X���PV��T�       T!�     @�
     X�
 �P�&P��        Q *      U�"     X)@U�P���T        T!�     @T�
     `	���P`B
�%        Q!*      U�"     `I
  PY��@e%        T!�     @T�
     ��@U%P�%$�j	        Q!*      U�"     ����*@&	)XI        T!�     @T�
      V*  @YIVB        Q!*      U�"      XU)@iHBR�P         T!�     @�
      h��
 eH���T         Q!*      U�"      `�  d��h%         T!�     @T�
      ��V@e�V	         Q *      U�"       Vi)@i��UB         T!�     @T�
       h�fUYZ�P          Q!*      U�"      ���������          T!�     @T�
      
    ����
          Q!*      U�"     �����������          T!�     @T�
     �����������          Q!*      U�"     ��������
�         T!�     @�
     �(
hUUU���         Q *      U�"     �*�ZUUUU*��         T!�     @T�
     �
�    �
�          Q!*      P�"     �
j     �
*          @!�     ��
      �*     �*          �
 *    � (�"      �     @*         �� �    ���
      �     @*          �"*    
�

�"      �     @*         (*((�    �" (�
      �     @*         �� � *    *���"      �     @*         ��*�    *��*�
      �     @*         ��"� *    ��� �"      ��������*         
�(�    
(��
      ���UUU���         ( ��"*    � 
�"      �j�fff��*         ��( �    V����
      � ���
@*         X	
�**    V� X�"      �      )         X%�`%�    ����
�      �      )         ����*( U� ��*(VUUUUU�FUUUUUiUUUUUUUUU
 ����  �PU����     �      )        �BUe���" U%Ue���VUUUUU�FUUUUUiUUUUUUUU�PT����
 U)EU����YUUUUU�FUUUUUiUUUUUUUU�UU���" U	EUe���VUUUUU�FUUUUU�UUUUUUUU%U����
 UIEU����YUUUUU�FUUUUU�UUUUUUUU%UU���" UIUUe���VUUUUU�FUUUUU�UUUUUUUU%UU����
 UIUU����YUUUUU�EUUUUUU�UUUUUUUU%UUU���" U	UUe���VUUUUU�AUUUUUU�UUUUUUUU%TU����
 U)UU����YUUUUU�QUUUUUU�UUUUUUUU�TUU���" U%TUe���VUUUUU�QUUUUUU�UUUUUUUU�PU����
 ��TU����������������������������RUe���"  �VU��*(     �      �         ZU���� U����
�PUUUUU�QUUUUUU�UUUUUUUU����*(             �      �        P     X  PPUUUUUU@ P �Q P P�P P P@UUUUUY  T        P@T@�T@T@T�T@T@T      X  E@P P TPEP�EPEPE�EPEPE@P PX  @PT@T@E @ �@ @ @�@ @ @PT@TX  U EPEP@UUUU�UUUUUUU�VUUUUUUU EPEX  UU@ @ TUUUUU�UUUUUUU�VUUUUUUUU@ @X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX                                UUUUUUPX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUX                               PUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUUQQUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUTQUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUEQUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUQQUUUUUPX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUQQUUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUU QUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUETQUUUUU X  UUUUUUUUUUUUUUUUUUUUUUUUUUUTQUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUUUUUX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUUUUUPX  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUUUUUUX  ,UUUUUUUUUUUU���UUUUUUUUUUUUUUUUU  �_UUUUUUUUUUUUUUUU � pUUUUUUUUUUUU��U5 �?�UUUUUUUUUUU����W�  �WUUUUUUUUUU�����U �\UUUUUUUUU��� �_=  �sUUUUUUUUU��0  ��� �UUUUUUUUU�? � �W= ��UUUUUUUU���������WUUUUUUU�������UU=�_UUUUUUU��0�����_U��_UUUUU�_����W��?��UU�UUUUU������U����UU�UUUUU�����UU��?�_U=�UUUUU�����sUU����U��UUUU�������UUU���_�UUUU�����?��WU��? ��UU�_�������_UU�� ���UU5��_���?���WU�����UU��W���� ��_U��? ��UU��U��� ��_U������_��U��?   _UU������sU��UU�   �}UU�������U��WU�   ��UU����������_U�?   ��UUU�����p5\U=��  � _UUU�W��U�\\U   0pUUUUU�WUWW�     ��UUUUU�\UU�UU    UUUUUs5\UUUUU�    0�WUUUU��_UUUUU   ���UUUWUUUUUU50     �WUU�UUUUUUU��   �  <WUUUUUUUUUUU  �  ? �WUUUUUUUUUUU  0  ��UUUUUUUUUUUU5  �  �UUUUUUUUUUUU�   < � pUUUUUUUUUUUUU  ��WpUUUUUUUUUUUUU  �UU=\UUUUUUUUUUUUU�  pUU=WUUUUUUUUUUUUUU _UU�UUUUUUUUUUUUUUU=�UUUUUUUUUUUUUUUUUUU�UUUUUUUUUUU5UUUUUUUUUUUU��UUUUUUUUUUUUUUUUU�  UUUUUUUUUUUUUUUU  �WUUUUUUUUUUU��_��? \UUUUUUUUUUU���_ �?pUUUUUUUUUU�����  ��UUUUUUUUUU�?��U ��UUUUUUUUU��0�= ��WUUUUUUUU��� �� �_UUUUUUUU�� ����W=��UUUUUUUU�?��� �_��UUUUUUUU�������UU�UUUUUUUU�������_U5�WUUUUUUU��_��? |U5�WUUUUUU���W��� �W��_UUUUU���?<WU����_��_UUUUU���?_U��? ���_UUUUU���� _U��� �?�_UUUUU���� _UU���0�_UUUUU����UU��? WUUUUU������UUU����UUUUUU����?�WUU��?��W�UUUU����?�_U}U�����?WUUU������U�U�����?\UUU�_����U�}������\UU��W����_��U��U�W_�_�UU��?���WUU��_U5��_UU���  ��_UU��pU��WUU��  ��_UU���U��UUU��  ��UU5W�U��UUUU�   �UU5\�UU��UUU�0<  �WU�pUUU��WUU5 �  � WUU_UU���_UU    ��\UUUUU�p5\UU5    0��WU�UUU�\\UU�    0 ���UUUUWWUUU�   � � ?<WUUUU�UUUU    �  WUUUUUUUUU50      �UUUUUUUUUU��  � �? UUUUUUUUUUU  0 ��pUUUUUUUUUUU   �U�pUUUUUUUUUUU5   �W�\UUUUUUUUUUU�  0 �_�WUUUUUUUUUUUU �� UUUUUUUUUUUUUU=  p|UUUUUUUUUUUUUU��_��uUUUUUUUUUUUUUU�UU��UUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUU=|UUUUUUUUUUUUUUUUUU�WUUUU7UUUUUUUUUUU�WUUUUUUUUUUUUUUU� �UUUUUUUUUUUUUUU  WUUUUUUUUUU��U� \UUUUUUUUU����W5 �pUUUUUUUUU����_� ��UUUUUUUUU�?��U WUUUUUUU����_= �WUUUUUUU��  ��_UUUUUUU�� ����W��_UUUUUUU������U5UUUUUUU�?���? �U5UUUUUU����_����_�UUUUUU����_��?��UUUUU��?�WU�� ��_UUUUU���?<WU��3��UUUUU���?_UU�?���W�UUU���� _UU�����_?WUU���� _UU������?\UU����UUU���U��\UU������UUU��WU�W_UU�����WUUUUUU�_UUU�_��?�_U�UUU��pUUU�W��?�_U�WUU���UUU�U��� U��UU5W�UU�U����W��WU5\�UU�U�������_U�pUUU�UU��?  ��UU_UUU�_UU��   UUUUUU�_UU��    ��UUUUU��_U��   ��WU�WU���U�   ��W��WU����U �   0 _=�\U����U     �?\ \U���U     ��  WU�\�U5     < �UU�5\sU�?    ���UUu5\]UU�    �WsUUU5WUUU    pU_UUU�UUUU50  � ?\UUUUUUUUUU�   0 �_UUUUUUUUUUU   �UUUUUUUUUUUU   �UUUUUUUUUUUU5  0 �UUUUUUUUUUUU�  �?�WUUUUUUUUUUUU  ��WUUUUUUUUUUUU��__UUUUUUUUUUUUU�U|}UUUUUUUUUUUUUUU5�sUUUUUUUUUUUUUUU�0pUUUUUUUUUUUUUUUU�\UUUUUUUUUUUUUUUU_UUUUUUUUUUUUUUUU\UUUUUUUUUUUUUUU��WUUUUUUUUUUUUUUUUUUUU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUU�  �UUUUUUUUUUUUUU ? pUUUUUUUUUUUUUU� \UUUUUUUUUUUUU��?  WWUUUUUUUUUUUU5� �UUUUUUUUUUUUUU��  |UWUUUUUUUUUUUU� �WU\UUUUUUUUUUUU�? |UUpU_UUUUUUUUU����WUU��sUUUUUUUUU�?|UUUU�?�WUUUUUUU��WUUUU�|UUUUUUU���UUUUU��?�UUUUUU���sUUUUU����WUUUU?��_UUUUU���? ��U�����WUUUUU����� ����UUUUUU������? ����_UUUUUU������������UUUUUUU ����������WUUUUUUU ��������WUUUUUUUU= �������_UUUUUUUUU�������_UUUUUUUUUU����?��_UUUUUUUUUUU��_��}UUUUUUUUUUUU�U����UUUUUUUUUUUU�WUU��WUUUUUUUUUUU�UUU��?WUUUUUUUUUUUUUU���WUUUUUUUUUUU�UUU��WUUUUUUUUUUUU�UUU�?\UUUUUUUUUUUU�WUU�7pUUUUUUUUUUUU�WUU��pUUUUUUUUUUUUWUUWUUUUUUUUUUUU�UUU5\UUUUUUUUUUUUUUUU�WUUUUUUUUUUUUU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUU�  �UUUUUUUUUUUUUU ? pUUUUUUUUUUUUUU� \UUUUUUUUUUUUU��?  WUUUUUUUUUUUUU5� �UUUUUUUUUUUUUU��  |UUUUUUUUUUUUUU� �WUUUUUUUUUUUUUU�? |UUUUUUUUUUUUUU����WUUUUUUUUUUUUUU�?|UUUU_UUUUUUUUUU��WUUUUUUUUUUUUUUU���UUUUUWUUUUUUUUUU��sUUUUU\U�UUUUUUU���_UUUUUpU�WUUUUUU=��WUUUUU��|UUUUU���UUUUUU�?��UUUU����_UUUUUU���UUU���UUUUUUU���? ������_UUUUUUU����� ����UUUUUUUU������? ��_UUUUUUUU����������UUUUUUUUU���������_UUUUUUUUU��������UUUUUUUUUU �������WUUUUUUUUUU  ������UUUUUUUUUUU? �����_UUUUUUUUUUU�����UUUUUUUUUUUU�����UUUUUUUUUUUUU��U�?�_UUUUUUUUUUUU�_U���sUUUUUUUUUUUU�WUU���UUUUUUUUUUUU�UUU���UUUUUUUUUUUUUUU��UUUUUUUUUUUU�UUU��UUUUUUUUUUUUU�WUU�WUUUUUUUUUUUU�_UU�\UUUUUUUUUUUU5\UUs5\UUUUUUUUUUUU\UU��_UUUUUUUUUUUUWUUWUUUUUUUUUUUUU�UUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU              �(Uj����V�V�i��jUj�RUUUUUUUUPUUUUUUUUUUU�����Z��ZiZ�U��ZU��  TUUUUUPUUUUUUUUUUUj��e�V�UiUZi�U�Z��PUUPUUUUU @UUUUUUUUUU�UeU�Rj���ZieU�V��
TUU TUUUU  UUUUUUUU�UYV�BZi��iYe��U��BUUUUUPUUUUUEPUUUUUUU�V�ZU
ZYe����j��( PUUUUUAUUUUUTTUUUUUUUVfi�*i�Z���UUj�*UUUUUU UUUUUTUTUUUUUU@VYe�*dU�*�Vj�V�
UUUUUUUUPUUUUPUPUUUUUUHZ�Z���Zj �Z�V%�@UUUUUUUUUAUUUUAUAUUUUUUJ�V�B��Z�Z�*TUUUUUUUUUEUUUUTEUUUUUU
@���
U�Z�Ui�UUUUUUUUUUUUUUUPEUUUUUU(
 P *(`UeU���PUUUUUUUUUU TUUUQEUUUUUU�*��
��jJYeU�
TUUUU PUUUUTUUUQUUUUUUU ���*@��RIY�U�@UUUUU�BUUUU TUUQUUUUUUU��
U�P	e�U�PUUU  �
  TUUTUUQUUUUUUU �BUU�R)�j��BUUU�*����PUUPUUQUUUUUUUUU PUU�JTeJUU�
�*�RUUQUUUUUUUUUUUUTUUU*P���JUU�J!@U� RUUAUUUUUUUUUUUUTUUU�U��@UU�@ UU�TUU UUUUUUUUUUUTUUUU*  �*TUU�X�UU�V�UUEUTUUUUUUUUUUUUUUU���� UUU�X�UU V�TUEUUUUUUUUUUUUUUUT�
�*TUUU�X�ZU jRTUEUTUUUUUUUUUUUUUEU@
UUUU�XhU�RTUEUUPUUUUUUUUUUUUUAUUU@UUUU!X`UA�
RTUEUU@UUUUUUUUTUUUQUUUUUUUUU ZUhUQ�
RTUEUUUEUUUUUUUUUTUUUQUUUUUUUUU(VUhUQ�RTUUUUEUUUUUUUUU@UUUQUUUUUUUU(VU�UQ�RTUUUUUUUUUUUUUDUUUQUUUUUUUU�VU�UQ��RTUUUU TUUUUUUUUUU@UUUUUUU�UUhUU��BUUUUUUPUUUUUUUUUUEUUUUUUU��UUhUU��
UUTUUUQUUUUUUUTUUEUUUUUUU�jUUhUU��*TUUPUUUAUUUUUUUTTUUEUUUUUUU�ZUU�UU���TUUQUUUEUUUUUUUTTUUEPUUUUUU�ZUU�UU�PUUPUUPEUUUUUUTTUUEUAUUUUU�ZUU�UU�RUU@UUUQUUUUUUUUTUUEUEUUUUU�YUU�UU�VRUUUUUQUUUUUUUUTUUUEUUUUU�YUU�UU�jBUTUUQUUUUUUUTPUUTUUZiUU��YUU�VU`JUUPUUQUUUUUUUUTAUUUTUU�ZUU�UUV�VjUZa(UEUQUUQUUUUUUUUTEUUUPUU�UUU�UU�jU����`(UEUAUUQUUUUUUUUTUUUUQUUUUUhU��UeU����a UEUEUUUUUUUUUUPUUUUUUUUUZ��VU�UU�*�a!UEUEUUUUUUUUUUQUUUUTUUUU!V%ZU�VZU�"�a!UEUEUUEUUUUUUUQUUUUETUUZY�V�UUiU�UU��!UEUUUEUUUUUUUEAUUUUQTUU�Z�U�VUUQVUj��!UQUUUEUUUUUUPEUUUUPTUU��U�U�j��iUi��%UQUUUEUUUUUUAUEUUUUTTUUUjU�Uej��fUi��&UQUUUUUUUUUUQUEUUUTPUUUjU�VYVeU�Uj��&UQUUUUUUUUUUQUEUUUUQU �ZU�UVUUUUV�U�
UQUUUUUUUUUUUTUEUUUEUQU*�ZU�UZUQ�V�U�
UQUUUUUUUUUUUTUEUUUAUQU��VU��ij���Y�UU
UQUUUUUUUUUUTUEUUUQUAU���VUi��i��iZ�UU�TUUUUUUUUUUUUTUTUUQUEU� �VUj�QeQY�VU�TQUUUUUUUUUUUTUEPUUPUEU!D"VUj�UUUUUY�VU�PQUUUUUUUUUUTUEQUUTUEU E�UUb�UUUUUY%VU�RQUUUUUUUUUUUUEAUUTUE(U�VUY�QUeUY�UU�RUUUUUUUUUUUUUEEUUTUE
UYZU���i��iZ�U��RUUUUUUUUUUUUUEUUUTUE�B�U�U�Vfj��fVjU��PEUUUUUUUUUUUUEUUUPU�@�ViU�ZZUQ��ZU��TUUUUUUUUUUUUUEUUUQU�D�ViUejYUUU��fU��TUUZiUUUUUUUEUUEUUUAU�T�V�UU�ie�e��UUi�PUU�ZUUUUUUUEUUEUUUEU�T�V�YU��i��ijV�i�RUU�UUUUUUUUQUUEUUUEU�T�V�VU�ZEQ�ZUU�URUUUUUUUUUUUQUU@UUUEUU T�V�ZUUjjU��VU�ZURUUUUUUUUUUUUUUDUUUAUU T�ZU��Z���Zi��*VURi�UUUUUUUUUUUUTUUQUU U�ZU���ViU�U���UUR�jUUUUUUUUUEUUTTUUQUU(U�ZUUU�Z��i��VUUURUVUUUUUUUUUUUTTUUQU(U�ZUUUU�UFVYUUUUURUUUUUUUUUUUUUUTUUUU*U�ZUUUU�VUUZUUUUURUUUUUUUUUUUUUUTUUUU&U�ZU����QTY���VURUUUUUUUUUUUUUEUUUUUU&U�Ze������i���*fUBUUUUUUUUUUUUUEUUUUUU&U�Z�ZUUUjU�VUU�ZUJUU PUUUUUUUUEUUUUUUV��Z�ZUUi��Z�UU�ZUJZi��BUUUUUUUUEUUUUUUV��Z�VU�jiU���UUZ�J�Z� JUUUUUUUUEUUUUUUV��Z�V��VVUUV�ZUjUI�U!HUUUUUUUUEUUUUUU�V��Z�U&V�jU�ZUbViVIUUaTHUUUUUUUUEUUUUUU�T��Z�U�Ue�V
fU�U�UIUUaTUUUUUUUUE@UUUUU�T��ZiUiUe� fU�U�UJUU`�*UUUUUUUU@UUUUUaT��VbejUe	V�eU�f%VIUUh� UUUUUUUUUUUUU`TY�VZ�ZUe�U�eU�Z�VJUX� UUUUUUUUAUUUUUhTY��Z�fUeU�UeUeZ�Z*UZ� TUUUUUUUAUUUUhP���Z�UU�iU�iUUY�V*UZ��TUUUUUUUPTUUjP��Vi%VU�Z��ZUUb�U&U�j��TUUUUUUPTUU�VQ��Vi��UUYV�UU�j�U&UhZ��PUUUUUUTDPUU�PU��Uf���Ui��U��ZeV&UXZU�RUUUUUUT@@UU�TU��U�U��j��j��jUi�&�jU�PUUUUUPT P U�T��jY�UUUUUUUUUUUY�&�jU�RUUUUUP      �U��VZ�VUUUUUUUUUUZ���jUUUUUU@ @ T�U���VUVUUUUUUUUUUV���jU*PUUUU @UUUUU�U��fUUVUUUUUUUUUUV�U�jU�RUUUU  UUUUU�U��f�UU�UUUUUUUU�U�U
��URUUUUUUUUUUU�U��feUU�UU���V�U�U�U	��URUUUUUUUUUUU�U��feUU�UU���Z�UeU�U��URUUUUUUUUUUUVU��eUUU���Z����UaU�U(��URUUUUUUUUUUUV���iUUU�������jU`U�U���ERUUUUUUUUUUU�V��ZiUUU��Y����jUaU�U���URUUUUUUUUUUU�U���ZUUUU�������U`U�V����URUUUUUUUUU�U�V���YUUUU�����j�VeU�Va���URUUUUUUUUU�U`V���YUUUU���j���VUU�Ua���UUUUUUUUUU�VhV���YUUUUf��j���VVU�U����U*PUUUUUUUY�VXU�jYYUUUUf������ZVU�U����U�RUUUUUUUj�ZXU�jZUUUUUe����j�ZVU�Ua���URUUUUUU�j�ZXU��YUUUUUi��Z�Z��VU�Ua���ZUJBU�UUUU���*X���iUUUU�Z��jV��jUU�Ve��XUYBU�UUUU����Z���eUUUUU���jU��jUUUVeY�XUYB��UUU�����Z���eUVUU����jU��jUUVei�XUYJ��Z����UU�V�V�eUVUU�����Y���UUVee�XUY	��ZUUUUU��UU�jeUVUUU��������UUVUe�*VUU���jUUU����*aeUVUUU��������jUVUe�(VUY���� U  
    `�UVUUe��������UUUVU��(UUUY���i�UVUUe��������jUUVU�V�UUUY���          XUUVUUe��������eUUVU�U�UUY����ZUZUUe��������UUVU�T�VUU	             jU�UUe��������UU�VU�T��TUIUU�U�UUe��������UU�UU�Q�����JUU           ���UUe�"
  ���iU�UU�UaU��*@UU�ZU�  �ZU�UU�UiUUUUUU              ��*        �jUU���ZUUUUUUU   �jU�UUUUUUUUUU                          ����UUUUUUUUUU    QUUUUUUUUUUUU                           UQUUUUUUUUU      PUUUUUUUU                            UUUUUUUU       PUUUUUUU                            QUUUUUU         TUUUUU                            QUUUUU        UUUUU                              UUUU          QUUU                                UU           QU                                @U                             Q    @                            @                      @                                                                                                           @                                                                                                                                      @       �(Q)YU  �U�Ue��Z���B T �VP�@����U*YU�  � �Ve
j�Z�� BBe �Z ��P����e*YU� �jd�Re���V�� @VjEA�ZP��������*YU� hj��Re���V�� P�jU������������iYU� hjj�Re`�jZ�� @V�Z����U������hiYU��hjEZ�Reh�Zj�� Pf��VY���������Z�UU��jjEZ�Re!h�ZjZ�
 T�U����V�������Z�UU��j�UV�Re Y�V�V�F�d��U���Vi�V���*�V�UU`�j�V�bU`Z�V�V�V� ��jU�ZVUi����Z�U�UU`�j�V�bU`V�Z�V�V� ��jUUjZUi����V�U�UU`���%V�*�V�Z�V�V��d�ZUUjVUe�Zf�V�U�TU ����V�&`U�Z�V�Z��d�ZUUjVUUUZj�V`U�TU h���U�*`U�Z�V�Z�f�ZUU�VUUUZV�V`U�TU*X��fU�*hU�Z�VUZ� j�VUU�VUUUj	��V`U�PUX��jU�*iU�ZUUUi�VUVUU�UUUUjI��Z`U�XUXi�fUU*YU�VUUU��VUUUU�UUUUjiV�Z`U�XU
Xe�jUU
ViU�UUUU�VUUUU�UUUUj�V�ZhU��U�YUUUUUi�ZUUUUUU�ZXVUUUUUUUUU�jUU�&ZU��U�YUUUUU��YUUUUUU�j�VUUUUUUUUU�ZUU�&ZUU�T�ZUUUUU��UUUUUUU�j�VUUUUUUUUU�VUU�&VUU�T�VUUUUUUjUUUUUUU�j�VUUUUUUUUUUUUU�*VUU�T�UUUUUUUjUUUUUUU�j�VUUUUUUUUUUUUU��VUU�U�UUUUUUUiUUUUUUU�j�UUUUUUUUUUUUUU�fUUU�U�UUUUUUUYUUUUUUU�j�UUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUUj�UUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUUUUUUU�jUUU�T�UUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUZUUU�TYUUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUUUUU�TZUUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUUUUU�XVUUUUUUUUUUUUUUUUUZUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��FUUUTUUUTUUUTUUUTUUUTUUUTUUUTUUUTUUUQTU�VTUTUTUTUTUTUTUTUTUTUTUTUTUTUTUTUTUTEEEjEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEETTTjTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                                        QQQQQQQQQQQQDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �������������                          UUUUUUUUUUUU���                        UUUUUUUUUUUUUUU�                       UUUUUUUUUUUUUUUU*                                  @UUUU�                    PQ              UUU
                    ��               @U)                    &                T�                   �*                @U
                   �                 T)                 ����                 P�            ����VU�j                 PU�          ��jUUUUU!`                  T�
        �ZUUUUUUU �                   U�       �VUUUUUUUU UUUUUUUUUUUUT     @�
      jUUUUUUU  ��UUUUUUUUUUUUUU     U)     �VUUU     �*UUUUUUUUUUUUUU     T%     �UUUU     �*UUUUUUUUUUUUUEU     P�   �VUUU     @(UUUUUUUUUUUUUUU    @U
   �UUU       ���UUUUUUUUUUUUUUUU    @U�  �jUU       T� �UUUUUUUUUUUUUUUU    U� �UU       ��*�UUUUUUUUUUUUUUUUU    UU�ZUU       ���UUUUUUUUUUUUUUUTU    PU
�UU        �*  UUUUUUUUUUUUUUUUU   @U)TUU        �	UUUUUUUUUUUUUUUUU    U�TU         �	**UUUUUUUUUUUUUUUUU    U�PU         �	**UUUUUUUUUUUUUUUUUU    T�B          �)UUUUUUUUUUUUUUUUEU   TUJ          �)� UUUUUUUUUUUUUUUUUU   PU	          ����UUUUUUUUUUUUUUUUUU   PU)         Tb�V�UUUUUUUUUUUUUUUUUQU   @U%       TUbU�jUUUUUUUUUUUUUUUUQUU  @U�     @UUU��U"bUUUUUUUUUUUUUUUUUUQ   U�     UUUU��U�jUUUUUUUUUUUUUUUUUUU   U�R    TUUUU��UUUUUUUUUUUUUUUUUUUUUU   TUB   @UUUUU�XVUUUUUUUUUUUUUUUUUUUEUU   TUJ   TUUUUU�iVUUUUUUUUUUUUUUUUUUUUP   PUI @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUQ   PU	 PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUP   @U)@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  @U%UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   U%TUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUU   U�TEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   T�T@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQ   T�TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P�TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P�TUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUTUU   P�PUUUUETUUUUUUUUUUUUUUUUUUUUUUUUUUUU  P�RUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUQU  PURUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  @URUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQ  @UBUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   UJUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@UU   U	UUUUUUUUUUUUPUUUUUU@UPUUUUUUDUU   U)UUUUUUUUUUUUUQUUUUUUDUQUUUUUU@UU   U%TUUUUUUUUUUUUPUUUUUU@UPUUUUUUUQU   U�TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   T�PUUUUUUUUUUUUUUUUUUUTUUUUUUUPU�*� PUBUUUUUDUUUUUUUUUUUUUETUUUUUUUQU���PUJUUUUU@UUUUUUUUUUUUUTUUUUUUUPU)  
PU�jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU	PU	����ZU�Z����UUUUUUUUUUUUUUUUUUUUE	**Pe�      �*   UUUUUUUUUUUUUUUUUUUUU	**PU
*������ �
�UUUUUUUUUUUUUUUUUUUUU)
PY	*   (��������
������*��
������j*�*� ��(*�����������*                  � ���   ���������
������������������� ����������������������������������������*�������
   ������������������*��  ������"����* ���������������������*�����
 ����������������������6UUUUUUUUUUUUUUUUUUUU}UUUUUUUUUUU�UUUUUUUUUUU�_UUUUUUUUUUpUUUUUUUUUU0�WUUUUUUUUU5� \UUUUUUUUU� �UUUUUUUUU�  WUUUUUUUUU�0\UUUUUUUUU=�pUUUUUUUUU0 sUUUUUUUU� 0 pUUUUUUU�� � \UUUUUU}�� sUUUUUU�\ �pUUUUU_��  pUUUU�p5   pUUUUU��0 0  pUUUUUW�    pUUUUU5\   pUUUU��p5   \UUUUW���  \UUUU5\���  WUUUU�p5�<��UUUUUU��0�  �WUUUUUW\ �_UUUUU5� \��UUUUU�  \����UUUUUU�������UUUUUUUU�����WUUUUUUU?�WUUUUUU�0 � WUUUUUU5��  �UUUUUUU0 �UUUUUUU� �UUUUUU� � pUUUUUU=�0 pUUUUUU�� \UUUUUU0<0_UUUUUU���?�UUUUUUUp?���WUUUUUU�_� �WUUUUUUUU?��_UUUUUUU����?\UUUUUUU�?3��|UUUUUUU5���?�UUUUUUU5<�=� WUUUUUU���? \UUUUU�  �  \UUUUU  0   \UUUUU  0   WUUUUU  �  �UUUUUU�����WUU6UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��WUUUUUUUUU��\UUUUUUUUUU�UUUUUUUUUU0 WUUUUUUUUU5� |UUUUUUUUU5� �UUUUUU_UU�� WUUUU�pUUU0\UUU�W�UU� �\UUU5\WU5  \UUU�p5\}5 0 WUUUU��p�5��\UUUUW� �3 <\UUU}5\<3  \UUU��p5 <  \UUUW�5    \UUU5\7    \UUU�p5    \UUUU�� �   WUUUU? ��   WUUUU5  W�? �UUUUU��?\�pUUUUUUU��?  �UUUUUUUU� ��WUUUUUUU���_UUUUUUU3����UUUUUUU��?��UUUUUUU5�33��UUUUUUU�0����UUUUUUU5? <�UUUUUUU�0 �UUUUUUU �  pUUUUUU�  3 pUUUUUU5 0 \UUUUUU� �0 \UUUUU� 0� WUUUUU� ��WUUUUU� ���?UUUUUUU����UUUUUUU��0 �UUUUUUUU����WUUUUUUU�?���WUUUUUUU���?\UUUUUUU�����sUUUUUUU|0�UUUUUU��s� WUUUUU=  �   WUUUUU     WUUUUU    �UUUUUU  0  UUUUUU������UUU;UU_UUUUUUUUUUUU�pUUUUUUUUUUU�W�UUUUUUUUUUU5\WUUUUUUUUUU�p5\UUUUUUUUUUU��pUUUUU�UUUUUW�UUUU�_UUU}5\WUUUpUUU��p5WUUU0�WUUW�5WUUU5� \UU5\7WUUU� �UU�p5WUUU�  WUU�� WUUUU�0\UU? WUUUU=�pUU5  WUUUU0 sUU��?\UUU� 0 pUUUU��UU�� � \UUUUUWU�< sUUUUU\U\� �pUUUUU3p� ��  pUUUUU���  �  pUUUUU5��     pUUUUU�0|    pUUUUUU�    pUUUUUU �   \UUUUUU5 ��  \UUUUUU� ���  WUUUUUUU <��UUUUUUUU �  �WUUUUUUU5 ���\UUUUUUU�  �?sUUUUUUUU ��?sUUUUUUUU ��?sUUUUUUUU5 ��?�UUUUUUUU5 0���UUUUUUUU� ��3�UUUUUUUUU �UUUUUUUUU � WUUUUUUUU5    WUUUUUUUU�    WUUUUUUUUU?   WUUUUUUUU�� �\UUUUUUUU�?�?pUUUUUUUUU�� ��UUUUUUUUU����UUUUUUUUU���?�UUUUUUUUU���?pUUUUUUUU�����_UUUUUUUU�?��UUUUUUUU_����UUUUUUU��3����WUUUUUU5 ����\UUUUUU5  �?�sUUUUUU5  <���UUUUUU5  ��? �UUUUUU�   �  �UUUUUUU  0  |UUUUUUU�   �WUUUUUUUU����U8UUUUUUUUUUUUUUUUU}UUU_UUUUU�UU_UUU}U�UUU�U�WU]U�U�UUU�U�UU{U�_�WUUuUU��WUUWUU}�_U��~U�U_Uu_�WՊ��U�W}W�_�U����_�\�U�W}U����^U_�U�WU몮�zU�W��ժ����U��W�Uի����U�_�U_������W}�\u�_������W�UW��_������W��W��_������W��W��\������W��W�UW������Wu�W�U������W�W�W��������_�W�W�׫�����W�]�W�_����z�]�U�WU����~U�U�W�������U�U�WU�ת���WU�U�WU������UU�U���W=��_���UU�����>���UUu��þ����UWUUUUU���SUUUUUUU����WUUUUU���(*���UUUUU���S�_UUU��U����\��UUU5_U?��U=WUU�U�_���U�_UU�U�ת���W�_UU�U������_�_UU�Uu����^W�UU}U������\U_UU}U������_U_UU}U������U_UU}U������_U_UU]U������_U]UUsU}����W_UsUUU}U��zU_UUU}U}U��~U_U_UU�UuU��_UW�_UU�W�UUUU�\�wUU�W�UUUU�_�UUUU_�_UUU�W}UUUU}��UU��U_UUUU�U�_U�W�WUUUU�UU}U_U�UUUUUUUUUUUUUUUU4UU�U���U�UUUUU�U}�W_�WUUUU}�W�~�U_UUUU_�����_}UUU�����^��UUU�5�����5�WUU���������_UU���ꪮ�_U�_}�����^_�U5W�����_5W�U_�����{}�U��_�����~��W��W��芪x��W��W�����z��W��U�����z��W�uU��ꪪxU�W��W�����~��W��_�����^��_�U�����_�_�����������W�U�������W�W�U���<���]�_�UU���_U�_}UU�����_UU_���  �U��\���������WUU�?����_UUUUU�.�:UUUUUUU?���>UUUUU�?���8�_UUU�����>��UUU�_�����U�_UU�U�  �W�sU�_U�����_U�UU_U���^U}UU�_���z�UUU}Uת���uU_UU���������_UU��߮�����WUU��ߪ�����WUU�Wߪ���}�WUU�U�����}�UUU5W_���}5WUU�W_���W}�WUU�W_���W}�UUU�_����s�UUUU�UU�_UUUU}U�W�U_UUUU�UU�_U�WUUUU�WUUUU�UUUUUU_UUUU}UUUUUU]UUUU]UUUUUUuUUU�UUW�U�\�U����5�5��5�
��������_                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      U���W�U���_�U����U��p�U�  �U���������?�����?w����?w����?w�����wU����uU���uU5��\uU�  _]U���]U���]�����W�����_����?p3�0p����\���_���u� p5 WUp��UUpUUUU�_UUUxUU�UUUUUU����������UUUUUUUUUUU�UUUUUU����������UUUUUUUUUUU�UUUUUU����������UUUUUUUUUUU�UUUUUU����������UUUUUUUUUUU�UUUUU��   ��   ��UUUUUUUUUU�UUUUU��   ��   ��UUUUUUUUUU�UUUUU��   ��   ��UUUUUUUUUU�UUUUU��   ��   ��UUUUUUUUUU�UUUU����� �� �����UUUUUUUUU�UUUU����� �� �����UUUUUUUUU�UUUU����� �� �����UUUUUUUUU�UUUU����� �� �����UUUUUUUUU�UUUU�     ��     �UUUUUUUUU�UUUU�     ��     �UUUUUUUUU�UUUU�     ��     �UUUUUUUUU�UUUU�     ��     �UUUUUUUUU�UUUU��������������UUUUUUUUU�UUUU��������������UUUUUUUUU�UUUU��������������UUUUUUUUU�UUUU��������������UUUUUUUUU�UUU���    ��    ���UUUUUUUU�UUU���    ��    ���UUUUUUUU�UUU���    ��    ���UUUUUUUU�UUU���    ��    ���UUUUUUUU�UU� �            � �UUUUUUU�UU� �            � �UUUUUUU�UU� �            � �UUUUUUU�UU� �            � �UUUUUUUU�U�    ��    ��    �UUUUUUUU�U�    ��    ��    �UUUUUUUU�U�    ��    ��    �UUUUUUUU�U�    ��    ��    �UUUUUUUU�U� �            � �UUUUUUUU�U� �            � �UUUUUUUU�U� �            � �UUUUUUUU�U� �            � �UUUUUUUU�U� �     ��     � �UUUUUUUU�U� �     ��     � �UUUUUUUU�U� �     ��     � �UUUUUUUU�U� �     ��     � �UUUUUUUU�U���  �      �  ���UUUUUUUU�U���  �      �  ���UUUUUUUU�U���  �      �  ���UUUUUUUU�U���  �      �  ���UUUUUUUU�UU��   �    �   ��UUUUUUUUU�UU��   �    �   ��UUUUUUUUU�UU��   �    �   ��UUUUUUUUU�UU��   �    �   ��UUUUUUUUU�UUU��   ����   ��UUUUUUUUUU�UUU��   ����   ��UUUUUUUUUU�UUU��   ����   ��UUUUUUUUUU�UUU��   ����   ��UUUUUUUUUU�UUUU��        ��UUUUUUUUUUU�UUUU��        ��UUUUUUUUUUU�UUUU��        ��UUUUUUUUUUU�UUUU��        ��UUUUUUUUUUUU�UUU������������UUUUUUUUUUUU�UUU������������UUUUUUUUUUUU�UUU������������UUUUUUUUUUUU�UUU������������UUUUUUUUUUUU�UU���        ���UUUUUUUUUUU�UU���        ���UUUUUUUUUUU�UU���        ���UUUUUUUUUUU�UU���        ���UUUUUUUUUUU�U�����      �����UUUUUUUUUU�U�����      �����UUUUUUUUUU�U�����      �����UUUUUUUUUU�U�����      �����UUUUUUUUUUU��������  ��������UUUUUUUUUU��������  ��������UUUUUUUUUU��������  ��������UUUUUUUUUU��������  ��������UUUUUUUUU�  �����������������UUUUUUUU�  �����������������UUUUUUUU�  �����������������UUUUUUUU�  �����������������UUUUUUU�    ����������� �����UUUUUU�    ����������� �����UUUUUU�    ����������� �����UUUUUU�    ����������� �����UUUUUU�    �          � �  ��UUUUU�    �          � �  ��UUUUU�    �          � �  ��UUUUU�    �          � �  ��UUUUUU�  ��������������    �UUUUUU�  ��������������    �UUUUUU�  ��������������    �UUUUUU�  ��������������    �UUUUU������������������    �UUUUU������������������    �UUUUU������������������    �UUUUU������������������    �UUUUU�   �    ����������  �UUUUUU�   �    ����������  �UUUUUU�   �    ����������  �UUUUUU�   �    ����������  �UUUUU�    ������� ������ ����UUUU�    ������� ������ ����UUUU�    ������� ������ ����UUUU�    ������� ������ ����UUUU�    �    �  ������    �UUUU�    �    �  ������    �UUUU�    �    �  ������    �UUUU�    �    �  ������    �UUUU�   �      �  ���� ��  �UUUU�   �      �  ���� ��  �UUUU�   �      �  ���� ��  �UUUU�   �      �  ���� ��  �UUUU�    ������  �         �UUUU�    ������  �         �UUUU�    ������  �         �UUUU�    ������  �         �UUUUU��                 ���UUUUUU��                 ���UUUUUU��                 ���UUUUUU��                 ���UUUUUUUU�����������������UUUUUUUUUUU�����������������UUUUUUUUUUU�����������������UUUUUUUUUUU�����������������UUUUUUB      ��p          �                  �    ��@0     ��p�p    ��� �@   �~� ��   ���8q   ���p �   �p ���   �8���  �>����  ����� ���� p � ����8� /0 ������ .0 ������ Np ������p ��p�p�� ����0��� ������ ������ �� `���~���  ��np��   �r/p��  ?��p�� ����0�� ����0�0����>�>0�����~P����  �~����  �~��� ������ ��p�� ��p�  � �p�  � ���  k ��� ,���q  �0��2  �P" T�"  ��" �ZBB  �" '�D�  !$ X��   �( ���   �  F     @     @ �@     @ B@     @@f�      @@~�      @�V{      ���q      ���      ���!     ���     `��      4        �                                              �     _            :       R      �`     ��     ��     |�     ��     �     �     `     �    �    �0    �t0    �p    � �    @  � �0  � �   � �    �     �     � b    � 	B   ��   ��  `� �� 0 ��   ��� �  ����b  �o� `  �x @ ��0��@��0 @@���� �p�`�p� 0�   0�   0�   0�   �   �   �    �     �   � 0   � 0   � 0    � 0    � p    @ p    @ p    @ �    @ �      �     �     ��    � � @  p ! @ p�   p   0  8  8  �02  �p!  ϐ�  ϐ  ��*  �(  �(  `(   (   (   (              �       @   P     �    @	    �
  @
  @   P D   P ��  0     � @      @      ��      p  �(UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�jTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�jUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�jUQUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UAUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UIUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UJUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VJUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ���JUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����
UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUAQ���TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQ@��zUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ��jQQUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUU ժ~AAUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ��^EEUEEQUUATUUUUUUUUUUUUUUUUUUUUUU@��^EUUQUUAU�APUUUUUUUUUUUUUUUUUUUUUU@��^EUUPUUU�AUUUUUUUUUUUUUUUUUUUUUU@��^EUUUQTU�UUUUUUUUUUUUUUUUUUUUUU@��^DUTQAEU�AAUUUUUUUUUUUUUUUUUUUUUU@��_DUTTUT�AUUUUUUUUUUUUUUUUUUUUUPi�_U  EPi	UUUUUUUUUUUUUUUUUUUUUPY�WU  PDE�UQUUUUUUUUUUUUUUUUUU P��_UT   P T�EUUUUUUUUUUUUUUUUUUUD P��UP    @@@�ADUUUUUUUUUUUUUUUUUUT�o�UP@UUU UAV�TQTUQUUUUUUUUUUUUUU T�k�U@   @U T�j(@TUTUUUUUUUUUUUUUUUE T�Z�U@   @ �oTETTUUUUUUUUUUEEUA U�Z�VA    T @�EUUUUEUUUUUUUUUUUQT U�V�VA    @��@iP@@TTEUUUUUUUUUQT@ @U�VZ      �V�UUUUUUUUUUUAQQ @U�Vj      �k)@ @AUQDQUUUUUUTUT @AAU�Vj      P�	T   APUEUUUUUU  P@AU�UjT      d�@�  QTUUUUUUQE  PA�mU�P      �U�PDUUQUUUUQ  @UPA�iU�P     �Z(  U  @DUQUUTT     \A�jU�V@     ԫ	P @ AUAUUU T   _@UjU�Z      Y��   UUUQ T  �U@U�UU�[    ��u@)@  @P@TQEU@   pU@U�UU�kP     �Z�    TQTD     U T�VU��      �j)    T A AEU     @  P�VUz     �իPJ   @ T D Q@        @�[UP     �Z� �    @ DTQD          U}U      ���P
@     P           TUU       ��V� P    P @ EE          @UU       ��j	      P           TU        ��P        P@ @           @U         �        P                       ��P        @@    @UUU                �U         T     T��                         @@   ����                           P   @����_                               ������                      @   P@    ������W                     �@  @A    䫯���o                     �R       �ꫪ��                  �*�Z       �������   @�            ���j   P    �������   �U          
 ]U��   @    ������   �UU          )T ��V   @    �ꪪ���   hUU�        �  P�j       �����~  YTUUVe        �  @Uj   h   ������^  @V�j�U�     @~   T�    h   P�����  �U�UUU�     ��   P�    `  @�����  `UiU�VU     T��    Pe   �   �����  `UiUeYUE    T��    @e   �   ����  hUZUYeU�    T`�    @U   �   P���V   hUVUY�Ue�    T���
�
@U        U��   jUZUY�Ui�    TU`%`%@e    Z     UU   jUi�eeUY�   �eU`%`%@i    h           �U��UU�U�   �e}@@@i    h          �U�VVUeU�   ��u   @Z    �          �VVjYUiU�  @��v   TZ   �          �ZZUiUjU�  @��z   TZZ    �j          �ZZU��Z��   @���� �ZY  U  �         �jiU��V��   @��Z(�@�Zi  E �V         ���UUiUU*    ��Z(�@�Vi  UQ  j         ��UUUUU*    ���+  P�V�  U   �         ��Ve�U�*   PU�Zi U�V�  U ��        ��j��Z�
    T�k�P��V�  UA  ��j         ��j���    @y��RU��ZU  UU  �Z       ��Z��*      �u�RDQ�jUY  UUA  ���      @��jU�       �WZ����VY  UU  ��Z      @���U*        𿚢���Z  UUT    �k     @����
         <�j�껪  UUD  ��     P���           ��� *   UUU  ��     P� ��              *     UUA@A   �Z     ��                       UUUT   �[     �*                       UU@Q  �[    ���                       UUUUUA �[   ����                      UUU  �   �k��>                      UUUPE �   ��i��                      UUUUU  |   �����                     UUUU@  \    ����?             
       UUUEA     �����            �*�
     UUU      �����R          ����
     UUUUEU @   �*����Z         �*���*     UUUU  P   ���   �i         ��(���     UUUUE    �Z%   h�U         ����    UUUUA    �V��*P�_        �@U�o    UUUU @  ��_���\�z       @��TU_    UUUUA @   ��W����_Uz       Pj�    UUUU    ��U����WU�W       TU@�U�Z    UUU    �~U�j��VU�]      UZQ�Vj   UUU    Z_�^U�ZUUU      �jA �Z�   UUUU     �W��WU�jUUU     @�����   UUUQ   �VU��UU��UUU     P ����
�Z   UUU    �UU�~UU��ZUU       �JUU�Z��  UUU   `UU�_UU��VU      ��WU�j�  UUUU @  @UU�WUU�jUU      @�� @U��  UU @    UUUUUU�ZU      P �z  U�V [  UUUU@    PUUUUUeUU      ��_  P�jl UUU  �   @UUUUUUUU      ��   @��  UUUE�    TUUUUUU      P�_ �� U�   UUU �    PUUUUUU        �W���
P�   UUUD �Z     TUUUU        �_ �*PUo   UUU  j      UUUU        �U ����@U}  UUU j     @UUU        �U  ���� U�  UUU  �      TU        UuU  ���� T�Z UUU �                 PU  ���* PUU UUUE �                  T   ���
 ZUUU UU  �Z                    �
 ���UUU UUU  �j          @UU      �    �UU  UUU ��V         ���e     �    �UU  UUUU  ��V       P����         }U   UUUA  ���V      P�����Z        @WU   UUUU  ���j     �������        TU    UUUU Q  ���U    ���� ��              UUUE   𪪪VUUUU���?   �j              UUUUU  ����������:    ��            @UUUU   𫪪������      �j           �UUUUU    ��������
      ��V           �UUUUEU    �������       ��         @�UUUUU              P    ��Z        �*UUUUUQ                   ��        �*UUUUUQPA             ��j       �
UUUUUUQ           @TT    ���V      @�UUUUUUU     @PA   ���     �� UUUUUUUUE @@    UT  ���j   ��* UUUUUUUUEQ @PEUQT   ���Z @U��
 UUUUUUUUUUQP@ UUUED    ���UU��� UUUUUUUUUUQEQDAEUUUT   �������
 UUUUUUUUUUUUEAEEEQEUUUUUE   ������ UUUUUUUUUUUUUUEUTUUUUUUUU    �����   UUUUUUUUUUUUUUUUUUUUUUUUUUA    ��j   UUUUUUUUUUUUUUUUUUUUUUUUU          UUUUUUUUUUUUUUUUUUUUUUUUUUEA         PUUUUUUUUUUUUUUUUUUUUUUUUUU@       UUUUUUUUUUUUUUUUUUUUUUUUUUUU      TUUUUUUUUUUUUUUUUUUUUUUUUUUUUA @ P@ @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUTD    PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU A PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUP    DDTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUA TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUD DDUUUU2UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U]UU]�UU�UU�UuU���WU�UU�UuU�U�UU�UU����u�UU�UU��Uu���U]�U]�}U]���]�U]�]WU�U�U]�U]�]WW�u�U]�U]�]�Wu��U\�E�_wU]UpD]�]�U_U���W�U\�]WU5]]G\�U]�_WuqM]W]�T]]15]G���]U����?L UU@DT     UU       DPG 0PUu ���? u��4p7P�W0 �u� 3� q�w �?3 �|� � <��03 ��� 0��0�03 ��p�  ?���p��  � 0��5�  0  ?��10  �  0����00��  030 ��?00�    �? 0                                                                                                                                              0  0��?���?� �  �        � ��   <� <�<�0��00<00C   30 3��0� 3��00 �0k<0? � ��_W000 0 <p^�000  0�U�0030  0`Uk030�  0`uk0<0  0h�Z         hUV         jUZ         jUi&UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUAUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTDUUUUUUUQUUUUUUUUUPUDQQUUUUUUEDTUQUUUUUTUUTEUUUUUU@tEDD]u��UU5Q���u��UDpU�Q]t��_ 0P�Tu��U 0  ���_uU]EU5 �T@@�Ww ��� �u��U�? @���C4u 0  �U  0�� 0  �@0QT 0  ���?4��W 0 �� U�3 C 0 00�@?0 0 0 0 ����@��C      4          T A         @           @                     P           P                                                            "             P@             @A                                          P              @              @                                �   ��    0    0   � 0���      �� �� 0   ���? �  � 0   �   � ��?   �  ����0� 0   �  0  �0� 0   �  ��0 ��3   ��� �  �3   �   �� ��3   �   � ��3   �   �� ���3   �   � �� 0   ��� � �� 0   �   � �� 3        0 ��                                                                                                                                          "                                                                                                                                         �  0    �    ��? 0 � ��     0  �       �     3 ��   ������� �     �����0�     � 0 ��    � 0  3�   �     3�    ��? ����3�    ��0�?� ��    ��0 �  �    ��0   � �   ���������            0                                                                                                                                         ?���           ���           ���           ���           �~           ��^            ��            ��            ��            �            �V             �             U                                                                                                                                                                        0           00          ��          �0      0�<� �   <�0 � �   ��� �  Z � 0�� �  [� 3  �� �  [  3  �� �  [ ��  ?�� �   ��  3�� �   0  ��� �    �������     �3 ���  �   �  �  �                                                                                                                                                                                                                                                                                                                                                                              $UUUu}UUUUUU�UUUUUU�W�UUUUU=W�UU�U�__UUUW�WUU�U ��UU}U  �WUWU� �UUW�3 �pUU��   \UU�<   pUU5 � �WU5 ����UU��0�_UUU�0 �WUUU�  �_UUU<��WUUU���_]UU��?�W}UUU����W�W�?�_U_�?��_�����U���?  �]��?�U������p���U���U�UU����]�UU������UU�����UU]���?UU}����_UU�W�_�UU]�_��UUU����UU$U}UUu}UUU�UU�UUU�U�WUUUu��?��U�_5���UuU� �_Uu=��UU�� U�   ��U�   0|UU    _UU����UUU����WUU5�<\UU  ��WUU_�UUU����_UU�u���WUU�W���_UUU��?�WUU��?��_]U_���W�U��� _�_���  |�_UU? _UUU??_��UU���sU�UU���_��UU���U�UU����w�UU��?���UU�����UU�����U��U�W�_U��W�w�UU����_UU$��U}U�WUuU��U�UUu���UU�����sUU��? �]U�  �  �WU   ��WU   �UUU�   _UUu� �|UUU}�  �UUUU  _UU]�  �UUU�� ��WUU ��UUU��UUU��?�_UUUu���WUU�U���_UW�_���W�WU���_�_����WU_��� _�]�<  U�5? \��U5??WUU����_��U����_U�U��?���U5��?���U���?��U�����?U�����_��_��W�_��WU�wUUU���_UU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �(��� U�ZQ)YU  �U�Ue��Z���B T �Vj��PY�jU*YU�  � �Ve
j�Z�� BBe �Zi� ��ZU�ie*YU� �jd�Re���V�� @VjEA�Zi� ��ZU���*YU� hj��Re���V�� P�jU���i� ����j��iYU� hjj�Re`�jZ�� @V�Z����� �Y���ZhiYU��hjEZ�Reh�Zj�� Pf��VY��� �i�jUjZ�UU��jjEZ�Re!h�ZjZ�
 T�U�����U� ��jUUjZ�UU��j�UV�Re Y�V�V�F�d��U����U! ��ZUUVV�UU`�j�V�bU`Z�V�V�V� ��jU�ZV�U! i�ZUUUU�UU`�j�V�bU`V�Z�V�V� ��jUUjZ�U! Y�VUUUU�UU`���%V�*�V�Z�V�V��d�ZUUjV�V% Y�VUUUU�TU ����V�&`U�Z�V�Z��d�ZUUjV�V�Y�VUUUU�TU h���U�*`U�Z�V�Z�f�ZUU�V�V%�Z�UUUUU�TU*X��fU�*hU�Z�VUZ� j�VUU�VUZ$�U�UUUUU�PUX��jU�*iU�ZUUUi�VUVUU�UUj$�UUUUUUU�XUXi�fUU*YU�VUUU��VUUUU�UU��UUUUUUU�XU
Xe�jUU
ViU�UUUU�VUUUU�UU���UUUUUUU��U�YUUUUUi�ZUUUUUU�ZXVUUUUUUU���UUUUUUU��U�YUUUUU��YUUUUUU�j�VUUUUUUU��eUUUUUUUU�T�ZUUUUU��UUUUUUU�j�VUUUUUUU��eUUUUUUUU�T�VUUUUUUjUUUUUUU�j�VUUUUUUU��eUUUUUUUU�T�UUUUUUUjUUUUUUU�j�VUUUUUUU��eUUUUUUUU�U�UUUUUUUiUUUUUUU�j�UUUUUUUU�jjUUUUUUUU�U�UUUUUUUYUUUUUUU�j�UUUUUUUU�jVUUUUUUUU�T�UUUUUUUUUUUUUUUUj�UUUUUUUU�jVUUUUUUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUUjVUUUUUUUU�T�UUUUUUUUUUUUUUUU�YUUUUUUUUU�VUUUUUUUU�T�UUUUUUUUUUUUUUUU�ZUUUUUUUUU�VUUUUUUUU�TYUUUUUUUUUUUUUUUU�ZUUUUUUUUU�UUUUUUUUU�TZUUUUUUUUUUUUUUUU�ZUUUUUUUUU�VUUUUUUUU�XVUUUUUUUUUUUUUUUUUZUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUTUUUTUUUTUU��FUUUTUUUTUUUTUUUTUUUTUUUTUUTUTUTUTUTQTU�VTUTUTUTUTUTUTUTUTUTUTUTUTEEEEEEEEEEEEEjEEEEEEEEEEEEEEEEEEEEEEEEEETTTTTTTTTTTTTjTTTTTTTTTTTTTTTTTTTTTTTTTTDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                                        QQQQQQQQQQQQDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       
                                                                              *                                       b                                      �*                                      ���                                     V�*                                   �"VU�*                              ����Z FUU�*                            �jUUUU�@UU�*                          �ZUUUUU� PUU�*                        �jUUUUUUZ  TUU�                       �VUU  @�Z   TUU�                      �ZU     h    UU�*                     jUU      �`    TU�                    �VU       ��
    @U�*                   ZU       �"     TU�
                 �V       @
*      UU)                �VU        �&      PU�                jU         &       U�              �VU          �&       TU
              �U          j)        U)              h           Z        T�              Z          $�        P�            �V          (U�U       @U
            �U           	�UU       T)           �V         @��VUU       P�           �U        UU�VUU      @�          ZU       @UUU�U�VEUU      U
         �V      @UUUUUUUfZUUUU      T)         �U       TUUEUU�UfUUUUU     @�         j      @UUUUU�UUUUUUU     @�       �V      UUUUUUUUUEUUU      U       hU      TUUUUU�UUUUUUUU     T       j     @UUUUUUU�UUUUUUUU     T
      �V     TUUTUUUUUUUUUUQUU     P�     �jU     @UUUUUUUUUUUUUUUUUUU    P�    �jU    PUUUUUUUUUUUUUUUUUUU    @�   �UU     TUUUUUUUUUUUUUUUUUUE     U   ZU     UUUUUUUUUUUUUUUUUUUUUU     T
  �VU     @UTEUUUUUUUUUUUUUUUUUUU    P)  �U     TUUUUUUUUUUUUUUUUUUUUUU    P�  ZU     UUUUUUUUUUUUUUUUUUUUUU    @� �VU    @UEUUUUUUUUUUUUUUUUUUUUTU     ��U     PUUUUUUUUUUUUUUUUUUUUUUUU    TjU     UUUEUUUUUUUUUUU@UUUUUUUUQ    T�VU     @UEUUUUUUUUUUUUUUUUUUUUUUU    �U     TUUUUUUUUUUUUUUUUUUUUUUUEUU     jU     UUUUUUUUUUUUUUUUUUUUUUUUUUU    VU    PUQUUUUUUUUUUUUUUUUUUUUUU   �VU     PUUUEUUUUUUUUUUUUUUUUUUUUUUU   �U     UUUUUUUUUUUUUUUUUU@UUUUUUUUU  �ZU    @UEUUUUUUUUPUUUUUUUUUUUUUUUU� hU @ PUUUUUUUUUUUUUUUUUUUUUUUUUUUU���ZU    TUUUUUUUUUUUUUUUUUUVUU������* (�V@  UUUUUUUUUUUUU@UUU������    �
(��U@  AUUUUUUUUUUUUUUDUUU      ����*��jUA @PUTQUUUUUUUUUUU@UUU���� �����((�������jUUUUYU������jUUUUU���������*�        �������     ��
�ZU    ��*�"��(�������
       �*        �����������*���������     ������������  ��*   �����
(�*�����������������������������������* ���������������  ������������������
�����������*  �
�����������*�����������������������������������������(P�@������� U�ZQ)YU  �U�Ue��Z�� ��P����j��PY�jU*YU�  � �Ve
j�Z��P�������i� ��ZU�ie*YU� �jd�Re���V����������i� ��ZU���*YU� hj��Re���V���U������i� ����j��iYU� hjj�Re`�jZ������������ �Y���ZhiYU��hjEZ�Reh�Zj��V��������� �i�jUjZ�UU��jjEZ�Re!h�ZjZ�Vi�V���*��U� ��jUUjZ�UU��j�UV�Re Y�V�V�Ui����Z��U! ��ZUUVV�UU`�j�V�bU`Z�V�V�Ui����V��U! i�ZUUUU�UU`�j�V�bU`V�Z�V�Ue�Zf�V��U! Y�VUUUU�UU`���%V�*�V�Z�V�UUUZj�V`�V% Y�VUUUU�TU ����V�&`U�Z�V�UUUZV�V`�V�Y�VUUUU�TU h���U�*`U�Z�V�UUUj	��V`�V%�Z�UUUUU�TU*X��fU�*hU�Z�VUUUUjI��Z`UZ$�U�UUUUU�PUX��jU�*iU�ZUUUUUUjiV�Z`Uj$�UUUUUUU�XUXi�fUU*YU�VUUUUUUj�V�ZhU��UUUUUUU�XU
Xe�jUU
ViU�UUUUUUU�jUU�&ZU���UUUUUUU��U�YUUUUUi�ZUUUUUUUUU�ZUU�&ZU���UUUUUUU��U�YUUUUU��YUUUUUUUUU�VUU�&VU��eUUUUUUUU�T�ZUUUUU��UUUUUUUUUUUUUU�*VU��eUUUUUUUU�T�VUUUUUUjUUUUUUUUUUUUUU��VU��eUUUUUUUU�T�UUUUUUUjUUUUUUUUUUUUUU�fUU��eUUUUUUUU�U�UUUUUUUiUUUUUUUUUUUUUU�jUU�jjUUUUUUUU�U�UUUUUUUYUUUUUUUUUUUUUU�jUU�jVUUUUUUUU�T�UUUUUUUUUUUUUUUUUUUUUU�jUU�jVUUUUUUUU�T�UUUUUUUUUUUUUUUUUUUUUU�jUUUjVUUUUUUUU�T�UUUUUUUUUUUUUUUUUUUUUUUZUUU�VUUUUUUUU�T�UUUUUUUUUUUUUUUUUUUUUUUUUUU�VUUUUUUUU�TYUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUU�TZUUUUUUUUUUUUUUUUUUUUUUUUUUU�VUUUUUUUU�XVUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUTUUUTUUUTUUUTUUUTUU��FUUUTUUUTUUUTUUUUTUTUTUTUTUTUTUTUTUTQTU�VTUTUTUTUTUTUTUTEEEEEEEEEEEEEEEEEEEEEEEjEEEEEEEEEEEEEEEETTTTTTTTTTTTTTTTTTTTTTTjTTTTTTTTTTTTTTTTDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                                        QQQQQQQQQQQQDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������                         �UUUUUUUUUUUUUU                         jUUUUUUUUUUUUUU                        �ZU             �
                     �jU                                  �UU              (JU                  �U               �
�                 �V                "                �Z                 **�                �U                 (b�                j                 �����               �V                 U�����
             �U     @QUUUUUUUUUUUU��XU��            Z     UUUUUUUUUUUUUU���UU�
          �V    PUUUUUUUUUUUUUU��TUU�         �U    TUUUUUUUUUUUUU �� UUU
         h    @UUUUUUUUUUUUUU ��V  @U�
        Z    UUUUUUUUUUUUUUU ���j  TU�      �V   PUUUUUUUUUUUUUUU 	�(�  @UU
      �U   TUUUUUUUUUUUUUUU@�*
�   TU�     �U    UEUUUUUUUUUUUUUU����    TU
     �U    UUUUUUUUUUUUUUUU����j    @U)     h   @UUUUUUUUUUUUUUUU��
�`     T�
    X   PUUUUUUUUUUUUUUUU�  (�h     @U�   Z   TUUUUUUUUUUUUUUUU&   �X      UU
   V   TUQUUUUUUUUUUUUUU&�� �      PU�  �V   UUUUUUUUUUUUUUUUU&����       T� �U   @UUUUUUUUUUUUUUUUU�  ��       @U
 `U   @UUUUUUUUUUUUUUUUU� h!        T) h   PUUUUUUUUUUUUUUUU�Z�Z       P� Z   PUUUUUUUUUUUUUUUUUZ��ZUU      @�*V   TUUUUUUUUUUUUUUUUUU��!hUUU      TV   UUUUUUUUUUUUUUUUUU���ZUUUU     @�V  @UEUUUUUUUUUUUUUUUUU��TUUUUU     �U  PUUUUUUUUUUUUUUUUUUZ�VUUUUUUU    @aU  PUUUUUUUUUUUUUUUUUU�*VUUUUUUUU   @`U   TEUUUUUUUUUUUUUUUUU  VUUUUUUUUU   @hU   TUUUUUUUUUUUUUUUUUU�*VUUUUUUUUU  PX   TUUUUUUUUUUUUUUUUUU �VUUUUUUUUUU  X   UUEUUUUUUUUUUUUUUUUUUUUUUUUUUUU Z   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUV   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUV   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUV  @UTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUV  @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUV  @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUV  PUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�V  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U   PUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U   TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U   TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U   TUUUUUUUUUUUUUUUUUUUUUUU@UUUUUUUUUU�U   UUUUUUTUUTUUUUTUUUUUUUUUUUUUUUU�U   UU�ZUUETUUETUUUUETUUUUUU@UUUUUUUUU�U   U�
hUUTUUTUUUUTUUUUUUUUUUUUUUTUaU   U� �UUUUUUUUUUUUUUUUUUUUU@UUUUUUETUaU   �*��UUUUUUUUUUUUUUUU��UUUUUUUUUUTUaU   ���UUUUUUUUUUUUUUU��UUU@UUUUUUUUUaU   �
��UUUUUUUUUUUUUUU	�UUUUUUUUUUUUUbU   ��`UUUUUUUUUUUUUUU��UUUUUUUUUVUUUa   �
��UUUUUUUUUUUUUUUU�`UUUUUUUU�����j   ���UUUUUUUUUUUUUUUU�����������    `   �*��UUUUU�UUU�U�UUU��          ���
��
��*� ��
����������������������������*      �
(                �������     ���������������������������� ����������"�  *�����
 ��**  **    **  ���������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUU  PUUUU�?�SUUUU���CUUUU���OUUUU���OUUUU���OUUUU���OUUU0�PUU�����UU?��� ?T�������TU?0<<T�????�Pu<0SuS�?�L1S�_ 0@�TU_���C=P�?<��S}�<??�3_]����0\}��C��3_UP0PUP�P� UUU�C�CUUUU�O�PUUU @  TUU��O��TUU��L��TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   TUUUU���TUUU���PUUU ���@UU?����U����<Tu<�����PU?����S�<���P��333�S]��3?? S� �  �P��� ?�TU���<P�?��� �S}� � �3_]����0\}����0\$UWUUUuU}�UU�w_]�UU�u]}�UU�w_�?UU�WU��?|UU��?|U������U������UU����|UU����|UU��0|UU��<|UU ��@U������U��3��WU�3�_UU����WUU� 3�TUU��?TUU� ?�TUU��?TUU 3 UUU��?TUU�?�TUU����TUU��?TUU< UUU< TUU� 3�TUU����TUU< TUU<UUU   @UU����OUU����LUUU���TUU���PUU���SUU���SUU���SUU���SU �� @�<���O�033�@���3?O��� �1 ���0�??���?<����?����?<� � <������<� � <� ��� ��PU��SUU��PUU� <PUU� <PUU� SUU���SUU� <PUU� <TUU    UU���?U#UU���TUU���PUU���SUU���SUU���SUU���SUU��PUUU<��TU@033@��3?�O��3�@��� O���1 ���0�??���?<����?����?<� � <������<� � <� ��� ��PU��SUU��PUUU� <PUU� <PUU� SUU���SUU� <PUU� <TUU   PUU� �CUU�� �UU���?UU1333UUUUUUUUUUUUUUUUUUUUUUUUUUU  TUUUU���TUUUU���PUUUU���SUUUU���S UUU<�<UUU��� U�U����T����?<�T�����3�T�_��<�?T�����U�U �? T�������TUu�� 3 TUu]��?UUu} 3 TUUU����TUUU�?�TUUU����TUUUU��TUUU� ?UUUU  TUUU���TUUU�  <TUUU�  <PUU�� SU������SUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�W�?�OUUUW���P�_���?�SW���?�P����?<SU�����S? �?���P�������P�����?S� ��?W3������T��� ?�<T<����<P���� S�������SUUUUUUUUUUUUUUUUUUUUUUUUUU  PUUUU�?�SUUUU���CUUUU���OUUUU<�OUUUU���OUUUU���OUUU�?�PUU�����UU��3��?T��3� �TU�?0<T�<  �Pu 00 S��?��P� 0 �TU���<P�?<��S}�<??�3_]����0\}����3_U  0PUP� � UUU��CUUUU��PUUU    TUU����TUU����TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  TUUUU���TUUU���PUUU ���@UU?���U����<Tu<�����PU?�����S�����P����<�S]���<? S��� �P��� ?�TU���<P�?��� �S}� � �3_]����0\}����0\UUU��?UUUU���?TUUU����TUU_��TUU]���TUU_���?TUWU��? T��?���T��?<3�T�UU53��P]�_��?�S}u]U��SUU����?PU���?�@Uu}U���OU�]U�@UU�W���SUUUU�@UUUU���OUUUU��OUUUU��<OUUUU�?�CUUUU��PUUUU��TUUUU PUUUU��SUUUU��SUUUU��PUUUU��@UUUU�LUUU����O	UU��?UUUUU��?TUUUU����TUUUU�?�TUUUU��?�TUUUU����TUUU ��? PUU���?�SUU?<3?PUU��<3��SUU������OUU��3��UU��?00UU�  3 �UU� ���T�� ? ��P��<����S}�� 3��_]������\���?���_U  ��  PUU��?TUUUU< TUUUU< TUUUU� 3�TUUUU����TUUUU< TUUUU< UUUUU    @UUUU����OUUUU����LUUUU���SUUUU���CUUUU���OUUUU=��OUU�W=��OUUuW���CUUU���� T�������T]}�3��P]_U3���SUW����SU_wU��PUU����TU���� PU��W���SU��U� PUUuU���TUU�U � PUUUU���SUUUU��SUUUU��SUUUU��PUUUU= TUUUU= OUUUU� 0 UUUU���?UUUUU� ?UUUUU= UUUUU= TUUU� <�TUU��<��T#UU���WUUUU���WUUUU���_UUUU=��_UUUU=��_UUUU���SUUUU���SUU�U���PUU�U�3� U��3��?U��?��� TW_UU�0�T��_U�3�T��]U��?T�W�?��UU��� 3 TUu����TUu}� 3 TUU]��?UUU} 3 TUUU����TUUU�?�TUUU����TUUUU��?TUUUU�UUUUU�SUUUU5 @UUUU�?�OUUUUU?�OUUUUU�UUUUU��3TUUUU���TUUUU��TUUU���TUU����TUU���TUU���PUU���SUU��SUU��SUU���SU ��� @�����O���<�@����<O����1 ��0�?����? � ��?����?<� � <������<� � <� ��� ��PU��SUU��PUU� <PUU� <PUU� SUU���SUU� <PUU� <TUU    UU���?UU1333U#UU���TUU���PUU���SUU��SUU��SUU���SUU���PUUU���TU@��<@���<�O����@��� O���1 ���0�?��?�? � ��?����?<� � <������<� � <� ��� ��PU��SUU��PUU� <PUU� <PUU� SUU���SUU� <PUU� <TUU   PUU� �CUU�� <UU���?UU1333U!UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U=UUUUUUUUUUU�U=W�OUUUUUUUUU���T�3UUUUUUUUU�����<TUUUUUUUU�����PUUUUUUU������SUUUUUUU�����PUUUUUUՏ����pUUUUUUկ��ϣ���UUUU�����������UUU���߳������WUկ��������Ã_Uռ�������3���^Uճ��������ˏ{U������<�:����U�������*��/zU��������*�+?_U����2���+��+?WU믪��<�+?�*<UU뭪��<�-?���UU}��
��<�-?���UUU�*���<z5<���UUի��|�<_�<���WUժ�_�<UU��_�WUU�U�_U�WU�WU�_UUUU�WU�U_UUUUU�U��U_]U_}UUUU�U�W��W}�U�!UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU]UuUUWUUUUUUUUU}U�U�_UUUUUUUUU�U�U�_UUUUUUUUU�U�W�sUUUUUUUUU���W�|UUUUUUUUU�����|UUUUUUUUU�����UUUUUUUUU�����_UUUUUUU_��Ï��PUUUUUU�_��Ϗ��sUUUUUU�_��Ϗ���UUUU����������UUU���߳��+��ˏWUկ���#��+?�ˏ_Uժ���#��*?�
�^Uի���0��*?�+?{U��������*<�+?�U���������<�/?zU���������+�\U����2�����\U믪������TU뭪*�������WU}���_������WUU���w5�0��/�_Uի
�]U�u�
Uժ�_W��U_ML_}UU��UU�W��W}UW�                                                                                                                            DUUUUUUUUUUU����UUUUUUUUUUUUUUUUU   _UUUUUUUUUUUUUUUU5 � pUUUUUUUUUUU���U� �?�UUUUUUUUUU�����WU �WUUUUUUUUU�����U �\UUUUUUUUU�����U�  �pUUUUUUUU��0 �U �UUUUUUUU���� �U� ��UUUUUUUU����? �_U��WUUUUUUU��������UU5�WUUUUUUU������? �WU5�WUUUUUUU�?������_U5�_UUUUUU��?�_���?�U��UUUUUU��?�WU����U���WUUUUU��?�UUU���_���_UUUUU����WUU��� �����_UUU���_UUU���?����sUUU���UUU��?������UUUU���UUU���0�W���UUUU����WUUU����U��UUUU��?�WUUU�����U��UUUUU��� _UUUU���U�WUUUU���UUUU���_U�\UUU�_���UU�_���WUs5\UUU����?�WU�U��UU��_UUU������_U��UUUUUWUUUU����� ���WUUUU�UUUU�����������_UUUUUUUUU������?����UUUUUUU�W����� ����UUUUUUU��W����  ��_�W�WUUUU���UU��  ��W�_�\UUUU��UU��   �U���pUUUU�UUU�    �UU��pUUUUU�UUU5    �UU�_UUUU���UUU5    �UU�UUUUU5p�WUU     W���UUUUU5\WUU� �W�_WUUUU5WWUU3 �_�WUUUU���UU��� ??\�s5WUUUUUUUU���?���p���UUUUUUUUUU���?���sWUUUUUUUUUUU�����?�sWUUUUUUUUUUUU�����pWUUUUUUUUUUUU�� ��0pWUUUUUUUUUUUU� �0 pWUUUUUUUUUUUUW�3\WUUUUUUUUUUUUW WWUUUUUUUUUUUUW� 3WWUUUUUUUUUUUU]5�0 WWUUUUUUUUUUUU]5   �UWUUUUUUUUUUUU]50  ��UWUUUUUUUUUUUU]500����UUUUUUUUUUUUUu5���0��UUUUUUUUUUUUUu� ����UUUUUUUUUUUUUu� <�p�UUUUUUUUUUUUU�U3�puUUUUUUUUUUUUU�U \uUUUUUUUUUUUUUUW5?�WuUUUUUUUUUUUUUU]����U]UUUUUUUUUUUUUUu}�?\_WUUUUUUUUUUUUUU�W W�UUUUUUUUUUUUUUUUU��WUUUUUUUUUUUUUUUUUU WUUUUUUUUUUUUUUUUUU5�UUUUUUUUUUUUUUUUUUU�pUUUUUUUUUUUUUUUUUUUU_UUUUUUUUUUU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUU��UUUUUUUUUUUUUUU���_UUUUUUUUUUUUU����UUUUUUUUUUUUU��  UUUUUUUUUUUU?   pUUUUUUU�UUU��   �U��UUUU��WU��   ���pU�WU5��U��   < 7�W5\U5�_=   � ���U p�     �� ���5 ��00     ����< �� 00     ����������0    ��������Us�     ���������U}U 0   ��������UUU?�   ��������UUU�?   ���������UUU�?   0 �?�����UUU�       ����UUU�   �?   ����UUU��  �U��� ����UUU��  �U�_U���?UUU=p� ����UUUU���UU_\U����UUU���_UU�WUU���_UUU���WUU�UUU�_�WUUU���UUU�pUUUU��_�WU��UUU=pUUUU5�����_UUUpUUUU\�����UUUU��UUUUW�����UUUUUUUUUU���_��WUUUUUUUUUUUu5pU�UUUUUUUUUUUUU�_���UUUUUUUUUUUUUUU5p�WUUUUUUUUUUUUUU5\WUUUUUUUUUUUUUU5WWUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU1UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU}UUUUUUUUUUUUUUUUU_UU}UUUUUUUUUUUUU��_��WUu�WUUUUUUUU� �7�UU�sU�WUUUUUU=�< �� pU\UUUWU����  \� pUUU\U?��������p=��UUUp�������������WU�����������������_���������������� ���������������� ����� �����������?���� ���������������   �  ����������<   0  � ������? 0��0  �  �?���� �U��     ��� �WUUUU��� �  ��? UUUUUUUU�0   �?�UUUUUUUUUU��  �3|UUUUUUUUUUUU�? ��WUUUUUUUUUUUUU���_UUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUU_U�UUUUUUUUUUUUUU����UUUUUUUUUUUUUU5���UUUUUUUUUUUUUU5���UUUUUUUUUUUUUU���_UUUUUUUUUUUUUUU��WUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUU�UUUUUUUUUUUUUUU��pUUUUUUUUUUUUUUUs5pUUUUUUUUUUUUUUU]\UUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU1UUUUUUUUUUUUUUU���UUUUUUUUUUUUUU�  �UUUUUUUUUUUUUU ? pUUUUUUUUUUUUUU� \UUUUUUUUUUUUU��?  WUUUUUUUUUUUUU5� �UUUUUUUUUUUUUU��  |UUUUUUUUUUUUUU� �WUUUUUUUUUUUUUU�? |UUUUUUUUUUUUUU����WUUUUUUUUUUUUUU�?|UUUUUUUUUUUUUUU��WUUUUUUUUUUUUUUU���UUUUUUU�_UUUUUUU��sUUUUUWUWUUUUUU���_UUUUU\�\UUUUUU=��WUUUUU�5��UUUUU���UUUUUU��_UUU����_UUUUUU����UUU���UUUUUUU���? �����_UUUUUUU���������UUUUUUUU����������_UUUUUUUU����������UUUUUUUUU���������_UUUUUUUUU?�������UUUUUUUUUU�������WUUUUUUUUUU �������UUUUUUUUUUU  �����_UUUUUUUUUUU������_UUUUUUUUUUUU�U���UUUUUUUUUUUUU�U��}UUUUUUUUUUUUUUUU��_UUUUUUUUUUUUUUUU��sUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUU�\UUUUUUUUUUUUUUUUs5\UUUUUUUUUUUUUUUU��_UUUUUUUUUUUUUUUUWUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU$UUUUUUUUUUU��UUU�UU��WUU�_U3?\UUw��30pUUw��0�UUuw7 �_UUw �\UUu   \UUU=   \UUU5  �WUUU�  �UUUU� <WUUUU �]UUU��0sUUU�?0pUU��<���UU�����UU�����_UU5�?�_UU5��<�UUU=���pUUU=���pUUU� ��pUUU�0��|UU������UU=  _U� p�  �p�   �� p�      \U     WU=   ��UU� �WUUUU��UUUUUUUUUUUU$UUWUUUUU��U�UWUU�U��U�UUU����UU��? �WUU� 3 WUU�   ��UU 3 ��UU�  �WU��� �UU�00? _U�    |UU�   �WUUw  \UUUU30|UUUU=�<�UUUU���|UU�_=��_UUu]���UU�_� �_U]��  U]��� \U_�?�� U}U����_UU���U�U����_UU����WU�W����_U������WU��?���WU�����?WU������UU�����sUU��?��_UUU����]UUUu��UUU$UUU�W}UUU�wUU�_�WW��C�W]�  <�u5  ?��53  |}5  \W53  � 0 � 3 |� � _��  W�03  _�?   WU ��_U���U�3��_U���3W�_���_�����U����_����W��� _u��  �UU� U_��_�}?��U��0��U��  U��  \U_?< UU���_}����W�����WU�}��U-UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUWUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��uUUU��UUU��UUUUUU��UUUUUUUUUUUUUUUUUUUUUU����WU����UU��]}UU���WUUUUUUU����VWUUWU�_U�����������U������U����~UUUUUUUݏ����UU����翪��.Ŀ��+���������������WUUUUU�����������+������������8ȯ�������������_�����ꎫ������������"��*���" * : � (�������������*�
*(��� ���**2�� �  @�
(  (�2 �� �: �
�� �� ��    � � ��   "     �  � ���" (  �   ��*      �         �        ��    "�             @            PU ��  @�  TUU @U U@UAUU  P�TUEP @ UUU PUUUPUUUUUUUUUUUUUUUUUUPUUUUUUUUUUUEUUUUUUUUUUUUUUUUUU	UUUUUUUUUUUUUUUUUUU��UUUUUUU��]}UU�������U����������ȯ�������" * : � ( @�
(  (�   "       �         @UU @U U@UUUUUUUU	UUUUUUUUUUUUUUUUUUUUUUUU��_W_UU�����U����������������������
��*����
 
��   �0    �        P   P@PUPAUUUUUUUU	UUUUUUUUUUUUUUUUUUUUUU��_UU�WUU��zUU�_���(�WU��������*���������
�"*�� �(� 2        �          T   TPTTUUUUUUUUUUU	UUUUUUUUUUUUUUUUUUUU��WUUUUUտ�^UUUU��*
�UUUU���*��_UU�*��*������������� � ���   � �     �   U     TUUU  UUUUUUUAU	UUUUUUUUUUUUUUUUUU��UUUUUUU��WUUUUUU��~UUUUUU����WUUUU������_�����������2 �� �: �  � ���      �       UAUU  PUUUUUPUUU$UU�_UUUUU��UUUUU  _UUUU\�UU� � �uUU= <�]UU    WUU���? �UU���� UUuuu�sUUUWW��UU�����U�=�� ps���   \=�U  _�U �u_��W��W�3��UU��|�WU����_�|UU��UU�pU�?_UU��u?�WUU����]UU����UUU���_UUU��=�uUUUU���UUUUUU�UUUUU���UUUUU��UUUUU��_UUUUU����UUUU��}WUUU��__WUUU����UUUU���WUUU$UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUU�U��UU��U  _U50U\]� ��u=3= <�]7�    �?���? ��W���� ��uuu��?�UWW��w�������]��=�� p�?�   \=0�U �_���U �U��U��WU���UUUU3��UUUUU3��UUUU]<�UUU]��UUU��1�_UU��3�wUU����WUUU=���]U$UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUU]U��UUUuU �_WU�U\]��� ��u=�= <��?�    �����? ������� � uuu��UWW��W?�������0=�� p�0��   \50�U �_5��U �U�0U��W�UUU�<��(
UUUUUUUUUUUUUUUUU�WUUUUUUU� |UUUUUUU �WUUUUU�   \UUUUU=   pUUUUu��UUUU��u�}UUUU��WUUUUUUU5�UUUUUUUU5�UUUUUUUU=�UUUUUUUu?�_�]_UUU�� �0�|UUU�� � �UUU��   �UU��w < pUU��w  \UU��5�  WUU�|u�  �WU��_UU |UU��_UU��WUU��WUUUUUU���UUUUUUU��WU�WUUU�0�WUUUU�_�0�WUU���_5�WUU<���UUU��� �UUU=���?UUU� ����WUUUU���WUUUUUUU��_UUUUUU_��_UUUUUU_��}UUUUU}���UUUUU�����UUUUU�?��wUUUUUU?��UUUUU(UUU�U�WUUUU�U�_UUUUW5\UUUU�U�UUUU�U5�UUU� W WUU��U WUU��W= _UU5 \5 \UU5 W\UU5�U\UU��W\UU� \50\UU� \50_UU�W= WUUU_�WUUU��UUUU=  �UUUU� _UUUUU�WUWUU�=]U�UU]��wU�_UU�_UU�|U���U�pU��5�W��u?�|������p���u?0|��W _��=U��WU���U�UUU�_WUUUU��_UUUUU��UUUUU��_UUUUU����UUUU��}WUUU��_WUUU����UUUU���WUUU(	UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��_UUUUUU= �UUUUU� �_UUUU�  |UUUU= � �]UUU < �uUUU   ��UUU=�? wUUU���� _UUUUuu��UUUUUUU�WUUUUUU�_U�UUW�����u������=���� p���   \U���5  �_��3�� �U��|U=�U���_U��UU=UUU]UU��_UU��_U��WUU� |U?�UUU�0���UUU�����_UUUU���wUUUU=���UUUUU����UUUUUUU��UUUUUU��UUUUUU��_UUUUUU����UUUUU��}WUUUU��__WUUUU����UUU$UU�_UUUUU� �UUUUU  _UUUU \�UU� � �uUU= < �]UU    WUU���? �UU���� UUuuu�sUUUWW��UU�����U�=�� ps���   \=�U  _�U �u_��W��W�3��UU��|�WU����_�|UU��UU�pU�?_UU��u?�WUU����]UU����UUU���_UUU��=�uUUUU���UUUUUU�UUUUU���UUUUU��UUUUU��_UUUUU����UUUU��}WUUU��__WUUU����UUUU���WUUU UU}_UUUUU��UUUU�3 WUUU�0 \UUU=  pWUU=33�WUU�UUU33�UU�   �UU���p]UU���WU� 0�UUU� UUU��UUU����UUU��?�WU�<��UU5�� �UU�pUU5<� �UU��  �UU����UUU�?@UUU� �WU��U� � �U�0� ��U�3  �U?��U �0�U���� U���UU UU�}UUUUU��WUUUU� \UUUu� pUUU�  �]UU����_UU5000WUU��WUU  �WUU���uUU3�_UU? ��WUU� �UUU5? �UUU��OWUU��PUUUU PUU��� �WU� �|U� � pU�0� ��U�3��U? 0|U �<pU5��� U�?�WUU= �UUU� pUUU���_UUU� 0\UUU5?WUUU�  WUU$UUUUUUUUUUUUUUUUUUUUUUUUUUUUU_��UUU�\5?_UU=\=pUU��UU�  wU��� �U�� ��\U�5  0\U�� �<_U��? �U�5�U��  �_U��? �WU��� �WU�u=�?\U�W��|U��< \U��� \U� �  WU��� _U� 0\UU}� ?|UUU���UUU� \WUU= \WUU� �_UU� �WWUU5 |UUUU���UUU? ?�UUU5� �UUU����U$UU��WUUUU WUUUU�UUUU��UUUU��UUUUU=|}_UUU_��UU� �3 WU=��0 \U5<<  pW�<0�W�0�U��  �U�� ��U���p]=0�� �W�  �U� � UU��UU����UU���?�WU�7��UUU���UUU�?pUUU�0 �uUU� ��UU����UUU�?��UUU  ��UU�0 ��UU�0 �UUU�� pUUU5� \UUU?� \UUU0 pUUU?��U$U�����UU��� �WU��   _U����\UU�UU�pU��}_�U� ��UUU��0 WUU��0 \UU5<  pWU5<0�WU50�UU�  �UU� ��UU���p]UU�� �WU�  �UUU� UUU��UUU����UUU��?�WUU5��UUU�� �UUU� pUUU=� �UUU�  �UUU���_UUU�?�}UUU� �uUUU ��UUU uUUU�WUUUU|�WUU��\UUU \UU��?�_$	UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU}_UUUUUUU��UUUUUU�3 WUUUUU�0 \UUWUU=  pW�|UU=0�W5�UU0�U5�UU  �U5�U� ��U5�U���p]5�UU�� �W��W�  �UU_U� UU|U��UU=�U����UU��_��?�WUUW5��UUU�?�� �UUU�� pUUUu<� �UUUU=�  �UUUU����_UUUU�?�}UUUU� �uUUUU�� ��UUUUU= �uUUUUU UUUUUU�WUUUUUU|�WUUUU��\UUUUU \UUUU��?�_ U_��UUU�\5?UU=\=�UU��WU�  wU��� �U�� ��\U�=  0\U�� �<_U��? WU�5�U��  ��U��? �WU��� �WU�u=�?\U�W��|U��< \U5�� \U� �  WU5�� _U� 0\UU�� <�UUU���wUU  �U� puU� < pUU� ��UU�|��WUU\� WU�\� WU�|0_U��_��W U_��UUU�\5?UU=\=�UU��WU�  wU��� �U�� ��\U�=  0\U�� �<_U��? �U�5�U��  �_U��? �WU��� �WU�u=�?\U�W��|U��< \U5�� \U� �  WU5�� _U� 0�_U�� ?�]UU��\}UU  \uUU \�UU _uUU=�WUUU��UUUU�0�UUU����WUUU_UU����WU U_��UUU�\5?UU=\=�UU��WU�  wU��� �U�� ��\U�=  0\U�� �<_U��? WU�5��U��  �_U��? �WU��� �WU�u=�?\U�W��|U��< \UU�� \U� �  WUU�� _U� 0\UU�� ?�UUU���WUU� \WUU=? \WUU� �_UU5 �WWUU5 UUUU����UUU? ?�UUU� �WUU����U UWUUUUUU�_UUUUUU�UWUWUU���UU]UU=��}_]UU�����_UU�����WUU=���WUU���<�_UU�s=��_UU��<�UU�_���UU�����_UU�����_UU�_���WUU�_����U���uUU����_�UU?�uU�?�?�uUU��}UU=�?�_]UU��0�]UUU=���WUUU3��pUUUU��<�UUUU30WUUU���UUUU5000UUUU�� WUUU3pUUUU��UU UWUUUUUU�_UUUUUU�UWUWUU���UU]UU=��}_]UU�����_UU�����WUU=���WUU���<�_UU�s=��_UU��<�UU�_���UU�����_UUU����UU�]���UUUQ���WUUUC���TUUU���UUU5� pUUU  0\UUU� \UUU0�UUU50 WUU WUU0<�tUU��0UUU<<\UU50WUU�0� �UUU�����UUUU1sUUUU�0\UU$UUUUWUUUUU��]UUu���WUU����_U�����U5s�s�_U=C��WU�UU]UU�}_]UU=���_UU��?�WUU����WUU����_UU�<��_UUU�<�UUU���UU�??�_UU����_UUU���WUUU���UUU��UUU���_UUU=�UUU�3�UUU�?�UUU��_U�U�30�UuU����W�U����_uU����]}U���}_U5�0\uWU=��|�W��UUU �UU�����WU$UU�_UUUUU��_UUUUU��WUUUUU�?_UUUUU��WUUUUU5�UUUUUU�_WUuUUU��UU]UU���}_]UUU����_UUU��?�WUU����WUU�_���_UU�W=��_UU=_�<�UU|���UU��??�_UU�����_UUU���WUUU���UUU���UUU����_UUUU?�UUUU�?�UUUU��UUUU�?�_UUUU�0�UUUU����WUUU����_�UU����]uUUU��]�UUU��\]WUUU�\}WUU�� \�UUUU|UUUU���_UU$UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUWUUUUUU�_UUUUUU�uUUuUU���UU]UU=��}_]UU�����_UU���?�WUU5���WUU�����_UU�s=��_UU��<�UU�_���UU��??�_UU�����_UU�_���WUU�_���UU���UU�����_UUU?�UUU?�?�UUU��UUU=�?�_UUU��0�UUUU����WUUU����_UUU��?�]UUUU��]�UUU�\}uUUU<|��UU����WUUU�<�WUUU����WU$
UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUuUUuUUUUUU�UU]UUUUUU�}_]UUUUUU���_UU�uUU�?�WUU��]U���WUU��WU���_UU��_U=��_UU���U�<�UU��|U���UU5��??�_UU�������_UUU��U���WUUU��W���UUUU?W��UUU��_���_UUUU�=�UUUU���?�UUUUU��UUUUU?�?�_UUUUU�0�UUUUU�����_UUUUU����]�UUUU��?�}uUUUUU����UUUUU�\�WUUUUU<|UUUUUU���UUUUUUU�<�WUUUUU����WU UWUUUUUU�_UUUUUU�UWUWUU���UU]UU=��}_]UU�����_UU���?�WUU=���WUU�����_UU�s=��_UU��<�UU�_���UU��??�_UU�����_UU�_���WUU�_���UU���UUU����_UUU?�UU�?�?�UUU��UUU?�?�_UUU��0�UUUU����WUUU����_�UU����]uUUU��]�UUU��\]WUUU�\}WUU�� W�UUUU� \UUUU���UU UUUUUUUUUWUUUUUU�_�UUuUU��UU]UU���}_]UU=����_UU���?�WUU�����WUU=���_UU��=��_UU�s�<�UU����UU�_??�_UU�����_UU�_���WUU�_���UU�_��?|U�����_UuU�?�U�����Uu�?��UuU���_UuU?�?���}U�����_UU����WUUU����UUUU���UUUU�p�\UUU�||UUU� W=�UUU��W5�UUUUUU��WU UWUUUUUU�_UUUUUU�uUUWUU���UU]UU=��}_]UU�����_UU�����WUU=���WUU�����_UU�s=��_UU��<�UU�_���UU��??�_UU�����_UU�_���WUU�_���UU���UUU����_UU�?�UU�?�?�U�U��UuU?�?�_U�U��0�UuUU����W}UU����__UU�����UUUU��UUUUU3�pUUUU���UUUU��W�_UUU5�� WUUU����UUU���W�U���O�U���U���s�U�p�U������<  <��<<<<��<  <��<�<w��0�wU���uU��}U���_}U5  \]U���]����_�����_�����_����?p3  0p����\<���_���U�p5 WUp��UUpUUUU�_UUUU���WUU���OUU���U���s�U�p�U������<  <��<<<<��<  <��<�<w��0�wU���uU��uU���_uU=  |}U���}U���]�����_�����_����?p3  0p����\����_��=�W��5�WUp5�UU�_5�UUUU�UU���U���U����U����U �������� �w����w� �w�? �uU?<�uU��_uU= |]U� �]U���]����_����W����_� �p����s�����WWUW�UU�UUUU�uU�u���}��]�3�]��_U|WU�_WUpWU�W���W���W��W���U�pUU_UU(eUUUUUUUUYUbUYUUUUUUUUUUUUiU�U�UiUUUUeU�UeUUUUUUUUUZ�`�dUZUUUUeU�UeUUUUUUiU�U�Ui(eUUUUUUUUYUfUYUUUUUUUUUUUUeU�UeUUUUUUiU�U�UiUUUUUU�V%X%Y�VUUUUUUeU�UeUUUUiU�U�Ui ��? ��?�����?��3?����� ��? ��? <3 <3 ��$	UUUUUUUUUU��_UUUUUU= �UUUUU� �_UUUU�  |UUUU= � �]UUU < �uUUU   ��UUU=�? wUUU���� _UUUUuu��UUUUUUU�W]UUUUU�_U�UUW�����u������=���� p��?�   \� ��5  �_���� �U�U=���UU�� ���WU�?    _U�0     s�0   0p� ��    p��    |U��  ��_�� �� �U5 �  �_5    �|�    �?p��  0 < pU? �� U�  � �W���3  |UUU�� � \U$	UUUUUUUUUU��_UUUUUU= ����UU� �? _UU� �� |uU=��� pUU� � �UU<   ��U=   ��W�   � _U �    \U �  � \U ��? ��  0 �=�    � ��   � ��    ��     �      �    ��U     ��W    � _� �   0 s� 0   0p�<0 �� p�0�    |U�   �_���� ��U5 � � �_5 � ��|�    �?p��  0  pU? �� U�  � �WU��3  |UU]�� � \U$	UUUUUUUUUU��_UUUUUU= �UUUUU� �_UUUU�  |UUUU= � �]UUU < �uUUU   ��UUU=�? wUUU���� _UUUUuu��UUUUUUU�W]UUUUU�_U�UUW�����u������=���� p��?�   \� ��5  �_���� �U�U=���UU�� ���WU�?    _U�0     s�0   0p� ��    p��    |U��  ��_�� �� �U5 �  �_5    �|�    �?p��  0 < pU? �� U�  � �W���3  |UUU�� � \U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             (
UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUU5��UUUUUUU�0�WUUUUUU5���UUUUU���?�UUUUUU� WUUUU� � �WUUU� � <|UUU�<�0 �UUU� ��� �UUU5 � � pUUU�0<0 _UUUU<�pUUUU  pUUUU3�  \UUUU��0��WUUU� pUUUU=  _UUUU�� �UUUU� 0<�UUUU� 0<pUUUU� ���_UUUU� 0 pUUUUU�� �UUUUU  WUUUU5  WUUUU�0 WUUUU5 00�UUUUU50��UUUUU� � �UUUUU��?�UU(
UUUUUUUUUUUU��UUUUUUU}5 WUUUUU�� WUUUUU5 �\UUUUU5 00\UUUUU5 0\UUUUU�� \UUUUU5�� sUUUUU5 ��p�UUUU�  3� �WUUU� ���_UUU� �_UUU ��sUUU5 � �?|UUU5 ��UUU��0�0�_UU� 0p�0�uUU� �_0|�UUU�� 0�UUU��U��_uUUUU�U=��_UUUUW0|UUUUU5sUUUUU�����UUUUU� 0� WUUUU�  \UUUU�  \UUUU� �� pUUUUU pUUUUU��0pUUUUU�0�UUUUU �UUUUU� 00�UUUUU5 00pUUUUU5 0�pUUUUU ��\UUUUU0� sUUUUU pUUUUU����(UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUpUU�WUUUUU�UU�_UU�_ WU�UU� �WU�UU 0\U���UU \U���UU \U��U�0 sU���U���pU���WW  �U��WW�  0W��UWU�0\�UU5 � \� _uUU� W5��]UUU��U�3 WUUU U?�\UUU5���� 0\UUU�_50 0pUUUUU50 pUUUUU���|UUUUUU0 �UUUUUU5���UUUUUU50 0|UUUUUU5 0�UUUUUU�0��UUUUUUU0 WUUUUUU� WUUUUU� � �UUUUUU�� 0WUUUUU�0 < WUUUUUU����W(
UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUU\UUUUUU�� pUUUUUU=< pUUUUUU� �UUUUUU �U�UUUU ��� �WUU� �U��_UUp� �_UU �U��sUU 0W�?|UU50 W��UU��0�U0�_U� �0_�0�uUU�\0|�UU�� � 0�UUW��_uUU �U=��_UU�U0|UUU5p]U5sUUU�_]����UUUUU}?0� WUUUU�  \UUUU�  |UUUU= �� �UUUU�  �UUUUU��|UUUUU �UUUUU �UUUUU� 00�UUUUU5 00pUUUUU5 0�pUUUUU ��\UUUUU0� sUUUUU pUUUUU����!UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUuUUUUUUUUUUUUUuUWU}UUUUUUUUUUUUU��_U�wUUUUUUUUUUUU��_U�_UUUUUUUUUUUU��_��_UUUUUUUUUUUU�����UUUUUUUUUUU���_�_UUUUU��w���U����+WUUU�������W���+?^UU������_�W?���+?|U���UUUUU�w?��:?�U�_UUUU�����?�.<�UUUUUU��������<�WUUUUU��>��0�����_UUUUU��:������^UUUUUë�:��(����{UUUU����:�3(?����UUUU�����0���zUUUU�����<
ϯ��_UUUU��>���<�ϫ��WUUUU�����
�����UUUUU��p<�*���sUUUUUu��
x?�?���WUUUUUU���_?����WUUUUUժ��U?��ϫ��WUUUUUU��_U_UU_���_UUUUUU�UU�_UUUU�WUUUUUUUUU�_U�UU�_UUUUUUUUU��U��UU�UUUUUUUUU��W��UU_�UUUUUUUU�_�_}�W�W�W4UUUU�U��_�UUUUUUUUUU�_U�UUUUUUUU��U]U��UUUUU]U��UU{U��_U]UU]U�WU��WU�\U]UU_UuUU��~UUWU}UUWU�UՊ��U�_UuUUWU}U����_U_UuU�WU}U����^U_U�U�W��U몮�z��U�]�WUժ����UU�W�WUի����UU�W�UU������WU�W�UU��������}U�_�U�_������W�U�_�U�_������W�U�\uU�\������W�UUW�UUW������WuU�W�WU������WU�U�wU��������_U�UU_U�׫�����WU}UU_U�_����z�]U}UU}UU����~UU_UU}W��������Uu_UU�UU�׊���WU�wUU�WU�߯���UU�WUU���W=��_���UUUU�����>���UUUUU��þ����UUUUUUUUU���SUUUUUUUUUU��SUUUUUU�����(*�����UUU����������]UU�WUU����PUU�WUU�WUU_��W}UU�WUU�UU�_��~�U�WUU�U��ժ����W�_U�}��U����W��U�UUUU����^UUUU_U_U� ;�^U}U}U�\�_U���^U�]�U�W�WU����^U�W�U�W�]U����^U�W�W�WuUU����_UUW�UU_�UU����WU�\}UU_�UU��zUU�_}U�]��U��~U��W�UU}U��_��_��_U_UUuUUUUUUUUUUUWUU�UUUUUUUUUU�WUU�UUUUUUUUUU�UUU�UUUUUUUUUU�UU<UUUUUUUU�WUUUUUUUUUUUUUU_UUUUUUUUUUUUUU}UUUUUUUUUUUUUU�WUUUUUUUU�U�UU�_UUUUUUUUU�_UUUUUUUUUU��U]UU�UUUUUUU��UU{UU�WU]UUUU�WU��WU�\U]UU]UuUU��~UUWU}UU]U�UՊ��U�_UuUU_U}U����_U_UuUUWU}U����^U_U�UUW��U몮�z��U�]�WUժ����UU�W�WUի����UU�W�WU������WU�W�WU��������}U�_�U�_������W�U�_�U�_������W�U�\�U�\������W�UUW�UUW������WuU�WuUU������WU�U�UU��������_U�U�WU�׫�����WU}U�wU�_����z�]U}UU_UU����~UU_UU_U��=�����Uu_UU}UU�Ê���WU�wUU}WU�ϯ���UU�WUU�UUU=��_���UUU�W����~���UUU����þ����UUUUUU�U���SUUUUUUUUU����UUUUUUUUU��(*��UUUUUUU���S�WUUUUUU�Uݯ��\�UUUUU�\U?��U�]UUUU�W�_��~�U�WUUUU�U�ת���W�_UUUUU������_UUUUu�Us����^s�}WUU�_U_� ;�^}U�UUU�W�_���^�U�WUU�UU_����^}U�\UU}UU����^UU_UU}UU_����_}U�_UU}UU_����W}U�WUU}UU_U��zU}U�WUUU�\U��~U�U�UUU}UUsU��_UsU}UUU�UU�WUUUUU_UUU�UU�UUU�_�WUUU�UUU�WUU�W�UUUU�UUU�_UU�U�UUUU�UUUU�UUUUUUUUUUUUUUU�WUUUUUUUUUUUUU}UUUUUUUUUUUUUUUUUUUUU<UUUUU�UUUUUUUUUUUUUU}UUUUUUUUUUUUUU_UUUUUUUUUUUUU�WUUUUUUUUUUUUU�UU�_�UUUUUUUUUUUU�UUUUUUUU�_UU]U��UUUUU]U�WUU{U��_UUUU]U�UU��WU�\UUUU_UuUU��~UUWU]UUWU�UՊ��U�_U]UUWU}U����_U_U}U�WU}U����^U_UuU�W��U몮�z��UuU�WUժ����UU�U�UUի����UU�U�UU������WU�]�UU��������}U�W�U�_������W�U�W�U�_������W�U�_uU�\������W�U�_�UUW������WuU�\�WU������WUUW�wU��������_U�WU_U�׫�����WU�UU_U�_����z�]U�UU}UU����~UU}UU}W�����>��UU}UU�UU�׊���WUU_UU�WU�߯���UUu_UU���W=��_UU�wUUU�����>��U�WUUUU��þ������UUUUUUU���SU�UUUUUU����UUUUUUUUU��(*��UUUUUUU���S�WUUUUUU�Uͯ��\�UUUUU�\U��WU�]UUUU�W�_��~�U�WUUUU�U�ת���W�_UUUUU������_UUUUu�Us����^s�}WUU�_U_� ;�^}U�UUU�W�_���^�U�WUU�UU_����^}U�\UU}UU����^UU_UU�UU_����_}UU_UU�UU_����W}UU_UU�WU_U��zU}UU_UU�_�\U��~U�UUUUU_UsU��_UsUU_UUU}UUUUU�U�_UUU�U�UUUU�_U�WUUU�U�WUU�UU�WUUU�U�_UU�WUU�UUUUUUUU�_UUU�UUUUUUU�WUUUUUUUUUUUUUU_UUUUUUUUUUUUUUUUUUUUUUU!UUU�WUUUUUUUUUUUU�?WUUUUUUUUUUUU��_UUUUUUUUUUUU��_UUuU]UU_UUUU�UUU�U}UUUUUU�U�UU�U}W�_UUUU}U�UU���U�sUUUUU�WU�����|UUUU_U�_U������UUU�WUU�U������_UU�WUU�W������PUU�UUU�W������xUU�UUU�W��ϣ���UUUU�����������UUU���_�������WUU��~�����Ã_UU��z?���3���^UUë��?����ˏ{U�����<�:����U�������*��/zU�������*�+?_U��>�����+��+?WU�����<�+?�*<UU뭪�p�<�-?���UU}��
x�<�-?���UUU�*�_�<z5<���UUի��U�<_�<���WUժ�_U�|UU=�_�WUU�UUUU|UU�UU�WUUUUUUUUU�UU�_UUUUUU��W��WUUUUUUU��_�WWU_}UUUUUUU�U_�U�!UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�]UUUUUUUuUUUUU=�UUUuUWU}UUUUU��WUU��_U�wUUU�_�_UU��_U�_UUU�WU�UU��_��_UUU�UU�WU�����UUUUU�_����_UUU_UUU�U����+WU�WUUU�W?���+?^U�UUUU�W?���+?|U�UUUU�7?��:?�UUUU�����?�.<�UUU���_�����<�WUU��>��0�����_UU��:������^UUë�:��(����{U����:�3(?����U�����0���zU�����<
ϯ��_U��>���<�ϫ��WU�����
�����UU��0<�*���sUUu��
x?�?���WUUU���_?�W���WUUժ��U��ϫ��WUUU��_U_UU_���_UUU�UU�_UUUU�WUUUUUU�_U�UU�_UUUUUU��U��UU�UUUUUU��W��UU_�UUUUU�_�_}�W�W�W8         ��         � _=          �U�          CT          L�           3          �                                                          �           �                        �            0                       �                        @           pU           ��            p            �                                                   �            `            0                                               �           �u           `�           XU           XU           XU           VU           VU           VU          @VU  @      PV�  @U     TV�   X     UVe T`    @UVe@UU�U   TUUVY���UUPUUUU��PUUUUUUUUUUV����UUUUUUUUZ�PUUUUUUUUUU�z���UUUUUUU��~@UUUUU������_ �UU���������  ��     ���8         ��         � _=          �U�          CT          L                      �                                                          �           �                        �      @   �?      @   �
      `          `          `    @     `    pU     P    ��     h     \     �     p    @U
     �    PZ%          �`�          ��     �    @�     `    UP�     0    UU�         VU%         XU%         `U    �    �VU    �u     XU   `�     `U   XU     �UU   XU      VU  XU      XU  VU      `UU  VU      �UU VU       VU@VU       XUUPV�       `UUZV�       �UUUVe        VUUVe        XUUVY        `UU��        �VUV�         jUZ�         �V�z         ���~         ���_          ���          ���8         ��         � _=          �U�          CT          L                      �                                                          �           �                        �            0                       �                        @           pU           ��            p            �                                                   �            `            0                                               �           �u           `�           XU           XU           XU           VU           VU           VU          @VU  @      PV�  @U     TV�   X     UVe T`    @UVe@UU�U   TUUVY���UUPUUUU��PUUUUUUUUUUV����UUUUUUUUZ�PUUUUUUUUUU�z���UUUUUUU��~@UUUUU������_ �UU���������  ��     ���8         ��         � _=          �U�          CT          L�           3          �                                                          �           �                        �           �?           �
                                    @           pU           ��            p            �                                                   �            `            0                                               �           �u           `�           XU           XU           XU           VU           VU           VU          @VU  @      PV�  @U     TV�   X     UVe T`    @UVe@UU�U   TUUVY���UUPUUUU��PUUUUUUUUUUV����UUUUUUUUZ�PUUUUUUUUUU�z���UUUUUUU��~@UUUUU������_ �UU���������  ��     ���     ����       ����*      ������     ������*    ��������   ��������*  ���������" ����������� ����������*����������*���������������������� ���������������������� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������� �
       ���BUUUUUUU���@UUUUUUU( $��������������  �������������������������
  �TU�������������������������@U   �����������������������
     @�����������������������        ����������������������*        ����������������������
        ����������������������        ����������������������PU  TU  ���������������������*   U   P���������������������
��
  ��
���������������������
�������
�����������������������������*�����������������������������*���������������������� �������*��������������������� �������*P�����������������������������
  ���������*  ���������������J @U         U������*��������J   @UUUUUU P  ������*��������J              �������
��������
             ���������������*            ��������@���������            �������*���������B           ����������������
P       UU������   ���������� TU       ���  @U �����������*  @UUU�������RU  @��������������    �������     ������������������������*      ������������������������
     �������������������������
    P�������������������������    �������������������������  @U��������������������������TU   ��������������������������  ����������������������������������*  ����������������� �*UU����������������*PU   ����������������
     ���������������      @���������������       @��������������*        ��������������        ��������������RU  U @�������������� @U    ���������������� ������������������������B����������������������J����������������������J����������������������
���������������������
���������������������@  ���������
 �������� PU         @U��������   PUUUUUU  ��������              ��������B             ���������
            ���������*            ����������P           �����������T      @UU������������  UU       �������������
  PUUU������������������*    ������U���U����_�W��u��_���_���U���w�����������U�UUUUUUUUUUUUUUUUUuU�����_���U���w�����������U�U$UUUUUUUUUUUUUUWuUUU�_��_U�?�<sU�?��LU�?�<sU  �\U����_U��0\WU3<\WU�3 pWU�3pWU�3�_WU3\WU53�_WU�3|�_U���5pU?���pU0 0�pU? 0�|U 0�_U� ��WU��OWU??�W�?��W�?��W   @W�?���_���W����_UU�3 �W�� ?W� �  W�3���WU���U$UUUUUUUUUUUUUUWuUUU�_��_U�?�<sU�?��LU�?�<sU  �\U����_U��0\WU3<\WU�3 pWU�3pWU�3�_WU3\WU53�_WU�3|�_U���5pU?���pU0 0�pU? 0�|U 0�_U� ��WU��OWU??�W�?��W�?��W   @W�?���_���W����_UU���W���?W�   W�����WU����U(
           �    p  � �  `                  `�  @��  ��� ���0 ���p O>p �p��p�����>��������� ���� ���� ���� ���� ���p���p���0������  ���  ���  ���  �p  �                 @UUUUUWu�U�uUUUU]U��UUUUUUUU������u]����WWuUUUUUUUUUWu����UUWUUWWuUUUUUUUU��]w�uuUUUWU��UUUUUUUU]�UW�uuUUUWUUWUUUUUUUUUU��UW�]uUUUWU�_UuUUUUUUUU]�UW�UuuUUWU�w�_UUUUUUUU��UW����UUWUuW�UUUUUUUUUUWUW�UuUUUWU]W�UUUUUUUUUW�]�UuUUUWUUW�UUUUUUUUU��uu�UuUUUWUUW�UUUUUUUUUUW]��UuUUUWuU���UUUUUUUUUWW��UuU����UWUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUWUUUWUU�UUUUU]UU}U�������UUWuU�Uu��Uu]UUUU�UUWU��������u]W]UuuUUUu����_UUWUUuUUu]�_U]uU�����UW]UUWUUuUWuWW]U]�UUUU����_UUWUU��_u]�_UWUWUU]��UW]���U_UWuuWu�UW�������_UUUU���Wuu_]}UWu�U]�UuwUU�UUu]UWuuwWU�UU�U]�U]�UuW_UU��W�]�UUuUU�U]��WW_uW]uU]UWuWWWU]uU��_�}UW�uWU�U]UWuUw�UW�U�U��UUWU]WU�U]uWuU_u���WUUUwUUWUU��WUW�UuUWUUWUWUUU]UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUuuU�����u�UUUUUUUUUUUU���_]U]����uUUUUUUUUUUUUUuuU]U]��u�uUUUUUUUUUUUUU�U��������UUUUUUUUUUUU����]U]��UuuUUUUUUUUUUUUUUUU��]���]_UUUUUUUUUUUUU��W��]��uUUUUUUUUUUUUUUUWWW��]��W�UUUUUUUUUUUUUU��W��u�����UUUUUUUUUUUUUWWW]U���U�UUUUUUUUUUUUUU��W��u��U�uUUUUUUUUUUUUU]�U]U]�����UUUUUUUUUUUUUWUW�����u��UUUUUUUUUUUU�UU_]UU��U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUuuuU�UUUUWUUUUUUUUUUUUU����UUWuUUWuUUUUUUUUUUUUUuuU��������UUUUUUUUUUUUU��_UWUWU�_UUUUUUUUUUUUUU�]WU]�UUuwUUUUUUUUUUUUU�}�UUu�UU]�UUUUUUUUUUUUU�]�UUuuUUWWWUUUUUUUUUUUUU�WU�]U�UW�UUUUUUUUUUUU�UU�UUWU}UWuUUUUUUUUUUUUu��uU�]UUUWUUUUUUUUUUUUUU]�UUu�UUUUUUUUUUUUUUUUUU_W_U]UW��u]UUUUUUUUUUUU�UW]�WU���uuUUUUUUUUUUUUUUWU}UUuu�uuUUUUUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              $U��WUUU��_UUU��UUU���UU����UUU3��UU����WU�3WU�_UU 3_U�?  \U�� �WU��WU��?WUU��_U���WU5 <�UU < WU ��UU���WU�< <WU <_U  |U�   �W5   <�= �������0�U5�W?�U5�||U� s�_U� pUUUU�UU                        $UUUUUUUUUUUUU��WUUU��_UUU��UUU���UU����UUU3��UU����WU�3WU�_UU 3_U�?  \U�� �WU��WU��?WUU��_U����WU� <�UU5 < WU��UU<��WU0 <0 <p�0  |�  �����?�����0���  <0�U 0�U����                        $UU�UUUUU��uU]U���WU]U����UU�����sU533�pU���< \U�� 3 _U�0���UU�  �uUU� �uUu��uU��?�puU���3puUU5��uUU= ��UU� �UU�� �UU� �UU� �UU��}UU��UUU WU��WU���U� ���S3  3� ��   0��0��s�<?�p5   0\� W                            $UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUU��uU]U���WU]U����UU�����sU533�pU���< \U�� 3 _U�0���UU�  �uUU� �uUu��uU��?�puU���3puUU5��uUU= ��UU� �UU�� �UU� �UU� �U]��|u �� @0�0�0   �������<30p�00 _U���U                            $UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUU��uU]U���WU]U����UU�����sU533�pU���< \U�� 3 _U�0���UU�  �uUU� �uUu��uU��?�puU���3pu�  ��u3 ���_��    ��0��s�<?�p5   0\� W                            $UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUU��W]UUU��_]U����� ����3 ������    ��0��s�<?�p5   0\� W                            $U��_UUUU��UUUU���UUU����UUUU33sUUU����WUU�0WUU�<_UUU  \UU�?  \UU�� �WUU��WUU��?WUUU���_UU���_UU�0 �UUU�<��UUU���UU�0��_U50��UU5�?0|UU��?\UU=<0|UU���UU=  ��_U�� �UU� �  WU�����\U��p0\U5�s \U� p WUU�_��WU                            $UU��_UUU��UUU���UU����UUU33sUU����WU�0WU�<_UU  \U�?  \U�� �WU��WU��?WU���_� ��_�  �U= ? U���W5�0|U5� �U����UU� �UU 0|UU ��WU� UU5� �WU���|U5?�<�U=0��U�W�U= WpU��W�                        $U��_UUUU��UUUU���UUU����UUUU33sUUU����WUU�0WUU�<_UUU  \UU�?  \UU�� �WUU��WUU��?WUUU��_UU�0�_UU� �W�_�0 �U=��0 �W_5��|�W= <��U �|�W= ��\_5  �_=��  W�_u �_UUU��_UUUU�WUU����\UU��0\UU5�� \UU� � _UUU���WUU                            $U��WUUUU��_UUUU��UUUU���UUU����UUUU33sUUU����WUU�0WUU�<_UUU  \UU�?  \UU�� �WUU��WUU��?WUUU��_UUU��WUUU�UUUU�?UUU �pUU� 0pUU�� <pUU� ?�_UU� �WUU�   _UU�   |UU����_UUU� \UUU5��WUUU=<�\UUU \UUU= _UUU���WUU                            $U��WUUUU��_UUUU��UUUU���UUU����UUUU33sUUU����WUU�0WUU�<_UUU  \UU�?  \UU�� �WUU��WUU��?WUUU��_UU���WUU� �UUU� <�UUU� �WUU�� <WUU5��_UU5 <\UU= <\UU5 ��WUU=  �\UU��� _UUU��WUU��_�|UU��\�UU5 \�UU� _�UU��U�UU                            $U��WUUUU��_UUUU��UUUU���UUU����UUUU33sUUU����WUU�0WUU�<_UUU  \UU�?  \UU�� �WUU��WUU��?WUUU��_UUU��_UUU �UUUU0WUU�3�<WUU�0�<_UU�0��\UU����WUU��� \UU=�\UU� �|UU�?��UU��WWUU5�U�UU=�W?WU<W WU= W�WU��U��UU                            $UU��UUUUU��WUuUU��_UuU���?W�U���?_�U�����U��?� pU��� |U�� ��WU� ��UU�  �U��? ��U������UU�����U�<���U ����U? ���U��<�W� < W? ��W� �s�UU  |�UU  ��U�  ��U�?  ��UU�����UU�p]UU�5sU�s��pU� � pU�p� |UU�_U�_U                            $U��WUUUU��_uUWU��uUWU�����_������\U33s?\����7 W�0��W�<_UU  _]U�?  \]U�� �W]U��W]U��?W]UU��_]U����]U�0 ��_U�< �pU����pU����pU�� �_U5�� _]U5�? \]U50� |]U=�� \]U����_]UUU\]UU���WUUU���\UUU5�\UUU� WUUUU��WUU                            $U��W]uUU��_]uUU���UU���p�U������UU333 �U�����U�0�_U�<_WUU  _WU�?  \WU�� �WWU��WWU��?WWUU��_WU����WU�  3_U�  �0\U�  �\U�   �\U5  �WU5 ���WU5 ���WU=  �|WU�� _WU����pUU� \�WU5�_<\U��\=�\U0\�\U W� _U��UU�WU                            HUUUUUUU�U]UUUUUUUUUUUUUUUUUU��W]UUUUUUUUUUUUUUUUU���?_UUUUUUUUUUUUUUUUU���?WUUUUUUUUUUUUUUUUUU��?WUUUUUUUUUUUUUUUUUU��?WUu]UUUUUUUUUUUUUUU   TU�}UUUUUUUUUUUUUUU��?WU��UUUUUUUUUUUUUU�00WU�UUUUUUUUUUUUUU��WU5�WUUUUUUUUUUUUU�� �_5�UUUUUUUUUUUUUU��\� �UUUUUUUUUUUUUU���\?  WUUUUUUUUUUUUU�� �\ 0|UUUUUUUUUUUUU��7\ <�UUUUUUUUUUUUU�_�  �UUUUUUUUUUU���_5p   pUUUUUUUUUUU���?p   �UUUUUUUUUUU 0p  �UUUUUUUUUUU� 0 ��UUUUUUUUUUU� ��  ��_UUUUUUUUU�? ������UUWUUUUUU�?@�������UUWUUUUUU����� _U���s�_UUUUUU����� WU�����\UUUUUU������  WU����?\UUUUU�   �  WU?�3 WUUUU���? �?  \U?<��WUUUU���� �  \U?�|UUUUU=   ��   \U=  |]UUUUU   0?   |U�  p]UUUU��    �  p]��_]U�UU��      p��<\]U�_U3?  ���  p�?�\]Uw��300  ��?   �����]Uw��0�      ��7 <��]Uuw7 �   ���7 <��_UUw �   ����7���pUUu      �� �7���pUUU=     ���7� <�pUUU5  �  �� ��� <_U���  �  ��?0��� ���� � < �?<���  ����? �� 0�=�  <�|3  ��03?�? 0�� ��\3  �?0����00�0��?�\3 ��<���  ���� � ��\3������?  <? <0��3�\3��������� <00�\30�?�  �����0� �\30��<�  �? ���� ��\3<���0  �� ��������\3<���0  �����    �\3� ��0 ������?  ����3�0��< 0���3< �  �3���� 0  3< �����3�  0���3 ����3   0����� ��WUU3    ����� ��UUU��?���  ���� �?�uUU����    �?� ���UU ��������������?�uUU�������������� �_�UU���           ����uUU��������������������UU�����������������W�uUUU�����������������]UUU�����������������U�UUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUU��_UUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUU����_UUUUUU$UUUUu}UUU}UU�UUU�U�WUUUu��?��U�_5���UuU� �_Uu=� �UU�� U�    �U�    |UU    _UU=??�UUU����WUU����<\UU  ��WUU��UUUu���_UUUU���WUU�W���_]U]���W}U����_�W����W�W]�� _�_���  �U��< �UU�<_U�UU���s��U����_U�}������u���������������������������_�_U��W}U�WUU�wUUUUU��_UU$U}UUu}UUU�UU�UUU�U�WUUUu��?��U�_5���UuU� �_Uu=� �UU�� U�    �U�    |UU    _UU=??�UUU����WUU����<\UU  ��WUU��UUUu���_UUUU���WUU�W���_UU]���W�U����_�W�����U_]���_�_��<  UU�<�_�UU���WU�UU���wU�UU���_U�UU�?���UU������UU�����UU�����UU5����_UU���U�UU���]UUUu��WUU$UUUUu}UUU}UU�UUU�U�WUUUu��?��U�_5���UuU� �_Uu=� �UU�� U�    �U�    |UU    _UU=??�UUU����WUU����<\UU  ��WUU��UUUu���_UUUU���WUU�_���_]U}����W}UU�?� _�W��� |�W=��  _�_��< �U��?���UU���_U�U����s��}����_U�u������������������������7���������_�_U��W}U�WUU�wUUUUU��_UU$UUUUu}UUU}UU�UUU�U�WUUUu��?��U�_5���UuU� �_Uu=� �UU�� U�    �U�    |UU    _UU=??�UUU����WUU����<\UU  ��WUU��UUUu���_UUUU���WUU�W���_]U_���W}U��?��_�W����W�W]�� _�_��<  �U��< �UU�<_��UU���s��UU���_U�UU���U�UU������UU�����UU����?UU�����_U���W}UU��U�wUU�����UU$U}UUu}UUU�UU�UUU�U�WUUUu�����U�_5���UuU� �_Uu=� �UU�� U�   ��U�   0|UU    _UU=??�UUU����WUU����<\UU  ��WUU��UUUu���_UUUU���WUUUU���_]UUU=��}UUU� ��WU�<  ��W��< ��_U�<�|U�����_�uw���U�u_������UU���U�UU����W�U��3����U������UU?���UU�����_UU���W}UUu��wUUU����_UU$UUUU�WUUU�UU�WUUU]��UUUUW?�s]_U�U<��_UWU?  �UU����_UU=�0 ��WU�    _U=    �WU�    �UU���3 \�UU???�|�U����W�   �|�W�����W�WUw���UU_UU�?U�_�U���U�_�W��_U�W5 ���� ��U��� �U��� ��W��U��?���}u������U�������U�������U�??��U�����UUU������U�����WUUU���WU��wUU�UU��UUUU]UUU�WU$UUUUUUu}UUUUUUU_U�UUUUUU�W�WUUUUUUu�����UUUU�_5����UUUUuU� �_UUUUu=� �UUUUU�� UUUU�   ��UUUU�   0|�UUUU    _�WUUU=??�UUWUUU����W�_UUU����<\UUUU  ��WU_UUU��U�UUUu���_UU�UUUU���WU�?UUUU��_UU��UUUU���UU��UUU���WU��WU�� ��_U����� ��WU�����? ���������������}UUU������?]UUUU������}UUU��?���UUUU������WUUUU=���_UUUUUU�<_���WUUUU���UUUUU��UU�_UUUUU��UU�]UUUU?�uUU�_UUUU��UU�W$UUUUu}UUU}UU�UUU�U�WUUUu��?��U�_5���UuU� �_Uu=� �UU�� U�   ��U�   0|UU    _UU=??�UUU����WUU����<\UU  ��WUU��UUUu���_UUUU���WUUUU���_]UUU���}UUU��_�WU���|�W���� p�_u�� �Uu��3���}��U��]�������u�?�U�UU����W�U��3����U������UU���UU�����_UU���W}UUu�_�wUUU����_UU$UUUU��UUU�UU��UUUUW��_UUU����\�WU� |�W�U� �U�����WUU? <�UU3    �WU   ��UU=    |UU��� WUU���<_UU5�pUU5   ?_UU�?<��UUU�]?�UUUU���_�W�_����W}�� �_U_U�� U���? �U}}��  U�U��<��W=}W����U�uU����w��������������_�����?�������UU�������W��?����U�U�U���U_UUUU�UUUUUU�_UUUUUU�WU$UUUUu}UUU}UU�UUU�U�WUUUu��?��U�_5���UuU� �_Uu=� �UU�� U�   ��U�   0|UU    _UU=??�UUU����WUU����<\UU  ��WUU��UU�u���_UU�U���WUU�W���_UU�=��]U��?� _}U��� |�U]�<  p�WU�< ��_U�����_UU���UUU������UU���U?UU��<���UU��?���UU��?��|UU�<��U������WU����UUUU�_��UUUU����_UUUUU�ZUUUUUUUUUUUU��U�VUUUUUUUU�* �V%ZUUUUUUUU
   j
�UUUUUUU��
 `�UUUUUUU���� �"VUUUUUU
� � 
(�UUUUUU   
 � ��ZeUUU    
  �

�R	( �
� �  � �	 (    "*��`)( 

��*   
Z�� � �ijUU%�
 ��
�
 Z�UUU� ��*����VUUUU�
   � `
�eUUUUU)   �
h��UUUUUU�
 (Z�ZUUUUUUUUU)��VUUUUUUUUUUU�ZUUUUUUUUUUU	UUUUUUUUUU��VUUUUUU� jUUUUUU
 ��UUUU�   �VUeU	���UUU
   �jZU   ��� �� `U�� �ZU
 � `UU*(�
� XVU%  �* ZUU��
* �fUU��  hUUUU
  �ZUUUU)�*�UUUUU�j�jUUUUU�ZUUUUUUUUUUUUUUUUUU��ZUUUUUUUUUUUU* hiUUUUUUUUUU� ��VUUUUUUUU��  �ZUUUUUUUU)�    �UUUUUUUU     �VUUUUUUU
 ��*  ZUUUUUUU	�* �  ���VUUUU�(  �  * �UUU�
   �    �jUU)       *  �jU	 ( �   ��
 �� �
�� �V��jU  � �( �UUUZU	� �   �
hUUUUU�      V�ZUUUUU�*    �VUUUUUUUU� �
��UUUUUUUUU���jUUUUUUUUUUU�VUYUUUUUUUUUUUUUU��VUUUUUUUUUUU�� �VUUUUUUU�jU
  �VUUUUUU��� �� hUUUUUU�   � * �iUUUUU) �   � ���VUUU	��
 ���ZUU�
�  ��� � ��j	 �  ���    ��	�* �* ��(  ���  ( ���*   �"    � �� ��
   ��� � �j*��
   
�* ( �U�jU) �    ��
�UUUU�
�    hU�VUUUUU��   ZUUUUUUUUUU
 ��VUUUUUUUUUU��jUUUUUUUUUUUUUUUUUUUUUUU.
UUUUUUUUUUUUUUUUU�UUUUUUUU=�U��������W�        _�       �_�������WU������UU�����_UU�      |UU�      �UU�      �UU� �� UU� �� _UU� �� _UU� �� _UU� �� _UU� | _UU� |  _UU�    _UU� �_  _UU� �W�� _UU� �U�� _UU� _UU� _UU� ���� _UU�      _UU�      _UU� ���� _UU�������_UU��WUU��WUU��UUU��UUUUUUUUUUUUUUUUUUUUUUU�U}�UUUUUU�W_�UUUUUU��W�UUUUUU��U�UUUUUU��U�UUUUUU�U�UUUUUUU�U�UUUUUU��W�UUUUUU��W�UUUUUU��_�UUUUUUu�_�UUUUUU}��UUUUUU_���UUU.
UUUUUU�WUUUUU���_UUU���� |UUU5�� � |UUU5��< �UU� _<�?�UU� �   �WU�    �WUU  �?�UUU��  �WUU��   �WUU��    �W����  ��U��� ���U�  0��0�U�  <�  �W��<�   �WU�<0   �WUU<0�?��UUU0�?�UUU<�7�UUUU 0�7�UUUU  �?�UUUU   �UUU�� �UU� ��? ��U�       �W� �    �W�    �WU�_��   �UU�W�����UU�UU����_UUUUUUUUUUU��U_��UWU�U_���UWU�WW��UWU�����UWU�����UWU�����UWU�����UWU����UWU����UWU����UWU�U��UWU�U��U��UU�U�U�U.
UUUUUUUUUUUUUUUUUUUUU��UUUUUUUU5�_UUU�_UU5 ����|UU� 0    �UU�0    �UUU�    �UUU�����UUU=_���|UUU�_UUU|UUU_UUU|U��|UUU|U�  p���|U�  |   |U��|   |UU�|��UU}|���UUU||U�_UUU||U�WUUU�|UUUUUU |U�UUU |U��UUU�|U��UUU�|U��WU��|U��_U� |��? _U� |    _U� _   �_U��_   �WUU�W�����UUU�U����_UUUUUUUUUUUUUUU��UUUUUUU��UUUUUUU��UUUUUUU��UUUUUUU��UUUUUUU��UUUUUUU��UUUUUUU��UUUUUUu��UUUUUUu��UUUUUUu��UUUUUUu��UUUUUU��UUU������?��?�����������?�����������?��? �����  ?�? �����  ?�? �����  ?��������������������������������� �����?�  ?� ���� �  ?� ���� �  ?������� ��??������� ��??������ ��??�?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����??  ?��� ����??  ?����������?  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��UUU��WUU�5 |UU�- �W�  ��� ��*�_������W������UU����WUU���UUUU=  _UUU� �UUՀ
 �WU5(  �^U
   ^U�  �zU  ���U   ��_   ���+   ����
 ����������������_������W������UU����_UU����UU
UU�Z�Z�V��jU)����������jU�ZZU�jUU��UUU�V
UUUiUU�jUU�j�Z�Z���V)�������U��jU�jZU�ZU^( ��*                                ��:   �                                 8 ����                                ���� 
�                                "(���(�                                "���("���������������������������������""���"�   �   �   �   �   �   � "����""�(��"�(��"�(��"�(��"�(��"�(��"�("����"� ""� ""� ""� ""� ""� ""� � ����"�*��"�*��"�*��"�*��"�*��"�*��"�*����                        ���������������������������������������� ���������������������������������?��   ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��    "�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU"�    �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU"�    ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��    �UUUUUUUUUUUUUUUUU�WUUUUUUUUUUUU"�    "�UUUUUUUU�UUUU���_UUUUUUUUUUUU"�    ��UUUUUUUU=�UU���� |UUU��UUUUUUU��    �U��������WU5�� � |UUU5�_UUU�_U�    ��U�        _U5��< �UU5 ����|U��    �U�       �_U� _<�?�UU� 0    �U�    ��U�������WU� �   �WU�0    �U��    "�UU������UU�    �WUU�    �U"�    "�UU�����_UUU  �?�UUU�����U�    ��UU�      |UUU��  �WUU=_���|U��    "�UU�      �UUU��   �WUU�_UUU|U�    "�UU�      �UUU��    �WUU_UUU|U"�    ��UU� �� U����  ��U��|UUU|U��    �UU� �� _U��� ���U�  p���|U�    ��UU� �� _U�  0��0�U�  |   |U��    �UU� �� _U�  <�  �W��|   |U�    ��UU� �� _U��<�   �WU�|��U��    "�UU� | _UU�<0   �WU}|���U"�    �UU� |  _UUU<0�?��UUU||U�_U"�    ��UU�    _UUU0�?�UUU||U�WU��    �UU� �_  _UUU<�7�UUUU�|UUUU"�    "�UU� �W�� _UUU 0�7�UUUU |U�U"�    ��UU� �U�� _UUU  �?�UUUU |U��U��    �UU� _UU� _UUU   �UUUU�|U��U�    ��UU� ���� _UU�� �UUUU�|U��W��    �UU�      _U� ��? ��UU��|U��_�    ��UU�      _U�       �WU� |��? _��    "�UU� ���� _U� �    �WU� |    _"�    "�UU�������_U�    �WU� _   �_�    ��UU��WUU��WUU�_��   �UU��_   �W��    "�UU��UUU��UUU�W�����UUU�W�����U�    "�UUUUUUUUUU�UU����_UUU�U����_U"�    ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��    �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�    ��UUUUUU�U�W�_����_U����W}UUUUU��    �UUUUUU����_��_��_U�U�W}UUUUU�    ��UUUUUU��W�_��_��U�U�_]UUUUU��    "�UUUUUU��W��_��_���U�U�__UUUUU"�    �UUUUUU��W��_��_���W�U�WUUUUU"�    ��UUUUUU��W��_�����_����WUUUUU��    �UUUUUU��W��_��_��_�U��WUUUUU"�    "�UUUUUU��W��_��_����UU�UUUUUU"�    ��UUUUUU��W��_��_�����UU�UUUUUU��    �UUUUUU��W��_��_��U��UU�UUUUUU�    ��UUUUUU��W�_��_��U��UU�UUUUUU��    �UUUUUU�_��_�u�_��U��UU�UUUUUU�    ��UUUUUU�WU�WU�_�_��U����W�UUUUUU��    "�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU"�    "�U�����UU����W���U�_�U���U�W���    ��UU�U��_UU�W�W��_UU�_�U�U�U_�U��    "�UU�U��_UU�W�W��_UU�_�W�U�U}�U�    "�UU�U��UU�W�W��_UU����U�W]�U"�    ��UU�U��UU�W�W��_UU����U�U�U��    �UU�U��UU�W�����_U�������W�U�    ��UU�U��UU�W�W��_UUU���U��_�U��    �UU�U��UU�W�W��_UUU����UU��U�    ��UU�U��UU�W�W��_UUU���U���U��    "�UU�U��UU�W�W��_UUU���U�U�U"�    �UU�U��_UU�W�W��_UUU���U�U�U"�    ��UU�U��WUU�W�W��_UUU���U�W_�U��    �UU�U��UUU�W�W����UU��_���W�W�U"�    "�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU"�    ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��                                     �  ��������������������������������������� �                        ����"�*��"�*��"�*��"�*��"�*��"�*��"�*�����"� ""� ""� ""� ""� ""� ""� � ���""�(��"�(��"�(��"�(��"�(��"�(��"�("����"�   �   �   �   �   �   � "���("���������������������������������""���(���������������������������������"��� 
�                                "(�����                                ���  �                                 � ���                                ��:  ��?                                ��? U�UU�UU�UU�UU�UU�UU�UU�U��W5W?3_33_33\33_�W W�U=�U5�U5�U�U	�_=�_�W�U�W_=��_
p � ��r���  �� �@ p /�@� �@� D@L�LB@ %S! ����@�BL�@Q$@$@���B$S�B  �@�`tBp�,�(                                                                ����@ @��@��@��B������@@��@$@""�@/r�@ �@@  @`�������@O��� ��
U��UU�_U�
`�)��%��*��*8����%�����j�U�VU
U��UU�_U�*`�)��%��
��*�����%����j�U�WU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �(UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@                                        @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @                                                                                                                                                                                                                                                                                                                                                                                                                            ��                                    

 *                                   �� �                                   �   ��                                �   � 
                                �                                       (  �� (                             ���
 � �                            �* *  �   �*                            �   �*   (�                          �  *       
                        �� �
�  �
 
                           ��
� � �(�                            �  � �* �*                                 
�(  ��                               �      �
                                �     �                                 ��� �                                   ��
�                                     �*                                                           ��
                                    
�
(                                   �  �                                   (  *�                                 �
 ��
                                 ��                                 �  
�
((                                   ��                                �  ��                                 ���                               �

�   �                                ���   �                                  *���                                  ��   
                                   * �                                     � 
                                     ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �
                                     ���                                  ���� �
                               �����   �                               �" �   �
                              
 **(���                             ��
�
* �
                            ��� � � * ((                          �  �� ���� ��                          (*�"   �� ��                         �   ( ��*� ��                          
���  � ��                               ��
 ( �                                 ��� 
 �                               "* �(
�                                " ��
                                 ��  �                                   
 ��                                    � *                                     ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �(UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� XUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% hZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% �bUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�  �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU
 �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� �*�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� ���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�  � VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� (� ZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU� XUUUUUUUUUUUUUUUUUU
�hUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU

 `QQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQQ	( `U
�  DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD� `�  @@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@  `�  (                                  
 �
@ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @ @   �                                    ((                                                                         
        �*                         (�        (�                    ��*  � �       �
                   ����  
 �        �                    ����*            (�                 �_ZZ��  " (        
                 ����]�  
       �
                   n_Z_��
 ��       �� ��                �����U�
� �        �� ��                �_��o��+���        �����                �����f_/��"        �"��                �������� "         "��                ������o� 
"         ���                ��@�����
(�         �                  � P� �         �      �
             ����+��        � �    *(             仾~/��        � �   �            #����/��        �  
   � �           |���~/��        �
     �          WU���/�          
�
  �* 
          P�S�~/ (          *  ���          0 �P��/ (         ( �    � (          0<<���/  �       ��      �          0� ��+ ��       � �   (( �          0   �� 
*        �     �(             �� �         
     �             @��
("         �    (��            @ ��(*�        �   
���            @ ���
(*    
   �    �  �            @ ��
�   ��   �    � (�          |  @���
�    (�    
  �
�          �
 @���+��    �      (��          �� @���/��    (
        (              + @���? �    �           (            P}}�> �� ��
      (� 
            TUV徠�  �  (      �
            p uP����  �  �        
(�           �U]@�ꂀ� � � �       �*               �W @�ꋀ(� ����       �  �            p @�ꏂ�* �� �       ��"            � @��/�  �� 
�        (              @���   �                         @���*  
� (         �� (              ����*�    ((       � �
            �  Ъ����   
       �
 (            `  䪪��  �(        ( �            0  y����  �          * (               m���
*�  �         ��              @o���              �               �k���   
   �       � 
            � ey���*
 (� (       �             �uUzy���
 �  �       �             `ի^^n�� �   

       ��"            XU�W^n��         �
             XUU�Wk��� (         (            XUU�����+*� � 
        ��            VUU֖ۺ� � �  �        ��             VU��eۺ� � �  (         ��             VU���ں�              `�            @VU��ٺ��    
 "         ��    @      PV�ezٶ��("  (           �   @U     TV��^����� "  ��          `      X     UVe�W������   � �         ��   T`    @UVe�������
(  ���         ��  @UU�U   TUUVY������   ��         �  ���UUPUUUU��~e����   "           (  PUUUUUUUUUUV�_�j�����   "(          �  ���UUUUUUUUZ�W�ں����  � 
            PUUUUUUUUUU�z��������   �           (  ���UUUUUUU��~֫����   ��           �  @UUUUU������_�j�*  �   ��           �   �UU����������ڪ  (
   ��           "    ��     �����* �
�  ��           *            �V���*�   (*   �                       TU���
  � �   
                    @UUU����
� 
    
       ���         �VUU�����
             ( ��     ��ZZ�������* � �         �
  �*    ��ZU�����������*�    (      � �  �  ��j�W��������꿀  ��(          * �
 �� �����Uկ�������*� ��    
     �  �
 ������_�U��������
� �     
     (    (  �����V���������+ �
*    �     
    �  ������u鯪����ꪢ�    �     �   �� 
 ������������+說+  �
   �     �  � �( (<���������� �
 �   �        (  
������������<�  �� �            
  ( 
0 ��� ���/� �� �    �     �  �   ( 0��/ ����   
�* �
         �  � � ����  0��2�*   ���          
 
 � � < ��2 ���  � �
��          (   0 � ���5 �/  � �� ��            (� 
�U0/p� �� � �  
      �*  � �*  pU0.\U�� � �*         �
�*  
   �\U5�� WU02�) ���
��  ��   �*�   
WU����UU502p�*(  ��� �  �
 �* � 
 �� WU� 3�UU5�pU�  (
 �*  
   
� �   ��UUU3pUU��\U% �
��  ��
  
 (�*  ��UUU3pUU��\U)�   (j)  � (��  
( (�   ��UUU3pUU��\U	  � ��� �   �
* �����WU�3�UU��|U	� 
 � �  
  
(���� 
� WU� 3�UU5�pU	   * � � � � *��
� |U= 3 _U��W) � �   �
 � �
 � �"����� �� 00 ����*�     �  �  ��*�   ��   <�  ��  ��( ��    
*��� �  ��<   <   �� �*� �����   ��*�(* ��� ��   Of<  ��  
� �(  �  �  � ��*��? ���� �hf��+   � �  ��
 �  � ( ��*����f���?��������� �  �*( �   �  ���������ff��������     �  
� ��* (   jff ���Y  �j& 
�*     ���� 
   ����(XUUUUUUUUUUU�*   �       

 ��� �
  �����W�����w�- � �       (( �� � j�:�p� 7�p� ' � ��        � ��������01L��01L�� �           ��
(�� �p<O�S�T<O�S�T<	�            �   * � �Aj���Aj���A*   ��
        
   �
�*�����������������*   (�        � ��   �����������������    IUUUUUUUUWuUUUUUUUUUUUUUUUUUUU�_�uUUUUUUUUUUUUUUUUUU�?�|UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\U�uUUUUUUUUUUUUUUU  PU��UUUUUUUUUUUUUUU���\U5�WUUUUUUUUUUUUUU��0\U5�WUUUUUUUUUUUUUU3<\U��_UUUUUUUUUUUUUU�3 p���UUUUUUUUUUUUUU�3ps��WUUUUUUUUUUUUU�3�_s�  \UUUUUUUUUUUUU3�s= ��UUUUUUUUUUUUU53��p= ��WUUUUUUUUUUUU�3|��=   �UUUUUUUUUUUU����=   �UUUUUUUUUUUU?����=   �WUUUUUUUUUUU0 0��=0   WUUUUUUUUUU�? 0��=0  WUUUUUUUUUU�? 0�_?0  ��UUUUUUUUU�� ���?�? ��UU]UUUUUU�?� � �����wU]UUUUUU�?���� |U����UUUUUUU�?���� \U�����sUUUUUU�?���� \U133�pUUUUU�   � \U���< \UUUUU�?� ��  pU�� 3 _UUUU��3 �  pU�0���UUUUU�   ��   pU�  �uUUUUU=   0��   �U� �uUUUUU�  <    �u��uU�WU�      ���?�puU�U��0  <33  ����3puU��W���  ���    _��uU����<�     � � ���wU��� ?   ��?0 � � ?UU�=  0   ���3 � 0�UU�5   0   ��0 � ��UUU�   0   � � ���UUU�  �  �������}UUU�    �� �W �UUUU �  �<�0�W �zUUUU= <<3 ?< ���� 0�UUUU���� � �� �?0VUUU�?�������������00XUUU����� <�?�0`UU�����  �� 0�����`UU��?�?�  �? ���0<0`UU���<0?  �������?0 `UU�����  �  �0�`UU�����  ����� �`U�����  ����     XU	��?� 0������      XU����� �0����     �V� ��?�? �00  �     jU�   00 �0���<   ��UU%    00 �����<  �`UUU% � 0� ���<   �UUU%  � 0 ���<    VUU%   �?  ����?    XUU�   (   <��?    `UU�
  �00 �� �  �* �UUU)  �0? * 
�  � �UUU�  �  �   ���  `UUU�
 (     �     � XUUUU��             VUUUUU%           �& �UUUUUU�           j� ZUUUUUU���      ��UU�UUUUUUUUUU�    ��UUUUUUUUUUUUUUU��
 �VUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUIUUUUUUUUWuUUUUUUUUUUUUUUUUUUU�_�uUUUUUUUUUUUUUUUUUU�?�|UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\U�uUUUUUUUUUUUUUUU  PU��UUUUUUUUUUUUUUU���\U5�WUUUUUUUUUUUUUU��0\U5�WUUUUUUUUUUUUUU3<\U��_UUUUUUUUUUUUUU�3 p���UUUUUUUUUUUUUU�3ps��WUUUUUUUUUUUUU�3�_s�  \UUUUUUUUUUUUU3�s= ��UUUUUUUUUUUUU53��p= ��WUUUUUUUUUUUU�3|��=   �UUUUUUUUUUUU����=   �UUUUUUUUUUUU?����=   �WUUUUUUUUUUU0 0��=0   WUUUUUUUUUU�? 0��=0  WUUUUUUUUUU�? 0�_?0  ��UUUUUUUUU�� ���?�? ��UU]UUUUUU�?� � �����wU]UUUUUU�?���� |U����UUUUUUU�?���� \U�����sUUUUUU�?���� \U133�pUUUUU�   � \U���< \UUUUU�?� ��  pU�� 3 _UUUU��3 �  pU�0���UUUUU�   ��   pU�  �uUUUUU=   0��   pU� �uUUUUU�  <    �u��uUUUU�      ���?�puUUUU��0  <33  ����3puUUUU��� ����    W��uUUU��<�0   � � ���wUUU� ?�0 ��?0 � � ?UUU5  0 ���3 � 0�UUU5   0? ��0�� ��UUU�   0�   ��� ?���UUU�  � �����?��}UUU�  �3  �� 0�� �UUUU ��� �<�00 � �zUUUU= <�  ?< �0 �  0�UUUU�0 � � �0 ? �?0VUUU�?�< �����0����00XUUU���  <�?�0`UU�����  �� 0����`UU��?��� �? ?�0<0`UU���?0< ������?0 `UU���?� � <�0�`UU�����  ������ � �`U���� ����?�?      XU	���?  0��?��      XU���?  00����     �V� ���� 00� ��      jU� ���?< 0���   ��UU% 0 �� �0��?   �`UUU% � <�* �����    �UUU% ��̯  0���?    VUU% � 0
  0�?�     XUU� �3�   0���     `UU�
 ���  ��2�3  �* �UUU)  �   * ���  � �UUU�  �  �   < ?   `UUU�
 (     �     � XUUUU��             VUUUUU%           �& �UUUUUU�           j� ZUUUUUU���      ��UU�UUUUUUUUUU�    ��UUUUUUUUUUUUUUU��
 �VUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUIUUUUUUUWuUUUUUUUUUUUUUUUUUUU�_�uUUUUUUUUUUUUUUUUUU�?�|UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU  PUU]WUUUUUUUUUUUUUU���\UU_UUUUUUUUUUUUUU��0\UU�UUUUUUUUUUUUUU3<\UUUUUUUUUUUUUUUU�3 pUU�UUUUUUUUUUUUUU�3pUU�_UUUUUUUUUUUUU�3�_UU? |UUUUUUUUUUUUU30PU� �UUUUUUUUUUUUU53�_U� _UUUUUUUUUUUU�3WU� |UUUUUUUUUUUU���UU�  �_UUUUUUUUUUU��UU�   \UUUUUUUUUUU� �UU� �|UUUUUUUUUUU� �WU�  pUUUUUUUUUUU� �_�� 0pUUUUUUUUUUU� ��5� ���UUUUUUUUUU�� ?�<����WUUUUUUUUU �� � ���_UUUUUUUUU��� �� �W=��UU]UUUUU���?< pU���uU]UUUUU���? pU���|�UUUUU�?   0 pU��?���sUUUU=����� �U����pUUUU�?� 0�  �U�� � \UUU�  ��?   �U� �5 WUUU�     �  �W�  ��UUUU�  � <   ��? �U]UUU�?<    0   �����U]UUU5��  ���<   W����U]UUU=���   \<��WWUUU� ��  �� \���_WUUU00��  ��\���WUU�  <�����??� <�WUU�   ��  ��? � < WUU�  ��0 � �� � ��[UUU �?�0 ��?� �����`UUU  �0 ��� � �?�UUU= �3�0 ���  �0 VUU� ���0 �� � � �0 VUU��< ���� � <  �0 VUU���?�?���?� ����0 VU��?��? ��?�3 �0  VU����� �� 3 �??  VU���3���3 �� ����UU��������?   �UU��?��?�� �    �UU��?� ����  �����UU>���� �����       `U������� �����       XU% ����� ���      XU	 ���?�  �   � VU	   � ���?0    (�UU	  ? � ����    �jUU	 (�� ? 0�?���   VUU	 ����� �3���� � XUU	  � ?�  ��?    `UU	  ��  �    �UU%   
�3   ?�     �UU�   �    0 �    
  �UUU      ���    �  �UUU	            Z* hUUU�  �          �V� VUUUU
 
  �      �UU�UUUUU��   j	     �ZUUUUUUUUUU �V�*    hUUUUUUUUUUU	 �UU�����VUUUUUUUUUUU��ZUUUUUUUUUUUUUUU                                    �(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      PUUU                                   T                                    U   TU                                T      PUUU                                                                          TU                            P     @UU                              @     *                                 TUUUQU                                    T                                                                                                                                                                                       PUU                                    PU @U                                 TQ                                                                       @U     P@                              P    UU                            PU   @                              P     @   @            PU               U    @P            TUQ               UPU     P           TUUY                                 UUU]                                 UUU^                 @U@U@           UUUU                  @U PU            UUUU                                   UUUU                                   UUUU                                   UUUeU                                  @UUUi�                              @  @UUUi�                              PU @UUUj�                             PUQ@UUUj�6                             PUUUPUUUj�             
             jUVUQUUUi��           PUTi           �Z�UUQUUU��ZP          UUU�Z�          �ZUUUQUUU��Z           UUU�j�         �VUUUU              @UUU�j�         �VUUUVU%              @UUUej�         �VUU�VUU�
   @         @UUU�i�         �VUU�UUU��  @         PU�U�U�V         �VUU�UUUU�  P         PU�UeU�U        �VUU�UUUU�ZU          PU�U�U�U        �UUU�UUUU���U          PUiU�U�UU        �UUU�UUUUU��           PUYU�U�UU        �UUU�UUUUUY�           UUUU�U�UU        �UUU�UUUUUY�          �UUeUUU�UU       �UUU�UUUUUU�         PEUUUUUU�UU
       hUUUeUUUUUY�       @UTUUUUUV�UU*       hUUUiUUUUUU�      @   PUUUUVVUU*       hUUUiUUUUUU��    P     PUUU�VUU)       UUUUYUUUUUU��6           PU�ZUU)       UUUUYUUUUUU��5     PUU  @UU�ZUU)       UVUUZUUUUUU�b5      @ PUU�ZUU)      @�VUUZUUUUUU�ju      T UUU�ZUU)      @�VUUZUUUUUU�Zu    T  TUUU�ZUU)      @UUUUZYUUUUU�ZU   @   @UUUU�ZUU%      �UUUUZeUUUUU�VV      EUUUUU�ZUU�     �UUUUV�UUUUU�ZUU   PUU`UUUUU�ZUU�     �YUUUV�VUUUU�jUUU     �UUUUU�YUU�
     hUUUUi�jUUU���ZUU     �VUUUU�UUU�*    ��UUUU���UUU�����UU    �ZUUUUUUUU��
  ����UU����jU��������U��ZU��UUUUUU�������                     �������UU�����������(                  �                                      �                                 �    �
                                 �
   �)                                  ��  �%                                  ��
��                                   ��
��                                    �*��                                    ��`�                                     �z�  �*                                 Z~) |U�                                X}) W�                                 h})���                                  hu	�                                   �U\)                                   �U_
                                   �VUW                                   �Vu�                                    �Fe�                                    �Ee)                                    �E�
                                    ��
                                    ��                                    �U�                                     �U                                     �U                                     �V�                                     �VU                                     �VU                                     �ZU                                    �ZY                                    �Za                                    �VA             �                     �UQ            �*                      �UQ           ��        ��            `UQ          �j          �
           `UA         �jU            ��         `UQ        �jU              ��        hUQ    �*  ��V                ���
      XUQ   ���
�jU                T���      XUQ   �U���V                  T��     UU  �ZU�j                   T�
     UU  �V�_UUUU                  @U�    @U  j  @UUUU                   @�    @U �Z    PUU                   �   @U �V      T                   �
   @E �U       @U                   \
   @A �U        T                  T)   @U j        @                  P�   @T�j         U                  @�  PUQ�f         P                  �
  PUU�f                             T�  TWU5�Y                             P�
 T�U�ZY                             @U� TUT�VV                              U�*XUT�UY                               T�*ZUPe�                               P��VUQUU                               @U�VpAUW                                U�U�E�_                                TUG��                                 TUED�?                                 P�AUT�       TUU                @UU  @uTT�      @  P               U    _PT�     TU    @             P  PU \PT�     @     @P            P      \AU     P                  @U      PAQ          U            P       PAQ     @ U               T     @  PAP      P    @           P  TU   PPT      PU                  U     @TT           T               TU    @EPT       @UUUU                      @TT                                   @T                                    UE                                    @A                                    TQP                                    Tu                                    TE                                    TA                                    PQ                                    PQ                                    TU      �*                            TU ���
���                           \UE �����
                             \QE�ZU���                              \QEjUUUU	                              WPU�VUUUUU                             WPU�UU @U                             _TUiU    U                             TUUU    PU                           TUU       U                          |UUU                                   4UUU                                   0TUU                                   pPUU                                   pUUU                                   pTU                                    pTU                                    pTU                                    @TT               *               �
   @QT             �       ��*      �*   @Q@            �
        ��
  ���Z�  @QUP            �         ����Z��U�   AUT           ��U          �jUUUUUU�  AUU           �VUUU         @U @U�
 @EUU           ZU                  @�
 @UU          �U                    U� @UU      � �Z                    T�@UU     ����U                    P�
@U    �����j                     P�
 U   �VUU��Z                     @U
 UUU   jUUUU�V                      U) UUU  �ZUU @U                       T�UUU  �UU   T                        T��UUU  �U                             T��UUu �[                             PU�UUU �V                             @U�UUU�kU                             @U�UUU�VU                             @U�UUUjUU                               UUUUU�ZU                               TUUQC�VU                    PU         TUU�P�U                   T          PUUPU                  T  @U       @UUUTU                 @  @UU        UUEU��                 @   T   TU      TUEuQ�                  @       @     TUEMQ�                    PU          @UEMQ�                   P     @      UUA�                    U    @       WQE�                     T  U        WQE}                     @U           WACu                       UU         WECQ5                                   WEOQ%                                   ]E}P                                   EuT                                   EUU                                   DTU                                   TPTU                                   TAUU     �
 @               �        UUU �  � P���       $UUUU_UUUUUUUUUUUUUUUU�pUUUUUUUUUUUUUUUU5�UUUUUUUUUUUUUUU��WUUUUUUUUUUUUUU  ��UUU�_UUUUU�����0�_U��UUUU? ��?��0�W�  �_UUU? ?����0��pUUU  �����0� �UUU ��� ����<<?WUU  � ?��?��\UU  <����\UU��<<??��UU?<� ?<<<� ��UU  � <<<0< ��UU� � 00���� WUW �  <<� �  ��WU�U��5� �   �WUUUU_5<     < �_UUUUU5   �? ��\UUUUU��?�� �0<pUUUUU����  �� �pUUUUU�?� ����3�UUUU��p��UUU�� ��UUUU�? \UUUUUU� �WUUU� WUUUUUU=0p\UUU �UUUUUUUpUUU?pUUUUUUU5p��UUU�\UUUUUUU�p��UUU�WUUUUUUU�pU�UU� �UUUUUUUU= \U}UU pUUUUUUU� WUUUUpUUUUUUU5 WUUUU� \UUUUUUU5�UUUUU� \UUUUUUU5pUUUUU��WUUUUUUU��_UUU$UUUU_UUUUUUUUUUUUUUUU�pUUUUUUUUUUUUUUUU5�UUUUUUUUUUUUUUU��WUUUUUUUUUUUUUU  ��UUU�_UUUUU�����0�_U��_UUUU? ��?��0�W�  �UUUU? ?����0��WUUU  �����0� \UUU ��� ����<<_UUU  �?��?��UUU�<<����sUUU�<<<?���UUU� � 0<< < �UUU  � 0<0<��UUU� ��0� � �UUUW _� � � �UUU�U��U�� 0   WUUUUU_U��    0�WUUUUUUU=�     pWUUUUUUU=���� \�_UUUUUUU�<� � W�_UUUUUUU��< �U�|UUUUUUUU�U0pUpUUUUUUUU\U=?\U=pUUUUUUUU�\U�\U5�UUUUUUUU5 \U�\U��WUUUUUUU� pU5 \U��\UUUUUUU� pU?WU�pUUUUUUUU3pU�WUUpUUUUUUUU=�U� WUU�UUUUUUU��� �UUU��WUUUUUU50� �UUUU�WUUUUUUp� pUUUU�UUUUUUU\� \UUUUUUUUUUUU��_��WUUUUUU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUU����UUUUUUUUU�� jUUUUUUUUU�*�VUUUUUUUU��hUUUUUUUU�
(�VUUUUUU����XUUUUUUUU�
 `UUUUUUUU� @UUUUUUUU*  �UUUUUUUU�
��UUUUUUUU��_UUUUUUUU���UUUUUUUUU��_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��jUUUUUUUUU��VUUUUUUU�� jUUUUUUUU���UUUUUUUU�  �VUUUUUUU  jUUUUUUUU% ��VUUUUUUU� 
��ZUUUUUUU
��jUUUUUUUU� 
XUUUUUUUUU
��UUUUUUUUU��jUUUUUUUUU� ��ZUUUUUUUU��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUU�jUUUUU�_UUUU�ZUUU���UUUU��VUU% �_UUU�
hUU% ��UUUU)�VU	 ��_UUU�
hU	����UUU���U	 �U�_UU� V	�jU��UUU* X%�jUU�_UU�`% �UU��UU�*`� �VUU�_U���U jUU��U��U	(�VUU���*�U��ZUUU��� �UU
�UUUU�/`UU��ZUUU�� `UUU*hUUUU�XUUU��VUUU��UUUUU�jUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUU�UUUUUUUUUU��WUUUUUUUUU%�WUUUUUUUUU%�_UUUUUUUUU	 _UUUUUUUUU	 UUUUUUUUU� |UUUUUUUUU� �UUUUUUUU�  �UUUUUUUU� ��WUUUUYUU���WUUUUYUU%���_UUUUYUU%��j_UUUUYUU%��YUUUUYUU	�fY}UUUUYUU��UU�UUUUiUU��UU�UUUUjUU��UU�WUUVjUU��UU�WUUVjUU��UU�_UU�bUU�UUUU_UU�bUUiUUUUUU�bUUeUUUU}e��`UUeUUUU�e��XUUeUUUU����XUUeUUUU���"XUUeUUUUՋ� VUUeUUUU��VUUUUUUUU VUUUUUUUU? �UUUUUUUUU= �UUUUUUUUU� `UUUUUUUUU� `UUUUUUUUU�XUUUUUUUUU�XUUUUUUUUU�VUUUUUUUUUU�UUUUUUUUUUU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU0UUUUUUUUUUUUUUUUUU�VUUUUUUUUU�hUUUUUUUUU% �UUUUUUUUU	  UUUUUUUUU _UUUUUUU�  _UUUUUUU� ��_UUUUUUU% ��WUUUUUUU%���WUUUUUUU	���UUUUUUUU����UUUUUUUU�h�~UUUUUUUU�Z�UUUUUUUUbZU_UUUUUUU�hV�_UUUUUUU�XV�WUUUUUUU�ZU�WUUUUUUU%VU�UUUUUUUU�UU�UUUUUUUU�UU}UUUUUUUUeUUUUUUUUUUeUU_UUUUUUUUUU�_UUUUUUUUUU�WUUUUUUUUUU�WUUUUUUUUUU�UUYUUUUUUUU�UUYUUUUUUUU}UUZUUUUUUUUUUZUUUUUUUU_U�XUUUUUUU�_U�VUUUUUUU�W�%VUUUUUUU�W�)VUUUUUUU�U��UUUUUUUU�V��UUUUUUUU�V)�UUUUUUUU�Z
bUUUUUUUU���`UUUUUUU���XUUUUUUU�� XUUUUUUU�� VUUUUUUU�   VUUUUUUU�  �UUUUUUUUU  `UUUUUUUUU XUUUUUUUUU)�VUUUUUUUUU�jUUUUUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �(UUUUUj������V�i��jUj�U�U�V�UZ�RUUUUUUUUUUUU�����Z��jiZ�U��ZU�VUUZeUV�PUUUUUUUUUUUj��e�V�U�UZi�U�ZU�U�UYe�V�  @UUUUUUUU���UeU�Rj���ZieU�V��V�U��j�(TU  UUUUUZZ�UYV�BZi��iYe��V����Z�U��
UUUEPUUUUXU�V�ZU
ZYe����j��)���jUj��BUUUTTUUUU�BUVfi�*i�Z���UU��* ��U�V��PUUUUTUTUUUUH@VYe�*dU�*�Vj�V�
UU��J  �*TUUUUPUPUUUUU HZ�Z���Zj �Z�Ve�@UU�j���UUUUUAUAUUUUU�J�V�B��Z�ZU�*TUUU�� *@UUUUTEUUUUU�
@���
U�Z�UeU�UUUUU   PUUUUPEUUUUU(
 P *(`UeU���PUUUUUUUUUUUTUUUQEUUUUUU�*��
��jJYeU�
TUUUU PUUUUUTUUUQUUUUUU ���*@��RIY�U�@UUUUU�BUUUUU TUUQUUUUUUA��
U�P	e�U�PUUU  �
  TUUUTUUQUUUUUPU �BUU�R)�j��BUUU�*����PUUUPUUQUUUUUPUU PUU�JTeJUU�
�*�RUUUQUUUUUUUUQUUTUUU*P���JUU�J!@U� RUUUAUUUUUUUUAQUUTUUU�U��@UU�@ UU�TTUU UUUUUUUQAUUTUUU*  �*TUU�X�UU�V�PUUEUTUUUUUPEUUUUUUE���� UUU�X�UU V�RUUEUUUUUUEUEUUUUUUEU�
�*TUUU�X�ZU jRUUEUTUUUUAUEUUUUUUEU@
UUUU�XhU�RUUEUUPUUUUUUAUUUUUUAUUU@UUUU!X`UA�
RUUEUU@UUUUUQUUTUUUQUUUUUUUUU ZUhUQ�
RUUEUUUEUUUUUPUUUTUUUQUUUUUUUUU(VUhUQ�RUUUUUEUUUUUTUUU@UUUQUUUUUUUU(VU�UQ�RUUUUUUUUUTUUUDUUUQUUUUUUUU�VU�UQ��RUUUUU TUUUUUUUUU@UUUUUUU�UUhUU��BUUUUUU@UUEUUUUUUUEUUUUUUU��UUhUU��
UUTUUUUUUUUUTUUEUUUUUUU�jUUhUU��*TUUPUUUUUUTUUUTTUUEUUUUUUU�ZUU�UU���TUUQUUUUUUUTUUUTTUUEPUUUUUU�ZUU�UU�PUUPUUPUUUUUUUTTUUEUAUUUUU�ZUU�UU�RUU@UUUQUUUUUUUUTUUEUEUUUUU�YUU�UU�VRUUUUUQUUUUUUUUTUUUEUUUUU�YUU�UU�jBUTUUQUUUUUUUTPUUTUUZiUU��YUU�UU`JUUPUUQUUUUUUUUTAUUUTUU�ZUU��UUU�UUVdHUEUQUUQUUUUUUUUTEUUUPUU�UUUa�iUU�UUVdHUEUAUUQUUUUUUUUTUUUUQUUUUUU`�YUU�UUVeUEUEUUUUUUUUUUPUUUUUUUUUUh�UUU�UUVe(UEUEUUUUUUUUUUQUUUUTUUUUUX�UUU�UUUV% UEUEUUEUUUUUUUQUUUUETUUZiUX�UUU�UUUV� UEUUUEUUUUUUUEAUUUUQTUU�ZX�UUU�VUUUh UQUUUEUUUUUUPEUUUUPTUU�UZ�VUUeUUUUH(UQUUUEUUUUUUAUEUUUUTTUUUUZeUUUeUUUUXUUQUUUUUUUUUUQUEUUUTPUUUUVeUUUeUUUUXUHUQUUUUUUUUUUQUEUUUUQU UVeUUUeUUUUHUHUQUUUUUUUUUUUTUEUUUEUQU*T�VeUUUeUUUUHUUQUUUUUUUUUUUTUEUUUAUQU�P�UeUUUeUUTUHU(UQUUUUUUUUUUTUEUUUQUAU��R�ViUUUeUUXHU�TUUUUUUUUUUUUTUTUUQUEU�R�UiUUUeUUXJU�TQUUUUUUUUUUUTUEPUUPUEUaEB�UiUUUeUXBU�PQUUUUUUUUUUTUEQUUTUEU`EJ�ViUUUeUZRU�RQUUUUUUUUUUUUEAUUTUEhU
aViUUUeUZRU�RUUUUUUUUUUUUUEEUUTUEJU)aViUUUeUVVU�RUUUUUUUUUUUUUEUUUTUE�B�%aViUUUeUVVE�PEUUUUUUUUUUUUEUUUPU�@�&`UjUUUeUUVE�TUUUUUUUUUUUUUEUUUQU�D��hUjUUUiUVUV�TUUZiUUUUUUUEUUEUUUAU�T�&XUZUUUYUVUU�PUU�ZUUUUUUUEUUEUUUEU�T��XUZUUUYU�VUU�RUU�UUUUUUUUQUUEUUUEU�T��ZUZUUUYU�UUUVRUUUUUUUUUUUQUU@UUUEUU T�VZ�ZU�UUU�UVU�RUUUUUUUUUUUUUUDUUUAUU T�jZ�ZU�TUU�VU�Ri�UUUUUUUUUUUUDUUUQUU U�jZ�ZU�TUUeVU�R�jUUUUUUUUUEUUTUUUQUU(U�jY�VU�TUUeVU�RUVUUUUUUUUUUUTUUUPU(U�jZ�VU�TUUUVU�RUUUUUUUUUUUUUUUUUTU*U�jZ�VU�PUUUVUERUUUUUUUUUUUUUUUUUTU&U�jV�UU�RUUU�VUERUUUUUUUUUUUUUEUUUTU&U�jV�UU�RUUU�UUEBUUUUUUUUUUUUUEUUUUU&U�jVeUU�RUUU�UUEJUU PUUUUUUUUEUUUUUV��jVeUU�RUUU�UUUJZi��BUUUUUUUUAUUUTUV��ZVeUUUjUUU�UUU�J�Z� JUUUUUUUUQUUUUTUV���VeUUUYUUUeUeUUI�U!HUUUUUUUUQUUUUTU�V���UeUUUV��VUUaUUIUUaTHUUUUUUUUQUUUUTU�T���UeUUU� ZUU�UUIUUaTUUUUUUUUQUUUUTU�T���UUUUU�  hUU�UUJUU`�*UUUUUUUUUUUUTUaT���UeUUU&  `UU�UUIUUh� UUU UUUUUUUUUPU`TY��UUUUU&��`UU�UJUX� UUTUUUQUUUUQUhTY�fUUUUU&��`UU�U*UZ� TUTUUUQUUUUQhP��fUUUUU�  hUUPU*UZ��TUTUUUUUUUUQjP��fUUeUU� XUU`U&U�j��TUATPUUUUUUUQ�VQ��fUUeU����ZaU&UhZ��PUAPPUUUUUUUU�PU��eUUe�""
���h�U&UXZU�RUQAUUUUUUUU�TU��eUUe�PE��UQ`�U�&�jU�PEQ UUUUUUUU�T��jiUU%�TU��UUa�U�&�jU�RUP@TTUUUUU��U��V�UU%�U��EU`�U���jU     @UUUUUU U����UU%��     h�U���jU*P   PUUU���(U��f�UU%U������Z�U�U�jU�RUUUUUUUUUUU����f�UU�UUYYUU�U�U�U
��UB�����U������Z� �feUU�UU�����U�U�U	��UR    ��   �*��J�jeUU�UU�����UeU�U��UUUUU PUUU   @�jUUU���Z����UaU�U(��UB@@TUUUUUUUjUUU�������jU`U�U���EUUUUUUUUUUA`UUU��Y�����UaU�U���UBA@TUUUUUUiUUUU�������V`U�V����UUUUUUUUUUUU@ZUUUU�����j�VeU�Va���UR@@UUUUUUUUU�VUUUU���j���VUU�Ua���UUUUUUUUUUUUUUA@XVUUUUf��j���ZVU�U����U*AUUUU UUZVUUUUf������ZVU�U����U�UUUUUUUUUUUUU�ZUUUUUe����j�ZVU�Ua���U@@ QUUUUUUUU�YUUUUUi��Z�Z��VU�Ua���ZUJUUUUUU  U  ��iUUUU�Z��jV��jUU�Ve��XUYUUUTUUU���j�eUUUUU���jU��jUUUVeY�XUY  @UUU  ��UUU�eUVUU����jU��jUUVei�XUY���  ����U��eUVUU�����Y���UUVee�XUYUUU���jUUU  `eUVUUU��������VUVUe�*VUU�UUUUUUaeUVUUU��������ZUVUe�(VUY  D U       `�UVUUe��������VUUVU��(UUUi�UVUUe��������jUUVU�V�UUU              XUUVUUe��������fUUVU�U�UU�ZUZUUe��������VUVU�T�VU               jU�UUe��������VU�VU�T��T�U�UUe��������VU�UU�Q����               ���UUe�"
  ���jU�UU�UaU���ZU�  �ZU�UU�UiUUU                  ��*        �jUU���ZUUU   �jU�UUUUUU                              ����UUUUUU    QUUUUUUUU                               UUUUU        UUU                                UU         PU                                                                                                                                                                                                                                                            @                                                 @        @                                                                                                          @                      @                                                                                                                       @         �(U%                                      U% @DAQUUQEUT          @TUUQQUU%                ����     @ @   @  U% @          @    ����*      @      U% @         @    ������    @ @      U%            @   ��  �*   @ @      U%PQEUQUUUQUEU  �*TeU���  EQUUUUQU%              ��BUeU�*         �* @             �*TUeUU��"           @           ��BUUeUU��           @            ��TUUeUU�*          @PQUUEUTEE �*UUAeUU�* QUUUUTA          @    �JUU eTU��                 @    �JUUAeUU��                    @    �RUUUeUUU�                 @    �VUUUeUUU�          EQUQ@UUTUUA  �RA e@� UUEUUAU         @      �V �*e�J�                      �VA�*e�J�                   �RU�*e�JU�                   �VUJe�RU�      �*TQQUUDUTUUTEQ  �VUJe�RU�PUUUEUUUEU              �RU�*e�JU�                       �VU e@U�               @     �VAUUeUU�       �*      @      �R UUeUU�       U%PUQU@@UUUUEUE �VAUUeUU�UUEUAUUUU%         @   �VUUPeTU�       U%   @     @   �RU@ePU�       U%     @     @    �VUUPeTU�        U%                �VUUUeUUU�           U%                �����������          U������������������BUUUUUUU������������U%                �@UUUUUUU(           �*                 @UUUUU               PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P                 UUUUU                P                 UUUUU                P                 UUUUU                P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�* P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�* P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU% P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�* P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUU                            P@UUUUUUUUUU                            P@UUUUUUUUUU                            P@UUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUU@UUUUUUUUUUUUUUUUUUUUUUUU   P@UUUUUUUUUU@                          P@UUUUUUUUUU@                       �* P@UUUUUUUUUU@                          P@UUUUUUUUUU@                          P@UUUUUUUUUU@    ���
  ����   ���
     P@UUUUUUUUUU@           �       �* P@UUUUUUUUUU@           �       U% P@UUUUUUUUUU@ ���  ���*  ����  ���U% P@UUUUUUUUUU@ VUU  XUU%  �UUU  XUUU% P@UUUUUUUUUU@ VUU  XUU%  �UUU  XUUU% P@UUUUUUUUUU@ VUU���ZUU����UUU���ZUUU% P@UUUUUUUUUU@ VUU  XUU%  �UUU  XUUU% P@UUUUUUUUUU@ �jU  XUU%  �UUU  XUUU% P@UUUUUUUUUU@ ��  ���*  ����  ���U% P@UUUUUUUUUU@                      �* P@UUUUUUUUUU@ �����*��������*�����*   �BUUUUUUUUUU@                         BUUUUUUUUUU@                         �BUUUUUUUUUU@                         ����UUUUUUUU@                         ���UUUUUUUU@                         ����UUUUUUUU@                         �XbUUUUUUUU@                         ��h�VUUUUUUU@                         P�j�VUUUUUUU@                         P `VUUUUUUU@ �*                       P �"VUUUUUUU@                         P  VUUUUUUU@                      �* P���VUUUUUUU@        �����           P�*�UUUUUUUU@ �*      �    
           P�*�ZUUUUUUU@ V%      hPT)           P(
hUUUUUUU@ V%      HR�T%%        �* ���`UUUUUUU@ V%      HB�P%$        U% � ��`UUUUUUU@ V%      XB�P)$        U%��*���VUUUUUU@ V%      �F�P)$        U%����"VUUUUUU@ V%      �B�Q*$        U%�*  
*VUUUUUU@ V%      �F�Pj$        U%�&VUUUUUU@ V%      �F�Q*$        U%�**&VUUUUUU@ �*      �F�Qj$        U%�**�&VUUUUUU@        �F�Qj$        U%�(j)VUUUUUU@        �F�Qj$        �*�(� Z	VUUUUUU@        �F�Qj$         �����V�VUUUUUU@        �F�Qj$         � ���VUUUUUUU@        �F�Qj$         �*P�j	ZUUUUUUU@        �F�Qj$           P"b�VUUUUUUU@        �F�Qj$         �*P�jUUUUUUUUU@        �F�Qj$         ��R�UUUUUUUUUU@        �F�Qj(         � ��UUUUUUUUUU@        �F�Qj
         �* �UUUUUUUUUU@        �F�Q�          ���UUUUUUUUUU@         ����            P�UUUUUUUUUU@ �*                       P@UUUUUUUUUU@                         P@UUUUUUUUUU@                      �* P@UUUUUUUUUU@                         P@UUUUUUUUUU@ �*                       P@UUUUUUUUUU@ V%                       P@UUUUUUUUUU@ V%                    �* P@UUUUUUUUUU@ V%���
  ����
   ���*  U% P@UUUUUUUUUU@ V%    �           U% P@UUUUUUUUUU@ V%    �           U% P@UUUUUUUUUU@ V�  ����   ����  ���U% P@UUUUUUUUUU@ VU  XUU�   XUUU  `UUU% P@UUUUUUUUUU@ VU  XUU�   XUUU  `UUU% P@UUUUUUUUUU@ VU���ZUU����ZUUU���jUUU% P@UUUUUUUUUU@ VU  XUU�   XUUU  `UU�* P@UUUUUUUUUU@ VU  XUU�   XUUU  `UU   P@UUUUUUUUUU@ ��  ����   ����  ���   P@UUUUUUUUUU@                         P@UUUUUUUUUU@                         P@UUUUUUUUUU@                         P@UUUUUUUUUU@ QEDUUA         PU   P@UUUUUUUUUU@      @     ����   @'
UUU�UUUUUUUUU	ZUUUUUUUU%�UUUUUUUU�VUUUUUUUU
XUUUUUUUU)`UUUUUUUU��VUUUUUUU�XUUUUUUUU
`UUUUUUUU)�UUUUUUUU� VUUUUUU��XUUUUUUU

`UUUUUUU)(�UUUUUUU�� VUUUUUU��XUUUUUU�

`UUUUUU�*(�UUUUUUU�  VUUUUU�  TUUUUU�  �_UUUUU� �_UUUUU�*��UUUUUU* �_UUUUUU���UUUUUUU��_UUUUUUU��UUUUUUUU�_UUUUUUU��UUUUUUUU�_UUUUUUU��UUUUUUUU�_UUUUUUU��UUUUUUUU�_UUUUUUU��UUUUUUUU�_UUUUUUU��UUUUUUUU�_UUUUUUUU�UUUUUUUUU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUU����UUUUUUUUU�� jUUUUUUUUU�*�VUUUUUUUU��hUUUUUUUU�
(�VUUUUUU����XUUUUUUUU�
 `UUUUUUUU� @UUUUUUUU*  �UUUUUUUU�
��UUUUUUUU��_UUUUUUUU���UUUUUUUUU��_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��UUUUUUUUUU�_UUUUUUUUU��jUUUUUUUUU��VUUUUUUU�� jUUUUUUUU���UUUUUUUU�  �VUUUUUUU  jUUUUUUUU% ��VUUUUUUU� 
��ZUUUUUUU
��jUUUUUUUU� 
XUUUUUUUUU
��UUUUUUUUU��jUUUUUUUUU� ��ZUUUUUUUU��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUU�jUUUUU�_UUUU�ZUUU���UUUU��VUU% �_UUU�
hUU% ��UUUU)�VU	 ��_UUU�
hU	����UUU���U	 �U�_UU� V	�jU��UUU* X%�jUU�_UU�`% �UU��UU�*`� �VUU�_U���U jUU��U��U	(�VUU���*�U��ZUUU��� �UU
�UUUU�/`UU��ZUUU�� `UUU*hUUUU�XUUU��VUUU��UUUUU�jUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU0UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUU�UUUUUUUUUU��WUUUUUUUUU%�WUUUUUUUUU%�_UUUUUUUUU	 _UUUUUUUUU	 UUUUUUUUU� |UUUUUUUUU� �UUUUUUUU�  �UUUUUUUU� ��WUUUUYUU���WUUUUYUU%���_UUUUYUU%��j_UUUUYUU%��YUUUUYUU	�fY}UUUUYUU��UU�UUUUiUU��UU�UUUUjUU��UU�WUUVjUU��UU�WUUVjUU��UU�_UU�bUU�UUUU_UU�bUUiUUUUUU�bUUeUUUU}e��`UUeUUUU�e��XUUeUUUU����XUUeUUUU���"XUUeUUUUՋ� VUUeUUUU��VUUUUUUUU VUUUUUUUU? �UUUUUUUUU= �UUUUUUUUU� `UUUUUUUUU� `UUUUUUUUU�XUUUUUUUUU�XUUUUUUUUU�VUUUUUUUUUU�UUUUUUUUUUU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU0UUUUUUUUUUUUUUUUUU�VUUUUUUUUU�hUUUUUUUUU% �UUUUUUUUU	  UUUUUUUUU _UUUUUUU�  _UUUUUUU� ��_UUUUUUU% ��WUUUUUUU%���WUUUUUUU	���UUUUUUUU����UUUUUUUU�h�~UUUUUUUU�Z�UUUUUUUUbZU_UUUUUUU�hV�_UUUUUUU�XV�WUUUUUUU�ZU�WUUUUUUU%VU�UUUUUUUU�UU�UUUUUUUU�UU}UUUUUUUUeUUUUUUUUUUeUU_UUUUUUUUUU�_UUUUUUUUUU�WUUUUUUUUUU�WUUUUUUUUUU�UUYUUUUUUUU�UUYUUUUUUUU}UUZUUUUUUUUUUZUUUUUUUU_U�XUUUUUUU�_U�VUUUUUUU�W�%VUUUUUUU�W�)VUUUUUUU�U��UUUUUUUU�V��UUUUUUUU�V)�UUUUUUUU�Z
bUUUUUUUU���`UUUUUUU���XUUUUUUU�� XUUUUUUU�� VUUUUUUU�   VUUUUUUU�  �UUUUUUUUU  `UUUUUUUUU XUUUUUUUUU)�VUUUUUUUUU�jUUUUUUIUUUUUUUUWuUUUUUUUUUUUUUUUUUUU�_�uUUUUUUUUUUUUUUUUUU�?�|UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\UUUUUUUUUUUUUUUUUU�?�\U�uUUUUUUUUUUUUUUU  PU��UUUUUUUUUUUUUUU���_U5�WUUUUUUUUUUUUUU3sU5�WUUUUUUUUUUUUUU<|U��_UUUUUUUUUUUUUU  |���UUUUUUUUUUUUUU0\s��WUUUUUUUUUUUUU�\s�  \UUUUUUUUUUUUU� ��s= ��UUUUUUUUUUUUU5�?�p= ��WUUUUUUUUUUUU� ���=   �UUUUUUUUUUUU����=   �UUUUUUUUUUUU?����=   �WUUUUUUUUUUU0 0��=0   WUUUUUUUUUU�? 0��=0  WUUUUUUUUUU�? 0�_?0  ��UUUUUUUUU�� ���?�? ��UU]UUUUUU�?� � �����wU]UUUUUU�?���� |U����UUUUUUU�?���� \U�����sUUUUUU�?���� \U133�pUUUUU�   � \U�   \UUUUU�?� ��  pU00 _UUUU��3 �  pU3���UUUUU�   ��   pU3��uUUUUU=   0��   �U3  �uUUUUU�   <    �u��?uU�WU}�      ����uU�U�  <33  �����uU��W ���    _���uU��� �   �?�  � ���wU����    ��� � � ?UU�=� <0   ��� � 0�UU�5 � 0   � < � ��UUU�� 0  ���3 � ���UUU�0�0    <�����}UUU��  �  ��W �UUUU�� �<��W �zUUUU= <<3�� ���� 0�UUUU�����  �� �?0VUUU�?�����0������00XUUU����� �<�0`UU�����  <  �����`UU��?�?�  � � ���0<0`UU���<0?  �������?0 `UU�����  �  �0�`UU�����  ����� �`U�����  ����     XU	��?� 0������      XU����� �0����     �V� ��?�? �00  �     jU�   00 �0���<   ��UU%    00 �����<  �`UUU% � 0� ���<   �UUU%  � 0 ���<    VUU%   �?  ����?    XUU�   (   <��?    `UU�
  �00 �� �  �* �UUU)  �0? * 
�  � �UUU�  �  �   ���  `UUU�
 (     �     � XUUUU��             VUUUUU%           �& �UUUUUU�           j� ZUUUUUU���      ��UU�UUUUUUUUUU�    ��UUUUUUUUUUUUUUU��
 �VUUUUUUUUUUUUUUUUUU��UUUUUUUUUUU   @   �@L�!�B���� L� �,�"@�tB �@��"�"	�H�"�"� HH�!@ HH"�!����D"��LD"D@
 D" `	�B3���� H�8?� ���������������w�U�" �� "�U�w���������������PPPii�Z�P                                                                                                                                                                                                                                                                                                                                                              �����*�����*(    ((    ((�?�?((�?�?((<<<<((<<<<((���?((���?(( <<  ( <<  (�����(�����(<<<  (<<<  (�?<  (�?<  (  <  (  <  ��*<  ��*<     <  ���*���*(�((�((��((��((�"((�"(���*���*        ��������   <  ��*<  ��*<  (  <  (  <  (�?<  (�?<  (<<<  (<<<  (�����(�����( <<  ( <<  (���?((���?((<<<<((<<<<((�?�?((�?�?((    ((    (�����*�����*   <��*<��*<( (<(((<(�*<(  <��*<��*<  (<�*(<(((<( (<��*<��*<   <��������        ���*���*(�"((�"((��((��((�((�(���*���*T      @� ��  P    �@��  ���P    @����� "P    @� )D "P    @��""��&R    Т���B!�S    Q��� B!��    �B�@����P    9F��    ��    D� �����Q    @�� ��@�Q    @� B@�@    @� B �D    @�B�D    AP����BQ`"�    � �  @���                  ��@�  � �  ���@�� ��! �@�@�D AP�� �B�@�1L� *�� ��Q�B���@� �����C�!D���� �����DOw�@�� �Q�@�Q�8�@�@ �F����D! �� ��A�D����Q�! �B�A�D@ �Q�� �B�@�!Ǡ���Q�  ��D�!t!	@�ь�zB�D�$
 �@� ��(B���A����   � ��   @ �                   �@   @   �@! ��@(�.�  �A�DP�@�B  �BH���B�R�N�  D@*� KP�S0��@ ���j��`%@�1 BP��J�p`R�ȃ!B�E!�O�`���r��H !��A0� � N�	J�AR  ��� B� z�M�  D�� B@	 J�A�    ��� .�AJ�A  B!���" ARB��  B&�����r!BB�    ��  pB�                 �     ��   ��     @��  �� @  @@  �� ��  ��@  ��@��D@@  ����@0D@@  �� @0O�B ��@D@��������� D@@  �� @P ��@  �� @0 B@  @@  B�@  �@�  B��@  ���  *�@  ��`@@�  @@  0           @                  @  �           N� ��          @@ �!          @  �!          ���          H���0          L� � ��      HB� ��      HB�!��      HB $A��      �B $�          t"@$@          ""�$�          ��          �A`(           �            v      @� � @     �@�� ���@     @����!)@     @� �!)@     @��"��)@    Т��0����    Q���� %@     �B�@� #@    9F��  �!!@    D� ��$A��     @�� $�!@     @� $@!@@    @� $�!@�    @��!B�    AP����(-�`    � �  �                             !  ��,�@�  ���� ��H�  ��B � @��*�DDB �@@0-�(B��d@�10 �R!BD!@ȃ��R""!����r ��B���@P�  ��B(�@0�� ���B(�!@�  ��B��b!@���  ��(N�����  ��(@@@瀱  ���(�@A    �  �@  @�                   @  �   ""��@  �  �����!D@  ��   �DB  �B �� �@�L��B@��*�"�B0�B��@@!�bDB0�B @ ���DB��@��)�� �B ���  * ��DB �  @  * ��D" �  @��j ��D"  � @@��� ��O"  ��@��( ���  �����$ �@(A  ��`@��"  �  @                          @  	   � ��  	 �@�� @  	 ��@  ������ @@� �!��@ 0���B"@� 0��""@�"�������� �P@@  �0 b@ B �bB@��  ��B� �@   ���0@��   �@@�� A@ A  � A  � �   �  � �                   �        ���  �!  ""����Q@"���  M�@  R�爀!   ��O�  ��$��!P  A`@  �@$IA)�0-��� ��P,JB/�`@���B$"*"!`	O�  �R�B�q`��@  �R$B�
A0KO�  �Q$��
A  )A  �A$ �A  �! ��$ zq  	!��N��*  	�  "%$A���A  I�   �  �  �                          �   �� "@ O�.��` !��� �B�� ���B�   N�   DB���� � (Bhh!l1� �"�RM�D&D!p�� �"R$!O�@�!B�!�!!A��@�!B�!@!�!AR��@���Bd!p��1M򄐀��@BD!@@d!A���dD!@ @A@D�D%@@�� (�B%L @A ��   A&C @��0                   �            @ ��            � ��             B"            �J�            h!b"            D&^���        $@ ��        �!L���        @!D��        p�D            @@L�            @ D            @D            L L�            C D            !          �         ""   ����       M�` !�!""      �� ���!��      A`   ��    -� � �0�0     �"� �0    	 �"� �    ��@�!�!�     K@�!$A��     )@��$���     񀀄@$@�@      	��d$�A`      	@D��B�      I� ((*      �                     @� ��       �@�� �!��      @�����!      @� � �!      @��"����      Т��P�00    Q����� `    �B�@�� `    9F��  ��!`    D� ���$A0    @�� ��$�      @� ��$@      @� �P$�      @��`�      AP������(      � �  L      e      @�         �@�� ���@     @���*�D�     @� %�D     @��"!PD�    Т�� ��h!    Q���)�DD&    �B�@%'D�$    9F��  ""DR�!    D� ��*��R@!    @�� * DQp�    @� i!D�@@    @� ��DQ@     @�  DQ@    AP����  %6L     � �    C                 �        ��    ���  ��  ����Q!@�!��B"  @  R!@L�""J�O�  ��!B! ""b"0@  �@)�"""^�0�� ��P)B��""@ @���B)B� ""L� O�  �R)B�!""D @  �R)B��""D O�  �Q)B� !�L�  A  �A)B� �D  ! ���  D  !��NԈA�0��L�  �  "%@@�� D     @�                    �  H�  H�  �� ��H�  H�  @ �N�  N�  @� �H�  H� "� ��@ @ �� �!� �P0�P( ���H�0H�(�� ��DD$@ � K� K�$(� �@  @ "b �@ ��L� L�!�  @� �  ���@�@D�t  t ��pBB$  $ @.��/��  � �                           @ @�  H@�@�@�� �� ���D@@���	@��DB@� �B� L�@��"DB���H�BТ�(B ��DBQ����R� 	PDB�B�@R�/r �B9F��  BE!B
@DBD� ��BE!B	�D"@�� �B!!B�D"@� B�/rhO"@�   �@�  �
 (AAP�����   �� �                         @@�    � �@� @��D ���@� �� L� �D@ ���B� �DB��@�D.2	Bmw  
0@D""�@���
@�""�@N 	 �pD!""��BQ 	@P  D�""�NQ����0��D@.2�BQ H��Ǡ""��NQ (���t! �@BQ@ ���$��B@
 @�� �BQ��   ��   �J�                  �               �               �               �              ��              �R0            �R`            �R`            �B`            �"0            �"              �"              �              �              �A              ��              e                  ""   ����@     M�` !*�D�     �� ��%�D     A`   !PD�    -� � � ��h!     �")�DD&    	 �"%'D�$    ��@�!""DR�!    K@�!*��R@!    )@��* DQp�    񀀄@i!D�@@    	��d��DQ@     	@D�  DQ@    I� (  %6L     �    C                 �        ��    ���  ��  ����Q!@�!��B"  @  R!@L�""J�O�  ��!B! ""b"0@  �@)�"""^�0�� ��P)B��""@ @���B)B� ""L� O�  �R)B�!""D @  �R)B��""D O�  �Q)B� !�L�  A  �A)B� �D  ! ���  D  !��NԈA�0��L�  �  "%@@�� D     @�                    �  H�  H�  �� ��H�  H�  @ �N�  N�  @� �H�  H� "� ��@ @ �� �!� �P0�P( ���H�0H�(�� ��DD$@ � K� K�$(� �@  @ "b �@ ��L� L�!�  @� �  ���@�@D�t  t ��pBB$  $ @.��/��  � �                           @ @�  H@�@�@�� �� ���D@@���	@��DB@� �B� L�@��"DB���H�BТ�(B ��DBQ����R� 	PDB�B�@R�/r �B9F��  BE!B
@DBD� ��BE!B	�D"@�� �B!!B�D"@� B�/rhO"@�   �@�  �
 (AAP�����   �� �                         @@�    � �@� @��D ���@� �� L� �D@ ���B� �DB��@�D.2	Bmw  
0@D""�@���
@�""�@N 	 �pD!""��BQ 	@P  D�""�NQ����0��D@.2�BQ H��Ǡ""��NQ (���t! �@BQ@ ���$��B@
 @�� �BQ��   ��   �J�                  �               �               �               �              ��              �R0            �R`            �R`            �B`            �"0            �"              �"              �              �              �A              ��              e      @� � @      �@�� ���@      @����!)@�    @� �!)@    @��"��)@�    Т��0��    Q���� %@    �B�@� #@    9F��  �!!@    D� ��$A��    @�� $�!@    @� $@!@    @� $�!@    @��!B    AP����(-�      � �  �                     @     @    �@ ��  ��� ��)@@  �@D �� )@  �@L�  )@��  � � ���  � D.2�%@� ��D""�#@�� ��""�!@�  ��D!""���P  ���D�""�!@0  ���D@.2�!@  �@PǠ""�!@� ��@0t! ��!B���(�$��@P-�@�����   �       �                    �      � p� !    �� @��� �  �P@@ �H�  ��@���	@��*�"�@	@  �R@0
��!@����R�10� @  �Rȃ� �@r �B�r ��@��@��"�  � (�@p �"�� ���@@@ �"�  �# @@p@���  �"�@@@@���  I pB��@��A��  ".�@P  ���  �                            � @@,�    ���!�@��  ����Q��@�"  @  R)@��.�O�  �� �D$"0@  �@��	B%"0�� ��P �@���@���B �@��"! O�  �R����D�"! @  �R  �t�" O�  �Q��D�"  A  �A ��D�  ! �� �@D"!  !��N� ��D� A  �  "% �D �     �                �    @� @@  �P  �@�� ��$@  ��  @����D@�!�!  @�  O�!��@��"/2@��R0Т� "@  �!0Q���$"t@���Q�B�@$"DB� �� 9F��  ""O��`�" D� ��.�D@���� @��  �D@�#�  @� ��D@�"�R  @�  �B@� ��  @� ��@A ��  AP���� B�" B  � �     �                   � �       (� �!      ��F� !@�       �"�"!@�       B"��!B��      �"�)��"0    @�"�)B��`    @�2�)B�"`    p�"�)B��`      ����)B�"0    ���!��)B��      ��� �@)B��      ��� ����      ��A ��A��      ��.��@@��      ��  D @�@         @   �@L�!�B���� L� �,�"@�tB �@��"�"	�H�"�"� HH�!@ HH"�!����D"��LD"D@
 D" `	�B3���� H�8?� ���������������w�U�" �� "�U�w���������������PPPii�Z�Ph(                       Pn       @U                            ���
                                   ���*      TQU                         ����	                                  ����                                 ���U�                                 ���Z�j                                @�ZU�                                 �j��         �                 @ `U  �����        @�                 �jn� �����       @��A              @�UU  �i����f       e�j             �j��	 �������      �V�U  Q         �����[}$RЯ�ﯹ     �Z�TU P         ��������[E��C   �j�  P  PQ      ������������V��   @��   @        Ц��j�����ڪ����   ��    @P        Ц�����������k��  ��j      P P@     ��j�몪�ڮ�ӿ� ���      UPP      @���ꪪ�皪����j� @Z�       AU        ���ꫪ�ۚ���K[�yBj�     @      �ki�櫪�n^��ZE�.�Uj  X    @T      �U��ꫪ��y��@�[d�       TFPP@   @����ꫪ��皫땁֦Tn      @fT@PUP    �����������뻔۹i.U
  TP��!  @P     ���� ����nn�������� P��*   @    ���z �꿥������P���[�  P��[ P  T     ���/ ����������km�o��V� P��  @ @    ��� ���V꿮��������ZU� PV�P       ��� Ы�jU���뿩���U���Z.
 D     ���  𫺪Z����o����������*�]     ��  䫪�Ze�������[��Z�����GPT@U    ��  ������������j髪����.��R TU    ��  ����������������V���.��       ��  �ꫪ�[�����ꫪk�����?�j P      ��  ���������������Z�����
TU@     ��  @��j����������������Z  TU P        ��  �������鿫�@����k TUU    P     � P�������j���   ��j  TU  @   P      `�@i����������/         @UUUP          T���������꿪�          DQT   P@    h��j������ꪪ�          @T    PP   o������������        P   TU  @ @   �k� �j������j       UUUUQ @@@ P  PZ��  骪������    D@   TU@P     @j��~ P������Z��        @          啮�/���������j>         @U     T  @  �� �A�
����릩�       T       P ���  �e�[�����z        P         ���   }�_忕����            U    D��   ����������                T@��    ���n�����.                   ��o    �Vk[�￪nj�                   ��� @  ����������                   P��     �j������o                   @��    @�nU�������                   ��o     �������ﺪk                   ��    ���Z������/                   � @    �U��������                      @  @�U���������                  P  T   к����������                  PP �j�_����������                  E PA@VU��e������oU�                  UU P�PU��T������oU�                  TU@P�jUiyh��������                  PQ@ADVj)m��������                  U ��e���������o�/                  UUT @�*iZ��������Z�z                  TQUA P�������oj��                 UUEU   i �����������@ @            PTT@   ��A�������              TEEU T@U  ���������VA@           ETU  TU ������jU�  P             UUP TTU �_�����U�� @@  @         T@U U  ����������    DUE         U @PP U @����������   T          PU    PU���������ZY)      A       P P @    �Z��o��Zk�*         @       PP     ������j���k        @       UA     �����������                APU     �e�A������      @       PTT     �������꫺               TPU@UE  @O�z  ������                QQU PA  T��k  ������                QUPUP �����   ������                 UPU@  ����}�  ������                @@U  ����n�[Qi������                UUU  @Zi�������������                UU  E ��j[������j�����.                UPT@U���V���b`T�����:                ATAPEUUUU�Z����j(�������                UUUATUU�U�����m9������                PUUUTU ���U����n������               PUUPUUU � 4����￯���               @UUU ���  	 ���뿪���                UUP �  @ ���������                  @A $  U�   �z������                  U  ��  @������z               UUEUD $�  @    ����.@              TU P�j        �����P                TPU         ����TA              U UPPA   P    �����BUU              P  PQQ   T      i �PEU              UPUAU   TU        @PTQ              �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� |ȥI�	�G 1��dG�G

i"�� i��l  ��` ��`  �` G�` ��` F�` p�` ��` p�``�I�& 逐<�Hi��(d)$*���� �V���W �� wˀ��dI ������H�H��dHdG��I`�I�� �����Hi�������'�q�=�M�)�'����'�G 1��������' �ҩ������'��'�G 1���'Ύн8`����'�=�$�)�'����'�G 1��������' �ѩ������'��'�G 1���'Ύп8`H�ZH����\�]����\����&�'����&������m��8����m��h)���� ��6� ��.�)������������� ��� ���8z�h`1�'�1��-�1�!��!���!�������������#0.��0101��*+��2/��2323��('��()()��H�Z�?���L`��G���E� ��?�;��� �;�{���;�������;�������� Ԇ������
�8�� +�� ��?}�����>�;
m>��ˁ�ȹˁ��8
���ȱ���:�?�;���{��� �?�;�8���>�?� �8.>ʀ��.->�.L���8����N�;��C�8��<dGdHdIdQ�H d���h)��h <�z�O�O�И�i��i��  ����O��z�h`�H�H�H�H�H�H����������� �� wˢ �ψ���� �� wˢ �π�h�h�h�h�h�h�`Hڮ?��>� �>ʀ��?����
�>I�-��>��h`H�Z� �8�'I�����8�&���?��z�h`H�8�&I��8h`��H�8�'I��8h`����6��d������6��6��^��0 ^0 ^F [ ^[ �  � �  � � � �    H�Z����E��x�E��y�E��z��x8�<�(n��0j�x�y8�>�y�z�?�z�z�Q�yɏ�J�8�xI��;�8�yI��,�y��x��

��e�)m��l��?���������'�L��z�h`   	!�Z�z�M���E��y�E��z�y8�>z�`H�Z�?�����������y��y�� ���ɑ�Lz��?�;� �Lw��?� �8 0��>� �8�&I����LC��Z��)�P�?���{ ���� ����?�;�b ��2� �8�'I���> ����?���{��?���ǩ���� ���?�;���)?����0Ȁ����I�� ���?� �8 7���?�?��L���N��	�N �� w�z�h`����] h��'�\�8�&����] 5���\��&8�\��`H�Z�?����]��\�?���� h��1������ 5��!������ �
 ������ ���� ����\��]�z�h`H��\���0 ����� 1����\������h`H��\� 0�& ����� 1���:�\�����I�-�h`H��l���h`8��H���0� h`8��H��] ���-�]���p0ɏ��\�] ����� 1���8��]���h`H��]���l ����� 1���i�]���h`H�Z��ɑ�G���������m����}�~�?���|� ��i��8���� �ʒ���ʒ��z�h`H�Z��ɑ�<�}�}��2�} Ғ �� w˭��|�i�8����~�~�
�� ����z�h`��6��d��6��0 ^0 H�Z����ʈ��ʈ��ʈ���8�<�0&��0"��8�>���?����ɮ��L���������}��'� 0����k�[ɑ�q��Z��[���
��$hp�i�h	@�h <۩Z����[����X����.)��.�?�? ����; 7� ����?������L�z�h`Hک���
�  ����1��0
�ɲ���ݰߩ�����h`��(��P��h��v�*v�D��X��q4�q��H�Z,�pL�������������������������8�<�(S��0O��8�>���?���	�ɏ�/����)���"��,����� k� Ê� ��.������L4�z�h`,�0+������������������ ����	���`�*)�*�w�(� �)��,����,����,����&��' j�`��6��Y��o�J��J & 9 L k2 H�Z���z�����������(���(���(����8�<�(a� 0]��8�>���?���D�ɏ�=� �i��i� k�(� !�� �z�~� ?�8�3�_ɑ���� ����.��z���Ld������+�Nz�h`�+� ɑ�R� ����I��,����,���,�e�z�����8��������)���F���+� ɑ�� �����*��+�������������������8�`�N����N� ����H�Z�z� Ӎ� �}�8��^ W��>�	����������^8���>i
�� ��O�����>�_ �� wˈ�� �ϩ��_ �� wˢ �πڥh	@�h Ӎ�i <ۭ.)��.z�h`H�Z�i���&��*)�*�&$*8����)߀�0�*	��*��ii���	 ���>��GdHdIdQ���y�3�z���� �Ύ�� �� w�  �  ��2 ���>�Ϣ� ��z�h`�y��ڭ���h�`8������ 		 	 	  		 	  	� �e�e')�� ��i
���������Ȁ�����������~`H� �����e�)��� ����~�h`HZ� ���J�������J����zh`H��0	8���������J����h`  ��d 9� q� 9եh)��h�y������0�X�\����Y�]�����	�
�t�(��)d&�j�'��
�h���������������
�{�����O����������z��{����`kjik����     '� �������(��)�>����(��)��> a� �ХE	��E���&�q�'�m> �
 �Ϝ����2�a��&�e��'�i��(�m��) �� wˢ ������� �Тx ��`�]��̢ �Ϡ
� ������ �ܰ����� S�Lr�� ���8��$*�&�%*�*��$��$*0�&��*�*���������� �G���G��GdIdHdQ`������i���i	� k�`Hڮ?�;��1�8��*���� D��?�� �
ʀ���.)�
�.�.8��h`H�Z���� ��,.p�.	@�.8�z�h`Hڮ?�����&��� �Ѱ�&� 1��*�&�&��"�&m��)��&�� 	Ѱ�&� 1���&� �h`H�Z�?�������y��y�� ���ɑ�L�� А�5�?�;��+�*���� $� �� w˩ ��(�\�?��;� �8�t ���H���� �ܥO� ��P� ����J� �������; ���F�;�(� �)dVdW � �� w˩ ��������?�?�LR� s�����N��	�N �� w�z�h`Hڭ?� ���:)��H�i�h	@�h <�h� �%8�#����h:)�h��8����:)�����h`��ɑ�Q�{�L�
�{��� � ����H��H� �x��K��K� �x�x�x�2�	� �x�������`Hڭ
��ʒ���ʒ������I@�������h`�������J� ��v� ����`�����`����������J� ���J������ k�8���� �� w˩ �����J��P�  ^ܢ �ϥO����P����P�  ^�`���� Ӎ�� ��_ɑ�8����^i����`8�� ǎ :��% Mݩ��� �)@��  � F��j o� q� ̉ ܈ x� ��� �[ɑ���_ɑ��h�@�')��h <ۀ�h�@�	@�h� � Ӎ�����i <�  � �� B��H�Ћ�.)��.����� �  '�L �    	HڥE� �Y�J�K���� �� �
��C��?��O����O����O����,L�O�� mH��I D�,.0�.	��.8��h`H�Z�G�6�H,L0i��I ���M��� ���,.p�.	@�.8��H��.)��.z�h`H�Z�'�Y��Hi���&i8�I��	8�z�h`H�&�"�0 	��H��&h`H�&��	 ���H��&h`,L0 K�� 4�`H�H8�&0�L)��L	��Lh`,L�H��H`,L0���Hڭ+ɑ�M�Ii�+�H,Li�*��~�	��i��*���~�)���z�~����(�����)�h`� � � Hڭ+ɑ�D�~��8�z�z��3�z�~�~
�����(����)�~� 0i�~m*�*����+�h` ���
H�Z�/ɑ�A�O�O��7�O�I�I��"��L�m/�/����.�.��.�.����/�Iz�h`H�Z�����*�+ k����+8z�h`H�Z�G�	��H���'8�
���&$*0i���%�/ɑ�4����.i��.���/i���H8�	I����	��z�h`�I8�	I��.���	��8��		

				L� n��	L
�HڥE� ���x��
�x�M�ޭH� 0��֭|�0����
L
��L
���e)��Hi���&i8�I��
 ��<�C��7�	��_��.�
 ��%�G�� ���_���K����O���0��S��M�N��O n��h`�G���������	�[���W�8`H�&8�HI��8h`��~���������������������ȘИ֘�
� � ��� � � ��� � � � ��� � ��� � � ��� � � � ��� � � � � � ��� � � � � ����� � ��� � � � � � ��� ��   �� � �  �  ��          �   �   ��  �����   ���� H�Z�O�LS��M�o��O�M����>�N,L��L���L��N,L�����mH�H |��M�	� �� ��L��������	������_�N� �mI�I�k�
� ���b���N��mI�I,L����@����;��>�N�� �����mI�I,L�
������Ь�N,L�)���$�mH�H�M
��Q���Q���N
���Jȱ�K����N�M� �� w˭.)�.z�h`�{�M���	�M�����M��M�NLB�H,L�H�0�H�
�H� �H�LI��Lh`� �� �ܰ����� S�L/���%����3����+��	�X��	���dF��� ���������8��G�*�G�.��0����������
������GdIdHdQ`  ���� 9թ��.��L���F�E���y�#�i�h	@�h <� �� �� w˩�x��O�MdGdS�a�I��N��X�O�I������z�.�{`���&�q�'��H�a�I��O� �M .���M�
 �dGdIdHdQ��O� �� .��M��` ��(�M�	���M�
� `�,.0�.	��.���{8�` 0��H�� �ȭ��H�E� ����F �� n� .� �� T� ��� Ŗ�@ n� �� �� ���|�a�I��M�N��O .��)��(���x �����/�RL� ��� Y�� 㛰L��| `� `� m�,J0/��x,MP"�
$*��GdHdIdQ �ȩ,{� ���ML��,{� ����G ���O�I��X��M�N�a�I��OL����/��M��N�x �Ơ�&8�HI��	 `� ����� �G���/� �� �� .��M��� �� '�dhL��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������d 9թ� q��� 9ե% M�d��O��� ��:�'�������������� �� �� �� M��&���'�8�	�*)�*LZ��'�Y��$*0�
���GdHdI�0�� �� �� �ȥG��L�.Z^/[_,X\-Y]悥��
�L��d��  ���ɑ�L��)�L����)��

m��+���	� ��*��/���	���.�Ь[���	���Z���� ���n��� ���ڲ��� k���<���������'����� ��
��	�
�o��� ��i�����1��� �� w˥G��!�
����&i���
���GdIdH���\����L�� �� w�`ڊ
���������������������轑�������������������`�*
�&i��'i� ���X��X >��8,J#� >��-�����'���#�i�' �� j֢ �π� >��
,J0��X��`�8��'`H�Zژ�0 ��he��e�����0����`�����������������H�@�I�J� �-H�"ȱ-H�ȱ-H�ȱ-H��I����JNHNHNINI����8z�h`H�G$*0"��;�<e&i�a�2�$�+�1�*�O�#�\�"����<8e&�����+��I��V��8h`H$*0�<e&i�$�#�1�"�O��\���<8e&���+��I��V��8h`H�Z�O�O��E�O�+ɑ�>�<e&�d�2�&���)���K�(��	����K���*�'i�+�L=������������*�+ k������A�*,K08��*�*��0T�i�*�*�(0�C�I�iw�(��) �� wˀ-�G��'�
�#��,K0�
���GdIdH���\� �����+z�h`�'ɀ�i�' �� j֢ �π�` }�� 9թ��g�h��i�
�j� �k��z�!�{���$������������d��O�I�E	�E ����� <� �� `� �� � d� ���i��� gĥE)�E � �� v� �� ��$h0�&���'�Y�� }󩙢 � '�L[��
 � gĩ |� �� gĩ��h�'�\�n�]d}�n�^��_ �� wˢ ���\�^�n�
�^��_�
�n�^��_�\��ЩS�]�l�^��_��*�.�Z�+�$�/�H�[��(�,�X��)�-�Y �� wˢ �ϭ^�l�
�^��_�
�l�^��_�]8��]���ͩ��[ �� wˢ �ϩ��/ �� wˢ �ϩ��+ �� w�` ����]�l�^��_ �� wˢ �ϩ'�] �� wˢ �ϩJ�] �� wˢ ��d}�\�&����}�n�]�n�^��_ �� wˢ �ϩ4�x��y`$hp ]̐d}�h	��h��l� �� <�Lc��m�L��d|��	��4 �̀� �ͥo��ޥn�ڭ�ɑ�ө������\i�����Lc��o�&�\�����'�H�*I�
hi�&�
� ̀ 4� ��Lc�$|0���|�l�^��_ �� wˀR�\i0�&�8�0�&��)��5I��&��)��&�k�p��q����l�p��q���m�r��sdndo`H�Z�+ɑ�L��I�I���I�\i8�*0 �	���m���8�+0���+i$>��)����������������������(�)�+8��+0$�-�i <۩�p��q��m��r��sdndo� �����+�E	��Ez�h`H�Z��ɑ�O�O�O�
�E�O���� k���i$��Ɂ�% �� wˀ"�G���
��F	@�F�
�GdIdH� ������z�h`$h"p#�j�k 5ְ ]̐�h	��h�n�n� �� <�L9� �� �˥m�L��d|��Q��5��
��Lr�LT��o��n�,�p��	@��,�� �ͥmдL�� �ͥmЪ ��dh <� �� w�L9��o��n���	����\$}08��i�\ �ͥo��A�n�=,�8���G��/��z dΩ�z�"$}0 q� q� q©
�  �  �  ©�GdIdHL9��o�$} ̀ 4� ��L9�$|0���|�n�^��_ �� wˀ�8�\�&I��z����}�i�z�7L:�ͬ�d}�
iͬ�$L:���	�)�DL9���G��)�5�K)��E�j�p��q��m�rdndo,�p
����
�� �˩���s`�n�p��q��m��r��sdndo`��m�n�p��q��s��rdodn�� Ͱ�ީ�d 9ե% M� ��d����
��x�y�z�{�|��}��~������������� �� �� g� ��&���'�Y��*)�*L֬	)>ltvi*.Z^+/[_(,X\xyz{|}~	,M0E�G���&e<i� �Ī�������'�&e<8�� �Ī�����` q©
�  ©�GdIdH`悥���Xd��  l��<i��Ī�<�:�<8�0�Ī��,�ɑ�O��ڲ��������)��


�� ����в �� w�`�Ī8�<��Ȫ��p��� �� ���ڲ��� k�������������8������ �� w˥G���
��𙩀�M�&e<i8�Ī�i��� q������
�I�i���  �������GdIdH�M���\��ڊ
��Ԫ��̪��ܪ��䪅�쪅�����Ԫ��̪��ܪ��䪅�쪅�����`�&i��'i� ��� ��	��� �����8��'` }�� 9թ��g���h�
�z�(�{��i��j� �k�����������d� �� �� � X�$h0�Lů$h*p+�j�k 5ְ ]̐�h	��h���x� �y�g���  �� <�L֮ �� �˥m�L%�d|��\��<����L����L�Lﮥo��n�,�p��	@��,�� �ͥmЭLz��_�] �ͥmО ��dh <� �� wˀ��g�]�o��n���	��� �ͥo��)�n��#,����G�� dΐ$}0�
���GdIdHL֮�_�] �ͥo���n��	�G�� �L֮$|0���|�g�]���^� �_ �� wˀ� �����L׮���(���)�b�x���)�A��R�h��d�)�F�\�f�p��q��m��rdndo,�p
����
�� �˩���s`�+ɑ�&��p� �q����i�p��q���m�r��sdndo`��m�i�p��q��s�rdodn�� Ͱ��o��n�$}0 4̀ ̩g�] �̀¥}��$}�	��\ez��)���\8��*���+��(��)d�d� �� w�`�+ɑ�e�*�+ k��G��,�0�
���GdIdH�4����.����3d�惭*,�0
8��*0�
i�*�(� �� wˀ���+������`���
�d��v�(� �)�'�+�&��i
�8�
�* �� �� 7��+ɑ��� �� ���E� �����FdGdIdH �� ���&����'�Y��*)�* }�L��+ɑ�L�悥����d��*�+ k�v�+�B��e��)��+8��+�	�+i�+�*0:��.�(�7�&��*8�&I���	�*�&���)��*�*��*�*�
�*��'�* �� wˀ���+� ���E	"�E��Z��[` 'ϩ�d 9թ�% M� 'Ϝd&�F�'���(��)�@�* �� j֢2 �Ϣ ����)���m�(�i �) 	� �� j֥<�$�� �d*��&�*�'�p�(��) j֢ �ϩq�(��) j֢ �ϩr�(��) j֢ �ϩs�(��) j֢ �� �� j� �� (۩��(��) �� j֢� �ϩ�� �� '멫� � '�$! ;�L ���������������������������������                                 " "

       $$$$$$$$���������(8HXhx(8HXhx � �                     �������H�ZH� 'Ϣ ���&�1��'�б�(��)�Q��* j��� �ߩ�&��'�h�(�) РZ�Ȣ �� �ܐ	���z���zz�h` '� 鲩�&�G�'���(��) Т� ��`�U�+d&d'�(��)� ��&�&���d&���'�Å(��)� ��&�&������+`�2�
�	 �� '� 鲩�&�+�'�u�(� �)�X Х&i�&��� �� �Щ�&��'�t�(� �) Щ�&�/����>�'�s�(� �) �Z� �*�ą(��)�
���������� �����&ȱ�'� jր�z�
�� �� �ܰ�ɿ��/I�/LU����`�2�
����� ���� M�LU���/`�.�C�`�}�����޴���PPPXX``hhppxx����PXX`hpx����PPPXX`hpx������PPPXX`hhpxx����PXX``hhhhhpx��PPPPPX`hhhhpxx����PPPXX`hhhhppxx����PPPPPX`hpx��PPPXX``hhhppxx����PPPXX``hhhhpxx���� 'ϩU�+�{�(��)d'd& Х&i
�&�(��'i(�'ɠ����+�|�(��)�0�'��&�@�* j� �Щ
�&�@�' �Ϣ �� �ܰ�`���ͶSUN WU KONG has saved his master but then enter the GOSSAMER CAVE. Here, he fights with the SPIDER DEMON.|They move on continuing their journey. They arrive at the FIERY MOUNTAINS and fight with the PRINCESS IRON FAN. SUN WU KONG steals the manfruit and then challenges the BULL DEMON KING to fight.|The pilgrims finally rise to the skies of Western Heaven. They go to the GREAT THUNDER MONASTERY and meets the TATHAGATA BUDDHA. Delighted by their arrival, he handles them the scriptures in which they will propagate in the East and eternally grant their great goodness. To congratulate them for their achievement of conquering and the completing the journey to the West, TATHAGATA BUDDHA also assigns them new posts: TANG SAN ZANG as the CANDANA-PUNYA BUDDHA, SUN WU KONG as the VICTORIOUS BUDDHA, ZHU BA as the ALTAR CLEANER and SHA SENG as the GOLDEN ARHAT.|H�Z�
�����#轛��$ 'Ϣ ���&�1��'�б�(��)�Q��* j��� �ߩ�'�  ����&�� H�� ̹h�:��$�0�'i	�'Ɏ��Z�Z�Ȣ �� �ܐ	���z���zz$�0�e#�#� e$�$��z�h`� d�d�Z�#�|�'� ��-��ڕ������z��� ��8eڨ`��i�`���نڀ�H�Z ��8� 
�� \Ͻ,���,��� � �ϥ�Z���z�0e�� e����� ���&�&�&�(�d&�e'�'ɠ�d'z�h`���������$�,�4�<�D�L�T�\�d�l�t�|�����������������Ļ̻Իܻ����������$�,�4�<�D�L�T�\�d�l�t�|�����������������ļ̼Լܼ����������$�,�4�<�D�L�T�\�d�l�t�|�����������������Ľ̽Խܽ�        ����� � 333     �c�c�c� ��0��� 46��f6 �c��3� ��`     ����� ����  c���c   ��灁       ���   �         �� ��`0 �7��v6� ������� �6��6� �6�6� ��c3� �0�6� �`0�66� �6���� �66�66� �66��  ��  ��  ��  �����`��   �  �  ���� �f� � �6���0� �c66�66 �gf�fg� �d000d� �gfffg� �d`�`d� �d`�``� �d007f� 666�666 Á����� �3� vfc��cv �````f� 6w��666 6v���76 �66666� �ff�``p �66��� �ff��cv �6p�6� 祁���� ffffff� fffffÁ 666���6 6c��c66 fffÁ�� �3��`6� ������� 0`�� �� ��f            ���       ��3� ```�ff�   �202� �33�   �3�0� �c`�``p   �33��p``�fff � �����  �33�p`fc�cf �������   3��66   �ffff   �fff�   �ff�`p  �33�  ��```   �0�� �����   3333�   fffÁ   66��c   3���3   333��  ��`� ����� ��� ��� ������  �     ��c666� �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I��HeJ�(d) ����M�dI�H�H�L�dHdG��I`H�Z y���:H�Z y��2�+ɑ�+��G�G��!�,���J��M��L  ��I����Nz�h`H�Z�+ɑ�&������(��)�$*��e&�*�'8��+z�h` ����  ����  ���� H�Z y��V�+ɑ�w�I�I��m�I����
���������m*�*�+8��+� B���+�;H�Z y��3�+ɑ�,��G�G��"�L�J��M��L  ��I����N y�� q�z�h`����H�������
��M��(�M��)�h`H�H��I��8h`  x{�H�Z����� �������ȹ����ɑ�X����C� ��r��,=��09��q�ɔ���0(���� k�����G������ m�����������L����� �� w� 5��
 ��z�h`H�Z��� �������ȹ����ɑ�)��m����m��� �~��~ȭi�ȩ���гz�h`H�Z��e&)��������i8�&�
-��04� 0���)��� ��,�*����(�"�����(� ����� �(� �������(�~����z�h`��	��`H y���+ɑ���( ���*)�*�&� ��� 	ѐ�����
��Ξ��&h`H�*	��* y���+ɑ���( ���&��	� �ѐ����
�����&h`HZ�'��00��' ���'��'��'8��'zh`HZ�'�p�h0�' ���'��'8��'i�'zh`�� ����� � ��������������� ��
���  � ��� � ������$����)�,�/�4�9�=�A�F����� � ���	
������      � � � � � � 666


$$$   LA�H�Z��� ��
����
����������ɀ��� ���ߨ����J����S����

��n��
�n���n���n��	�� ����� � 1���������ɀ�����m��� H�������ɀ�����m�����z�h`H�Z�������Ξ��z�h`H�Z��m8�&
I��
��ͬ��Kz�h`��m	8�'
I����ͭ���K�K��֜K8��H�Z�+i���*i����m8�
I��
��	��z�h`��m	8�8�
I�������8��H��I���h`  ��d 9թ&�,�X�\� �-�Y�]������I��i�K����`� � 7� � 89���(���(�������dQ����ή����0�Q
��V����V��� 5����'��i�&�(7��0�Q
��\��(�\��) j֥&i�&�(��0/�Q
��b��(�b��) j֮� �� �Э�8����Q�Q�ЃL�� k������������ ���Z���
�.�8��i ��� �� � 5�� k�z��ԥh	@�h <�`�Ύ�� ����H�Z��� �� ��������z�h` �� w˭�
��\����\��� 5� ��`��
 �� �� w� 5��
 �� �� wˈ��`� ����� �� w� 5�` ��% M� h����&�P�'������(d) ��dI�*)�*�J�� ���Ύ�� �� ���& �� 5� w� �� �ϥ&�
0��	��( ���ܢ ���N�� �ܰ	�� S����� y��g�+ɑ�`��( ���W��
H�*)�*h���H�*	��*h����� � 3��/�� ��� y��N�� ��N�� ?��N�� ���N �� )� À ��,J0; ��� �� �����+(�7L[� d��/�G���H�� ���L[� �� m�,J� ���! ���ILއ�N�05�N U���I���,��'��' �� w� 5�,MP� ��dIdHdG�ML7��� �� ���h)��h �� w˥*	�* 5�)�* �� �� wˢ� �� 'ϩ �% Mݩ�&��'��(��) '� �Р ����&�х(� �)� ����&��'��(��)� ���� �ϩˢ� '�LB�H���#�
����I	����h��Ί���
�(�����������=����� 5�h`H�+��$*�&i� ��&�0��h`H�Z�/ɑ�9�(�4��(�.m~�.�*�)��.�/ k� m����/ �� w� �z�h`H�Z�/ɑ�=�,�� m��.��i�/���~����8�&��~���(�
�)z�h`H��8�&��)���	���h`H ���,�0�����h`H,����		H�E� �S�-�N��-�*�D�&8��I��06���)����*����*����*���*�+��,h`���0�� 楠����*��H�&8��I��8h`��Ƌʋҋڋ����؋����������������������������}~����������������    ��H�Z�,�L���*����,�*�� )����+,������m����9�	�,����+���&�� ����� ���� ������/���R�*
�����轨���+
����ȱ������+�*�	 �� w� �z�h`�.)�.�*��
 ����*��*�+L,�H�*���	�$��+������ D�,.0�.	��.8�h`H���� ���*M����,.p�.	@�.��-8�	�.)��.h`H�Z��:8�&	I����
ͬ�z�h`��i8�8�'	I����ͭ��8��  ���� 9թ��,��-���X��Y��Z�
�[���\��]��^��_�>�������������������(������/��i��������o���(�������*�+�
����������z� �{`H�&��0 	�����&h`H�&��	 ������&h`,� P�� 9�`̶�H�Z�(����*�+��,�
 	�������&�� $EP���'�
 ��ڢ
 ��� ���&���P� �� �������'�'�'�
�&� ��Ȣ�'i�'�& ����� �Ʃ2�-z�h`ڹs��( �� w˩�� 扢 ���` �� 9ե% M� y��h	@�h <۩(���
�[��_���� �ȥG� �!,/�/�̢� '� 9ե% MݥE)��E�� ��I�� 所 ���� �� �����- � � ފ L�,J0i �� ��}����� �� w� � ���"L$� 猐 e� e� e��-i
�- m�,J0',MP�$EP���(dVdW �� w� 扩 ���ML.���G� ���$EP�� ���E�@�㩀�/�ܢd �ϩ~�� ��dGdIdH �� 扠�(�� �ϭ������� �� w� 扈��*)�* ���d �� 'ϩ��(��)�
�&�<�'�
�& �� j֢2 �ψ��͢�$EP�΢� '�L#� �� Т2 �� �Т �ψ�� � ��`�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������d �d�ʢ�  '� 9ե% Mݩa��� �����(��)����������������������� �� p� B� w� ���E�&���'�Y��*)�* }�� 9թ��X��Y��Z�
�[���\��]��^��_������g���h�	�z�$�{�
�i��j� �kd������������}��\�h	��h���k�O�  �� <� �� � t� ��$g0�G�� gĥ*)�* ���&�� 	��& �� wˢ �π�@�g���h��z�$�{��i�<�j� �k����������� �� � Q� ��$gp�&���'�Y��*)�* }��Lj�$h%p&�j�k 5ְ ]̐�h	��h���k�O�  �� <�LW�,�0�	�z�$�{�Q�x� �y�O� �k���z��{�[�x� �y�W� �q�t�u�] �� �˥m�L��d|��Lr���Ly�����4��ML�����o��n�,�p��	@��,�� �ͥm�LW�L� �ͥm� ��dhdg <ۜ� �� w�LW��o��n���	��� �ͥo��4�n,�0��)���#,����G�� dΐ$}0�
���GdIdHLW�$|0���|�t�^�u�_ �� w�LU��~���2��� �����LX����.�~�
�¥)Jj��,�0�O� ��W� �p�q��r��s��L���2�����>�)Jj��,�p
����
�� �˩���s,�0��T� ���W� �r�p�q��mdodnd~`��m�O�p� �q��s��rdodn�� Ͱ�ޥo�$}0 4̀ � �̀ɥE	�E�N�O� �ϥo�,�n� ��a�
���`��Z�]i^�^� i �_ �� wˀ��do�n�n��0dn�,�o�o��$�n���  �ܩ��� �ܥO��P�
��GdIdH�5 �ܰ����O��O�O���OL���O���O� ���N�N���dmdodn�E)��ELW�$h*p+�j�k 5ְ ]̐�h	��h�z�x� �y�k��� �� <�L�� �� �˩k�]�m�L7�d|��L���L�����,�D�o��n�,�p��	@��,�� �ͥmЭ ��L�� �ͥm� ��dhdg <� �� w�L���o��n���	��� �ͥo��)�n��#,����G�� dΐ$}0�
���GdIdHL���o��ni��^� i�_ �� w�L���n�����L��do�nI�n$}0 4̀ � �����o���3��m���p� �q,�p
����
�� �˩���s��rdodn��o`�\8�&I�8�z�8����)���m���p� �q��s��rdodn�ǩ�m���p��q��s��rdodn�� Ͱဦ�o�E$}0 4� 4� 4̀	 � � ̥n��c�"���W����H����O�
���e��i�] �ͥo��	�n��L�L���~
���~-Hڥ=�@ ۩@�*���k��(�k��)�k��'�k��8�<�(	��0�& j֭��� (��h`()* /01234H�Z�=�)�<e&�G��� ������	������ �ɞ������8z�h`	Hڥ�E��A�=�=�<e&i�3�-�8�-����8�� �	�
�8�
�����i�8�'���'�h`L�H�Z�O����O�+ɑ���)���(�����(�*���G�r�'�Y�l�(�*�'i�g�J�+� ���*�+���K k�K��:��( �� w� w�,�0(����� ���΢� �ܥO��P�
��GdIdH�� �� �� gĀ����+z�h`�*�*�* �� wˀ�H$g�<e&�@�8�h`�� �d 9ե% Mݩ��g���h��z�$�{��i������������������� �� ٠ �� ���g)��� �����g���h��z�
�{���� �� k� �� �� ���&���'�Y��*)�* }��L�$h@pA��j8�<�(���:�j8�<�($��0 �\�h	��h�C�x��y�R���I� �� <�L�� �̭��]�m�fd|�m����$��L��L(� �ͥm�� ��dhdg <� �� w�L����8��]�o��n���	��� �ͥo���n��,��� A�L�� ��$|0���|�H�~�~��.�+ɑ�'�����!�����F�p��q��s��r��mdndo�$�d� d~�L�c� t��d~�I�^��_ �� w�`�o��n�,�p��	@��,�� �ͥm��L���L�� �ͥm��,L0-���L���)��d�8�<i(�\�l����d� t� ����L�� R6R!R.R<�p�q��s��r��mdndo`d}�\0�&����}`�+ɑ�+�*�+ k�&�G�� dIdH�
,K�G�����+����`����������Vd�惭I��I�����+i�+���1���+8��+�����*,K08��i�* �� w�`�`�+i�+��$}0�\8�&8��
�&8�\8���]8�'0%�
�J� ��\i�*�]�+����S����9I���"� ��\i�*�]i$�+����(����]i�+�����]�+�\$}ez�*�}�K��(� �)�d�d�`#-7A<72-(#

##-2A<-
(2<A7-#

#-7A7(
(2A2((2<A7(###(<A<7((2A77-##7AA<-$hp-�ąh��i�'�\��]���^��_dmdodnd}�� <�L��m�$dh�%��� ���]���\���O �� w�L"��~�~�����I��i��^� i�_�\�\������)����룍]�A��
� #������� #����d~ �� w�`�  T��ɑ�+�\i��]i
��Ғ�� �� ��=���d������`8`*.Z^��+/[_��(,X\�� ������L0�悥��
��d��  T��ɑ�oڲ��� k���1�]���,�0`��o��i��:����:�<����/�1�G��+�
�'��#�&i8��
���GdIdH���\� �������Ѓ �� w�`��o���i���&��:������(�π�ڊ
��n���b���z�������n���b���z�������`��ɑ�L"��O�O�
��O�������������� k������@���B��e��)���8����	��i�����
�����)�Ί�������� ���ЅO��P <� �� w�`�� �d 9� )� 9ե% Mݩ!�_��^�Z���[������g���h��z� �{��i��j� �k����������� �� �� K� ���g)���&���'�Y��*)�*L��$hXpY�j�k 5ְ ]̐H�h	��h$g�P�t��u�L�v��w�J�x��y��Y�t��u�U�v��w�S�x��y�o�t�u �� <�L�� �� �˩o�]�m��1�o��n�,�p��	@��,�� �ͥm�� �����LK�L����: �ͥm�0 ��dh <�$g���h��z� �{��i��j� �k�dhFg �� w�L����U�k�]�o��n���	��� �ͥo��4�n��.,�)���G�� ,��� �� dΐ$}0�
���GdIdHL����L���o��net�^� eu�_ �� w�L���n�����L��do�nI�n�)��\8�&�\0�!� ������\���� 4���� �����C���>��m�v�p�w�q,�p
�������������G������s��rdodn��o`��m�t�p�u�q��s��rdodn�� Ͱ�,�p�0��� }� ��� 9� q��O���g���h��z� �{��i��j� �k����������� �� �� �� �� ���g� �멀�g���h��z�$�{��i�&�j� �k��������d� �� \� �� �� �� ��$h0�&���'�Y�ީϢ� '��L}�$h*p+�j�k 5ְ ]̐�h	��h�;�x��y�k��� �� <�L^� �� �˥m�La�d|��$��L��!��LK���Y��Ly��	�L�L�� �̀��o��n�,�p��	@��,�� �ͥmНLF� �ͥmГ�k�] ��dh <� �� wˀR�o�6�n����p��q��s��r�W����M�������� V��\��k�] �̀�o�$} ̀ 4� ��L^��k�]$|0���|���^��_ �� wˀ�8�\�&I��z����}�i�z�`L_�ͬ�d}�
iͬ�ML_����)�)��yL^���G��)�\�h����)�j�L)��z����� V�� �p��q���W���p��q�
�m��rdndo,�p
����
�� �˩���s`���p��q������p��q������p��q�	��m�r��sdndo`��m���p��q��s��rdodn�� Ͱ�ޥo�I�n�
��	����;���W�0���M�(���\$}08��i�\�\��k�]�o ���o��] �ͥo��C�n��=,�8���G��/��z dΩ�z�"$}0 q� q� q©
�  �  �  ©�GdIdHL^��o�$�n�
��	�������\$}08��i�\ �ͥo��̥n���Lܬ�}���\$}ez�*�]i�+�&�(� �)d�d�`�+ɑ�e�*�+ k��G��,�0�
���GdIdH�4����.����3d�惭*,�0
8��*0�
i�*�(� �� wˀ���+������`~xvx~���`ZXZ`fhf�O�O�� ���LϮLЮ�O�/ɑ�Ll��&���)���K�'��	����K���.� �)���������/����,��-Lɮ ���_��)�����������/�)i��,� i�-,K0�.�.�.������.�.�.0	�(����/ �� w�`�G����
�����,K0�
���GdIdH���\�ϭ��������
��.�/ k�����`�������������������������������� " "

       $$$$$$$$���������(8HXhx(8HXhx � �                     �������H�ZH� 'Ϣ �a��&����'�!��(�A��)����* j��� �ߩ�&��'�h�(�) РZ�Ȣ �� �ܐ	���z���zz�h` '� :���&�G�'�Ѕ(��) Т� ��`�U�+d&d'�х(��)� ��&�&���d&���'�҅(��)� ��&�&������+`�2�
�	 �� '� :���&�+�'���(��)�X Х&i�&��� �� �Щ�&��'���(��) Щ�&�/����>�'���(��) �Z� �*�Ӆ(��)�
��J���J��� �����&ȱ�'� jր�z�
�� �� �ܰ�ɿ��/I�/L�����`�2�
����� ���� M�L����/`^������α��/�F�i�PPPXX``hhppxx����PXX`hpx����PPPXX`hpx������PPPXX`hhpxx����PXX``hhhhhpx��PPPPPX`hhhhpxx����PPPXX`hhhhppxx����PPPPPX`hpx��PPPXX``hhhppxx����PPPXX``hhhhpxx����d* '� �Щ2�'�@�*��������'�&�# ޳�	 M� �����$"Ls����$"PL�� �Щ�������'�&� ޳�	 M� �Щ�������'�&� ޳�	 Mݢ< �� '�d&�!�'d*���(��) j֩
 M� ��d����P �Х ��� ��� �� ������
�� M݈�� '�d&��'�ԅ(��)�(�* j� '� :��O��P��4� ��� ���
 �������� ��`HZ �d&�' �נ � ���(�� (�zh`HZ �d&�' �ץ��8�>�� ����(�� (�zh` �Э��(���) j֢ ���&���`H�&�
�'�� �&���'�A ���= ��hH)�JJJJ ��hH) ���  ���X ���= ���)�JJJJ ���) ���  ���Y ���= ���)�JJJJ ���) ���  ���	)�JJJJ ���	) ���)�JJJJ ���) ���
�&��' �ܰ�h`�
�i0�i7 ��`H�Z ��8� 
�� \Ͻ������ � �ϥ�Z���z�0e�� e����� ���&�&�&�(�d&�e'�'ɠ�d'z�h`Եܵ����������$�,�4�<�D�L�T�\�d�l�t�|�����������������Ķ̶Զܶ����������$�,�4�<�D�L�T�\�d�l�t�|�����������������ķ̷Էܷ����������$�,�4�<�D�L�T�\�d�l�t�|�����������������ĸ̸        ����� � 333     �c�c�c� ��0��� 46��f6 �c��3� ��`     ����� ����  c���c   ��灁       ���   �         �� ��`0 �7��v6� ������� �6��6� �6�6� ��c3� �0�6� �`0�66� �6���� �66�66� �66��  ��  ��  ��  �����`��   �  �  ���� �f� � �6���0� �c66�66 �gf�fg� �d000d� �gfffg� �d`�`d� �d`�``� �d007f� 666�666 Á����� �3� vfc��cv �````f� 6w��666 6v���76 �66666� �ff�``p �66��� �ff��cv �6p�6� 祁���� ffffff� fffffÁ 666���6 6c��c66 fffÁ�� �3��`6� ������� 0`�� �� ��f            ���       ��3� ```�ff�   �202� �33�   �3�0� �c`�``p   �33��p``�fff � �����  �33�p`fc�cf �������   3��66   �ffff   �fff�   �ff�`p  �33�  ��```   �0�� �����   3333�   fffÁ   66��c   3���3   333��  ��`� ����� ��� ��� ������  �     ��c666� อ�s�����E�SHU WU KONG goes into the Peach Orchid and jumps up onto the trees to collect the Golden-Hooped Compliant Rod. He passes the EAGLE'S SORROW GORGE and meets the GREAT WHITE DRAGON in which he has to fight.|SHU WU KONG defeats the GREAT WHITE DRAGON. A GOLD HEADED PROTECTOR appears and turns the dragon into a white horse to serve as PRIEST TANG SAN ZANG's mount for the rest of hid journey to the West.|When ZHU BA JIE loses, SHU WU KONG will replace him.|SUN WU KONG has defected SHA SENG and convinces him to become the third disciple of PRIEST TANG SAN ZANG and to follow them on their journey. The four of them then arrive at the Seven-Storey-High Temple in which monks plead for their help. Their treasures have been stolen and they will need to go to the DRAGON PALACE to retrieve it.|ZHU BA JIE has defected SHA SENG and convinces him to become the third disciple of PRIEST TANG SAN ZANG and to follow them on their journey. The four of them then arrive at the Seven-Storey-High Temple in which monks plead for their help. Their treasures have been stolen and they will need to go to the DRAGON PALACE to retrieve it.|SUN WU KONG defeats the DRAGON KING and collects back the treasures. They continue their journey and pass through the WHITE BONE DEMON'S CAVE in which PRIEST TANG SAN ZANG is captured by evil spirits. SUN WU KONG goes and rescues his master.|H�Z�
��Ը�#�Ը�$ 'Ϣ �a��&����'�!��(�A��)����* j��� �ߩ�'�  ɾ��&�� H�� ��h�:��$�0�'i	�'Ɏ��Z�Z�Ȣ �� �ܐ	���z���zz$�0�e#�#� e$�$��z�h`� d�d�Z�#�|�'� ��-��ڕ������z��� ��8eڨ`��i�`���نڀ�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xآ�����  � � � �  �Μ" ��& d d� � � � �������X�� Dϩ��+��X��N �ܰ������" b�����@�" �����!� �% M�L �� �% M� ��d���� �L ���LB�L#� ȩ� Dϥ��L����L �L[�� �� �ܰ����� S�Le����������$E�E����B�	�>�����6�����.�����&�������������Q��M���G�'�Y�A��G�2��������*������������������GdIdHdQ`����� ��L��L��H�$EPi�$Fi�	���i�S�h`�I� �H�$E0� ����#�� |���SL��LJĥI�� �� ��  ¥��	� 1���&�@�*�H��$E0����ȩ$�ĩ |����Iо �� �� q¥��	� 1���&����$Q`���� ٞ�:��� .��0����	�� Ǣ��&m��)��&�� 	ѐ
$hP 4�`�&��$Q04���� ٞ�'����	�� Ǣ��&��� �ѐ
$hP �`�&���I�$Fpn�H� q�$\0 d\�*	@)��*� |� �åI��9�E� �0������� �܀ ������ �ܥO��P�
��GdIdH�� �� ��`�Iй�Hе  �$\0����H��"�S �åG��F)��F��`�I�$Ep
�H��
��  �  ©@�*�/LJĥI��$Ep
�H��
�� q� q©��*���d۩�M�I��$EpK�H�� |��>���������I�e'd'0�' 4Ɛ���ۀ�����R ��dR��� �ƀ�H�� |������������I�U�S
���ȅ��ȅ�H

eH���W�(d)ȱ�M�$*ȱ�V�$*0ȱ�W�G��
���	ȱ����Q �� wˀ�M�dI�H�G���� �����`�I`dGdIdHdQ`�I�֥H�� |���� ��L�åI�C�H�� |��8��-�����*��&�����R ��dR�8�Y�'JI�eY�'��� �� �åI��	�H�� ��`�I��H�	�$F:�S �åI��6�H��0���+�+ɑ�#����(��)�&8��*�'8��+�E)?�E`�/ɑ���X���,��-�&$*0i�.�)���'8�0�/�I�O��8��.�	��I��H�	� $EP�S �åG��'�Y��' ��`�I��H�� |������� �� �åG�2����� A�� ���N�L��ЅO��P <ۥE	"�E��Z��[`H�Z���4� �0�=�,�<e&�%�@�!ɨ��'�S�*
�&i��'i� W��'��z�h`H�Z��=��9�=�5�<�7�/ɓ�+e&ɨ�$� �'�"� ���'�Z �� w�z���8z�h`� �����&$*0i�i��'i � ��3�'�Y�-�'�R$R�R)���R)��R��')��� �� wˢ �π�`H�Z���� �1�=�-�<e&�&�@�"ɪ��Z��,��� �(��� �)��� �9�Y�'$R8��'�� �z�h`$R0	 ����$R�'i�Y��Y�'�� ᡀ� {ƀ�$R0ҥ'�D� ���'��' �� wˢ �π�'�Y��'�')�� �� w� wˢ �ϥ<e&ɞ���L���*
�&i��'i� WL�	59b	=H� '� ۩ �*��(��)d&d' j֥
���ǅ&车ǅ'�����i�(� i�) j֢ �� �ܰ���ɿ�����дd�� (��h`H�Z�%� �� �% Mݥ*H� �* 'Ϡ��(��)d&d' j֢ �ϥ
���ǅ&车ǅ'�����i�(� i�) j֢ �ψ��h�*z�h`�E��*�Z�& �� w˥EI�E���
�Z���Z�[��E)܅EdZ` |ȥG

i� iȅl  ��` ��`  �` {�` <�` ]�` ��` ��` p�` ��` ��` �` y�`@�V�K�f�vɟɯɿ��������� �� �+�1�<�L�uʅʕʠʦʱ�������
���+�;�A�G�\�g��  �   ������ �     �   �  	 � 
��  �  �  �  �� � ���  �   �  � ���� �  � � ��           ��  ��   � � � � � �  � � ��� ��� � �  �  �� � � �  ����� ��� �  � � � �  � �  ������� d���e���f��� g� �h� �i���j���k���l���m� �m� � ������������ ����������� �������� ���� )���*��� .�  / � 0��  1�  2�  3�  4��5 � 6��7�  7�   8�  9� �:��� =�  >� �? �� ;   <   ;    G���H���I��� @� �A���B    �   � �  C���D���E���F  � ��  ��   +�  ,   -�   �E���&�TeV�&�'�UeW�' j֥T�&�U�'`�G����/,�P*�
,�0
 	��&�\� ���&�\ �� wˢ �ψ�ۜ�`�\8�&I�8�zI��8�I��� �ʀ��� 4�ʀ�`�\�(�&�\�\�(��8�( �ϥ<i����jdk�h)��h`�\ez� �\�\ez��<8�dj��jdk�h)��h`�h� �7�\�(�ɀ� 4̭\�'�"� ��\ez� ̭\ez�����}8�`�]�^�_dmdodn����d|�h� �)߅h�*)�	@��`�h��-�m����#���hI�h�� ��ƀ��h)��h� �� w�`��hI@�h �� wˢ �ψ��d ��` �ͥm�$�o��F$}0 4� 4� 4̀	 � � �$hP,�($}0�\8ez�&����&m��\��}I��}�8�`�h	@�h$}0�\��'�\�}I��}�߭\8�&���}I��z�i�z��d}ͬ�iͬ������� `�o��nep�^� eq�_ �� wˀ�s�do�n�n�r�dndm��o`$hsPq�m��k��g�\�] ��\ �� V� d� ݩ ���i <ۥi��i���h	�h��������������������m�s�r�x�p�y�qdodn`�\8�&$}3I��z��*�$}0$ͬ���]8�'I��{���ͭ��8�`�����$* 4̀ �`H�$h#P!�h�� ۢ �\�&�����}	@�* j� (��h`H�G�
�m� �� w�h`� � � � � � � � �ҍ � �( �) �* ��f`H�Zd �@�� � � � �������z�h`HڪJ)�! �Jjjj) 	�& �h`Hڪ)��)���J)�! ���� Dϩ ��h`H�$J)�! � D�h`ڢ(ڢ������������`HZ�dd
� �ψ�zh`HZ��d��&����e��e�zh`HZdd�
&&(&&���%+��%+�zh`H�Z �� ��F,�-� d.�,�0�  ��Z�.��ȥ��.�.z��0�� [���� ��z�h`H�(e � � e��0e�� e�h`H�,��H�Zd�� �ע�� � ���(�� >���� ��z�h` �� �� ��`H� ��	 �
 � � ��� � � ��	 �
 �� ��� ��� � h`H� ��	 �
 �@� � ��� � � ��	 �
 �P� ��� ��� � h`H�Z�:��6�8�K�6 �$D�;�	�6�:�6 � {�8���;� dѦ;�
�7 � d��7 #��:�:�(�d:��68z�h ��(`���������(���Z�:$D0� �� z� >����`H�Z�:��6�C�6 �$D�;��6�2�'�:��: � {�8���;� �Ѧ;�
�7 � ���7 *�8z�h ��(`���&�ȑ�������Z�:$D0� �� z� >����`H�Z�;�
�7�j���;�7�;�;�;�; ԩ�������ڢ(��������8��X��� ����� {� A��'�'�'�'�:��6 � {� i��68�>��>�?� �?z�h ��`�(�; ���e � �e�d��`H�Z�;��7�9�rɌ�
�;�;�;�;�d;�7 �d������ڢ(���������i��i ����� � A��'�'�'�'�:��6 � � i��6�e>�>� e?�?�;��7z�h ��`�;������ʩ( ���e � �e��@���`�8�'�
�:�$D0Z�
� z�� ��
����� >����`�8�'�
�:�$D0� �� Z�
�z�
����� >����`��� �y � � �   K x � �  K �� � � � � � � � � � �( b c } ~ � � � #$� � � � � � � � ��L)��LW��Lg��Lw��L���L���L��H�Z�6
�dD�

i�� iӅl ���7����Ӏ���Ӏ�����Ӏ�7����Ӏ���Ӏh�����Ӏ^���ӀX�����ӀN�âӀH�7��ǢӀ>���͢Ӏ4�ӢӀ.���٢Ӏ$�ߢӀ����Ӏ����Ӏ
��Ӏ��Ӆ�	��4ȱ�5������D��(�)�4�(�5�) �׆(�)z�h`                                                        H�Z�� ���e

����ԅ��8ȱ�9ȱ�6ȱ�7d:d; �$D0 �ϥ4�(�5�) aХ����X���Т�O�P <�d<d=d>d?d@dAdBdCd&�@�*����� �
��������E� ���������F����� ���o�
�V����q�����Y�' g�dhdmdodn ������J�����%z�h`�<��=`H�<��=�<h`�Z�<��=�����<��=�$*0d}�'����}�zI���\8��z`H�Z�&�-�'�. ��$*0d.��,:�.�*) �Lץ'�ɐ#I��-�T�, ���e � �e��-e'�d'�ɐ�4e-ɑ���8�'���-�&#$*0I���,m-:�.d&�,m-�0� L���(��e,�)�$*�,�.�.�(8�&��,�0�$*0d.��,�.�.�,�0�- �ץ*���8�>��.�/�0�1�/�.�1�0� Z�.� z$*0�.�ڪ����.�$*P)��*������)�� �)��)���)���=�ّ���0д [��Ф �ϭ-�&�.�'z�h`Hک0�' ���&e��@e��h`HZ�(�2�)�32&3� e2�2��e3�3�(e2�2�)e3�3� �2� ȱ2�ȱ2 \ϲ �-� ��� �,� ��zh`         0300<?<<03000300                  ����������������������������������������������������������������         0300<?<<03000300                           0300<?<<03000300                      
    
  "#  "#((*+,,./0023002388:;<<>?    
    
  "#  "#((*+,,./0023002388:;<<>?�������������������������������������������������������������������������������������������������������������������������������� @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��Hڢ �&�(�����h`Hڢ �(�&�����h`���H�Zd�[�� �� ���(�� >���� ۥ���%� ��J� �(�)d&�`�*� �9ۅ' j��&�&��N��O��PJfJfJfJf��x��x�[��f������ �0��ڢ� >�������������ʀ����?���������� >����$hP^�h��X�$�&���'����b���ɢ �(�) j֩\��Ӆ�����i� �#��ʩ���ʩ��� >Ј��������� (�z�h`H�eO�O�eP�P����O�А�ЅO��P <��h`H�eO�O�eP�PdOdP <��h`ڭ  ���$]0�����  ������]�d]8�`H�adb���ch`H�Z�c2�a
��݅d�݅e�b
eb��d��* ȱd�( ȱd�) �b�dc�* z�h`dc�* `��,�3�C�
/
 ?O_O �� `�o((�(� /X� H�Zd�d�


��腍�腎�腜�腝�腔�腣�腓�腢���������������Ȅ�d� V� �ޥ�	������������������Ȅ�d� �� (ߥ�	@������� � ����z�h`H�Z��)���$����d���	�� ��春�ŗ� V�$�P���d���	�� (�槥�Ŧ� �ޥ�������� � ����� � �ҍ � ��� ��)� z�h`������ȱ���ȱ���Ȅ�d�d���)
��M酙�M酚���%������ȱ�������$�Pd��� V߀Ȅ�d���`������ȱ���ȱ���Ȅ�d�d���)
��M酨�M酩���%������ȱ�������$�Pd��� d߀Ȅ�d���`��)?	@��$�!��)�������)���Ȅ������ƛ��d�`��)?	@��$�!��)�������)���Ȅ������ƪ��d�`H� d���)��h`H� d���)���h` ~    � � � � ~    ^ c i p v ~ � � � � � � � . 1 4 7 ; > B F J O S X ^   Y�Y�    ^ c > c   ��    ~ p c   �Q �    � c ~ � � � �    �    � �    ���         � � � ~ � � � � � �$     � � � ~ � � � � i c$  c    c S X p c c X c$  ~ ~ c ~ � � � � �$     � � � ~ ~ �  � �   �Qe, �e,>�Qe�Qe, �   e,>�Qe�Qe�Qe�Qe�Qe   �Qe�Qe�Qe�Qe, �, �    � ��Qe�Qe, �, �, �   > � � �> � � � �> � � � � � � � � }> �}>ez�	z����z��> � � �> � � � � � �> � � � � � � �� � � �> ~ � �z � � � �� �   � � � �> � � �> � � � �> � � � � �� � � �> �> �� � � � � � �� � � � � �� � � � �>� � ~ � � � � � � � � �> � � � > � � � �    � � � v> � � � >& � � �7>e>�e}e> } > � � �> � � � �> � � � � � � � � � � � � � � � � � � �    � � > � � � � � � � � � � � � � � � � � � � v> � � �> � � �    >>>>> � � �>>eeeeze>>  >>>>>> � � � � �>>eeee   z���z> ��zz��ee  �������zz>��zzzzz���eeeeezzzz������    �@�@�@�@	�`  �@�@�@�@�`  � � � � �@�@    �� �� ���>�z�z   e�� �� ���>�z�z   e�� �� ���>�z�z   e�� �� e�z�z��z�z   e�� �� e�z�z��z��    �    �  ���      �   � � �   ��  ���   �  �����}�  ���   �   � � ��  ���   �   ��� ���}  }}} �   �}   ��� ��   ��觧DD���误    ##DD    �����觧���觧���觧���觧���觧���迿����??���迿���觧��駧DD+�+鯯DD1�1駧DD=�=�//A�A�//E�E�//I�A�//P�t�����  ��1�j��  ��  r�  x�  ��  ��  ��  ��  ��  �  �  �5�5�h������5�5�5�h������  �5�5�h��"�@�X�"�@���  ��-�  ������@�  /�  5�  >�  J�  [�^�i��������
	�		�
�

		�		�		 �d*��X�D�Y�(�Z�b�[ 3��X�Z�Z����X�Z� �� 3��[�[�C��
 Mݩ \ϩ��  f꩐ f� �Ϣ� ��` 'ϭX�&�Y�'���(��) j֭Z�&�[�'���(��) j֢ ��`Hڜ � � �� ���� $0�� � ���h` V� d� ��X���/��/��� u�� $��/���� �� ʲ���L7������N�ЅO��P�� �ϥ
ei�� i�������% M�l �v�j�K�� �,��� ��� � � �_� �[�۬�H�%�� �% M�hZ��z� ¯��� 7��
 q���� ��`�* � � ��� �`H$0(����� I�)�� ���ƌ �ݥf��f� �ܩ�fh@Hڭ' ��	���$ �d�% �� �� �ܰ����d�hX@ 'ϩ� ��dd� �� Dϩ��d � � e�� e������� ����������d ��L���&�P�'���� �� ��Z�'������� ��#ȱ�$�8�#��� ��8�$��� ��$���#����&�O ���K ������&�F ���A ���I ���L ����CHECK SUM��F�'�
�&� ������ ����`ZH)�JJJJ ��hH) ��hz`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ������H�x������8�h�������(�X��������H�x������8�h����Ъ`*.Z^����+/[_����(,X\����H�Z �� "� ۩�������-���-��@�*����*��y��y�� ��� ��(ȱ�)������,����,�� .��.���О����	�� ���� ������ 1� (�z�h`H�&����'��	,�$  j�h`H�Z ��)�� �$�#H�Z ��)�ɀ��)0� ��)���)��z�h`8��H�Z ��)�����)0�0��)���)��z�h`8��H�Z ��)���)0��)�
�)�z�h`8���d���&����.����m��m����e��`T RV (V��X��f >h��p��r��y >�  �����Ș F� (����������� nLO�H�Z����=��$ p� 	@�  �� w˥(H�)H�*H���������%�(������������8�<�(c��0_��8�>���?���	�ɏ�?����9����2����������60����������� S� k� ���.�.���9�Lx�h�*h�)h�(,�0.$ 0��ɑ�I������ k�� ���E	��E��	���z�h`�Z��,��'��,����,���&H�'H�&�'$  j�h�'h�&z�`�i��Y��i��Y��`��������������������������� ���R�  ^�`�@�<�@8�<�= I��*�.�Z�^ΊΎκξ:���*�.�Z�^����:��`d�B�>�B�>�,��� �i��i����� [�� c�����`ɑ�8�`ɑ�i`H�Z�:8�&
I����
ͬ�z�h`�8�'
I����ͭ��8�������	�H�Z�G����e�H��_��H��WڥG����� $EPi
�����轡���$*0����轡�e&��轡�e'����8��	I��z��
���z�h`�8��	I��{������8��H�Z�8�&
I�����
ͬ�z�h`�m�8�'
I�����ͭ��8��(�� |�dH�S
���ȅ��ȅ�H

eH���(d)��$*ȱ�V�$*0ȱ�W �� w��&� �ϥ&)���Z�^�H�H��&�0�`���X��Y��Z�
�[���\��]��^��_ ��߅( a�`qppq���    '� ����&�q�'� �
 �Ϝ���&��'�!�(�%�) �� j֢ ������� �Т� ��` uuy\]^_ �� �ϩ����'��&�
����(轁�) �� j֢ �������� }��( aЩ �&dVdW��'�  I�� �ϥ'8��'��&� I�Ȣ�'i
�'�& I���� �Ʃ ���y�&�}�'�!�(�%�) �� wˢ ���(����� �Т2 ��`ڹs��( �� wˢ �ϥ&)���Z�^�`LӇHڥ���M�
�����
��������� �ܥO� � �P� ����J�[�+ɑ����[ ���h`��������+ɑ��#��!�(d) ���M	@�M��N��H�Z��4�!� �[0�#� �(�)� �� �� w� 5��2 ���(���dG��I �ŀ�J��GdIdHdQ�J�Nz�h`H�&�(�'�)�(�*�)�+�*�,)��*���&���'���(���) j֭(�&�)�'�*�(�+�)�,�*h`� ���i <ۥi��i`8`H�ZHd�� ����t�����t�����h Mݥ������% M�d�� ������������ V� �� �� (ߥ�	���z�h`H���+�/�[�_������������h`H�*)��*���&���'���(���) j�h`H,y!�*)L�*�H�&�I�'�J�(��K�) j�h`     �� ������   ���� ��  ��      �� ��     ������L ��    M ����  N       !   ����"   �� � ������#   ��  $   ��  Hڜ�


��Z����Z���譊�(�%���)�$*��Z��V��Z��W�h`�Z��V������H���&����Z�Z���(�Z�^�^�^���(�^h`H����(���mZ�^�������h`�`�X��Y�a�\��]��Z��^��[�_��`H���%���Z ���Z�^ ���^�X��\�X��\�h`�)���(`��`������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ � �� V� *� d� �� r� (� �� � :� �� Z�  � � �� n� 0� � �� s� o� %� ì � � � K� �� t� x� z� ۹ � K� �� `� 4� F� L�  �������ʙ��T�d���ޞ��x�>� �Ƣ��\�ڥ˧ǩ}��I�E�A�=�O��'�I�K��O�a��� ���Η�Й�\��T����&�ؤ2���"�����l��j�Ϻ�� �������α�Z��V�޸p�Ȼ�� �X���ż���Ž� ������� ����e�Ư��>�h�"�d���z� ���������ʸ ������f��,�����4�f� �������d�ʸ0� �	��	�	n�	z�	��	��	��	��	 �
��
�
�
Ȯ
�
�
�
Ĳ
Ƴ
ȴ
��
��
��
p�
R�
4�
 ����7�j���еV��A��Y��� ������$��~�ܽ ����Ү��n�<�
�ط0���� ����x��`�Ժ� ����Ү*���ĵ�H���4�޽ ����J�8�e�|� ����\����N���Һ��T��� ������ȴ��M� ����į������� ���̍����������±³µu����� ����������ʰ����������������й������ ���
�~�#�E�g�A���9���9���9�[�}���1�s�ݟ���â��������Ǩ��������ͭ�Y�[�]�_�	���-�o����A���͸ ���$�ބp�ĈҋX�ޒϔ����t�N�(���������̫��p� �ڀ������������������~�|�z�x�v���ʕ��0�R�t��$�F�h���L�z���v�D���ɫ�����׬��ʻ޻����޼� ����L��� �������Z���޸ ������ΰ�R���ܽ^�w��� ���ƀR���΁�r���֖(�z����.�@��������������������������������������������������������������������������������������������������������������������������E|c� ���