                                                           �?      p�      \�     l�     l�     ��     ��    �<��   ���?    Ϫ�;    ����    p���    p��?    ���     ��     ��?     ��>     ��     ��;     W~9     \s     �s     ��     �s9     ��?                                             �     �e>     p�     p�     ��     ��     ��      ��  �  ���  ��_50  ��[90  ����0  ���  �kU��  ����    ����    ����    ���z    ��C    �     \~     �_     �     ��     �o     W�9     ��?                                              �     �e>     p�     p�     ��     ��     ��      ��  �  ���  ��_50  ��[90  ����0  ���  �kU��  ����    ����    ����    ���z    ��C    �     \~    �_�    ��    ��    �o�    W�9     ��?                                              �?      ��     �e>     ��?     ��7      �      �     ��  �  ��   ���0  ���50  ��[�0  ���  �kU��  ����    ���    ����    ��     ��}    �N�   \~͕   �_Φ   �C�   ��}    �o     W�9     ��?                                              ��      \�     ��      ��      ��      �;      �      �     ��     �� �  ��   ��� 0  ��o�0  ����0  �U�  ��[��  ���    ����    ��     ��    \~�    �_     �}0   ��C�   �o͕   W�y�  ��?}<                                            �?      ��     �e>     ��?     ��7      �      �     ��      �� �  ���  ���50  ��[�0  ���0  �kU�  �����  ���    ���    ��}    ��C�   �Ε   \~ͦ   �_N�  �}    ��     �o� 0  W�9�   ��?                                          < ��   � p�   � \�   ��� �{�� � �� p� � �;\= \���� �����  \Ϫ��>  p���  ����   ����    ��    <��      ��     ��     ��     ��     �     \~     �_     �     ��     �o     W�9     ��?                �      �      W      �   �?��    ��p9 <�e>\ ���?��  ������ ��   ��>�  � �?   ���   \Ϊ�   ܽ��   \���   p��    p���    �:��    ��     ��     ��     ��     �     \~     �_     �     ��     �o     W�9     ��?                     �      0     �3     <00 �   ��     ���0  ��     �� �    ���    ��s5    �_9    ��[    ���     �?     ��     ��     ��     ��     ��     ��     ��     p�     �u     py     \~     ��    ���    ���     �_     ��         �    �    �    0��           ��    � �   ��W   p�ϕ   ���    p��    ���     ��     ��>     ��?     ��     ��>     ܺ?     |�?     ���     ���     ���    ��     �_     �p     \�     ��     �\     �\9    �ys:    ���     �                                                             �      �e     p�     p�     ��     ��     �� <    ���    ����    ���0   ����   ���    ��    ���     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?                                                          �   �    � �  �e: �  ��> �  ��? �  � ��  ��0�  �� �   ��?��   ���_�   ���V?   ����    ���    ��?     ��     ��?     ��>     �?     ���     W��     \s5     ��     ��?     �s�     ���                                                               �      �e     p�     �    ���   ���  p���� \��  00 ܫ��� �� � ���> � �����?0 ����_� ����U  ��?��  ��?�?   ��>     ���     p��     p9�     l��     ��:     ��?     �s�     ���                                                             �?      p�      \�    �_�    0���   �� �   ��   ���    W��><  W��>   ���� 0  ����     ���    ��?     ��?     ���     ���     ��>     ۿ�     Ws�     \�5     p�9     ��?     W~�     ���                                                               �      \6      ��      W�      ��      �?      ��     ���    W��    W��   ����?   ��>   ���?   ����    ���     ��?     ��>     �    ���;    ��\9     �s     �s     ��    ��s9    ���?                                                                    ��      \�     p�     �     p�    ���    \�    \�?    p��    ����   �����  0���   ����  �s���   ����  ���   ��  ���    p��    p9�    ���    �_    p�W:    ���?                                                             �?      p�      \�     l�     l�     ��     ��    �<��   ���?   Ϫ�;  � ����   �p���   0p��?   ���     ��     ��?     ��>     ��     ��;     W~9     \s     �s     ��     �s9     ��?                                                              �      �e�?<   p� �  �s���   �����   ����   �� 3   �� �?   ��|   ���W  �����  ����>    ���    ��     ��    ���    ���     ��    ���:    ��s9     �\     �     ?�    ��\9    ���?                                                    ��      l�     �_     �v    �s�    \��?    \��   p��   p���5   î���    ����   ��?   0 ��    ��     ��    ���    p�    \��;    \|9    ps�    ����   �9 �   |9 p;   W �9   �  p5      \                                                           ��      l�     �_     �v     p�     ��    ��?    ��    0��    0�>    ��?    \�?    �_U�     ���    � ��    ��    0��     ���    �Vz     oy     ��5      �7     �_?     p�     ��                                   �            � ��    � l�   � �_    �v   0�s�   0���?   < ��  � ��  w���;  0w����  0�վ��   ��� �0?���    ��_    ���   ���    p��    p�    �9�    �5\     ?\9    ����    \� �   �� \      �     ��                                                         �0��    � l�   �0�_    0�v   � p�   ����    �?    0��    0��    0�>    ��>    �_�?     \U�     ��      ��     ��     ��     ���    ���     ��     <�7      �7     �_?     p�     ��                                                      �     �[9     ��     p�     �W     �Z    ��� <   ��� �   �����   [���   ۿ�W:  �����  �6��   ���   �����    ���    ��W    ��w    ��\    s5�    _9�     ��   ��[5   �5 �   ��       [                                                                �     �[9     ��     p�     �[     �k�    ��00    ���    ���    ���    ��?0    �~�    �U5     ��   ���    ��?0     ��     ��W    ���    p��     ��<     �?      ��     �V     ��                 ?      ��      0      0      0     ���    �[��    ��?   p�   �[�   �k�5   ���p5  ���p  ��   ����  ����    ܾ�0   p�     ��     ���     ���    ��{    ��_9    \>p9    Wp   ���   �� l   � l=   l ��   \  ?   p5                                                                �    �[90   ��    p�0   �[0   �k    ���    ��00    ���    ���    ���    �~50    �U�    ��?    ���     ��?      ��     ��W    �]�    pm�     \�     �?      ��     �V     ��                                     ��      \�     �    ��]    |�     ��    0�    �V9    |U:    ��}�    ����    W���    ���    �p�   W��   ��   ���    ���5     ���     �9�    �;\    \9�    �\      �                                    ��      \�     �     pw     p�     ��      ��      |��    W�>   �]��0   ����0   ��ٗ3   ��~�    ��    ���     ��?     ��     \~     �s9     ۳9     ��     ��     ��9     ��?                                     ��      \�     �    ��]    |�     ��    0�    �V9    |U:    ��}�    ����    W���    ���    �p�   W��   ��   ���    ���5     ���     �9�    �;\    \9�    �\      �                                    �?      W�      ��     �|�     �5    � |�    � ̧   � �U    e9    ��y:     �n�    ���    W>��    �p�   < ��   ��   ���    W��5    ����    ��9�   ��;\    \9�    �\      �                                    �?      W�      ��      |�     ��5     �    � ̧   � �U   � |e9    y:    ��n�     ���    ����    pp�   \��   \�   � ��     ��5    ����    ��9�  0W�;\   �_9�  ���\      �                                    �?      W�      ��     �|�     �5    � |�    � ̧   � �U    e9    ��y:     �n�    ���    W=��    �p�   < ��   ��   ���   0W��5   ����   ��9�   ��;\    \9�  <�\      �                                     �     �U:      �;      �= <    w �    ���   �?��  �_��0  p�{��  �W���    |z�6    �_�    ���     ��     ��     p�     ��      ��      p�      �]     �y     ��9     \]9     ��?             �       p      \      | �    \�   p~�   p͟   ��u?   ���0    ��50    l�9    \�9     l�     ��     ��     \;      \>      W:      �>     ��     ��      �      �      \      \      �      �      ?      ���     �      ��      �    �U�0     �{     �}     w�      ��     �w>     \W9     \�9     p}:     p�     ��     p�     \U     \�     ��     ��     \�     \^     p]     ��     ��      \�     ��   �?�    � �    ���    |      \��    p}�    ���    ��w     �]     ��      [�     \�     \u     ��     \�     \U     |�     ��      w�     ���     �9�     �5�      7�      �\     ��     ��     �5�    ��                <       �      �    ���    \��    ��?    �]s    p�|    ���     ��     �V9     pU:     �}�     ���    ����    \��    Wp�   ���   � �     ��     ��5     ���     �9�    �;\    \9�    �\      �                             �?      W�      ��      |�      �5    � p�    ��   |�w  ��ץ_   ���u  ���W�  ���   0 ��   0 ��   [�  � ��     ��      ��     ���     �5�    �5\    �7�    p9�    �?\      �                             �?      W�      ��      |�      �5      p�     ��   �s��   �swW5   ϳW:  0��p�    ��    < \�   �  \�     W�     ��     ��     �_     �p    ��p    �9\    p?�    p�    �\      �               �          ��0    �U30    ���0    |��    p]=     �W     w�     w>      ��      \z     \y     ��      �?      W�      W�      ��     �_     �\    �5p    �9p    p\    p�    ��      \      �                                              �    �[5    0��    �z    0[    �o    0o�     �Z�    p[�    ��y     ��     ��      �?      W�      ��      ��    ��_    �    W>�     ��     7 �    ; W     �                                              �?      l�      �?    � �     �[5    0po     \�     \�     W�     W�     �~    ��    ��~    �i�      ��      ��    ��_    ��     W>�     �7     7 �    ; W     �                                              �     �Z5     ��     �w     ��     �[     W�0    ����    ��    ��_9<   p����   p�7��   �����   ���    {y<    |�     ���     p��     p=�     p7     ��    � W      �  �      0      0      0�      ��?      �� �   ��Z5   0\��    p�w    �y�     _[     l�    ��v     ��     p�     ��     p�     \�:     \��     ���     pu?     ��     p�      p�      p�      ��      W      �                            �?      \�      �     ��    �s�     \��    \��    p�Uz   pzUy  ��^j�    �o�   �[�   � �>      ��     �U�     �w�    \��    �_    �\    �p:    p��    \ �   � �   <  W      �                                    �?      \�      �     ��     p�      ��    ��    �U:    �u:    �]    �    \�    �_�>     ��;     ��     ���     p��    p��    �[^     �_           ��     \�      ��                    �       �?    � \�    � ��   � ̭    s�    0���   0< ��   ����  wsu�  w]U  0�uZ�  0��[�9   0\}�  �  ���    �_�?    \��     \��     p��     p�    �W    �5|    \9�9    �?�5      \9      �                          �        �?    0 \�    0�   0��   � p�    ����    �    �U9    �u9    �]    �    �_�     \�>     ��;     ���     �]�     p��    py�    ��y     ��      �     ��     \�      ��                              �      [5     ��     �z      [     �o     �� <   �j~�   �k]��   ��Uu�   ���]>   l[�   k}5��   [� 0   �_�   0�n5    ��5    ۳    ��p    ���    �?\    ll5    \�    l5      �                                        �      4     ��     �z           �o�    ��00    lU�    l]�    �u�    ��?0    ���    �V5     �Z     ��     {u    ��_    �^m    �m�    �k�     ��      ��      [5      �         �            0    �0    [50   ��   �z�    [�?    �o�5   ��p5  ��Us  �nU�   �k��  �k��   ����    �6      ��      �U    �V�6    �_�5    ���6    �5�6    �p;    k�   �� �5   �6 ��   ��  <    �                                        �      [50   ��    �z0    [0   �o    ���   �U30    �]�    �u�    ���    ��50    �V�    �Z>     [�     k[    ��_    ��V    ���    ��?     ��      ��      [5      �      �7W��7                                                                            �      �e     p�     �    ���    p���    \���   ���   ����   ��   ����    ���    ���     ��     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?                                              ?      ��      0�    ��e�    pu�^   pu�_   \��_   ���9   ����;   ����   ���   ����    ���     ��?     ��     ��     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?     �      00      �      �     ���   \=�_   \�\   W�p9   ��e�5   �s��9   �s��9   ����   ����   ����   ����    ����     �>     ��?     ��     ��     ��     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?      �            �      �     �� <?   W��   W���   ����   ��e��   �p��5   �p��9   ����;   ����   ����   ����   ���     ��>     ��?     ��     ��     ��     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?                                                                      �      �e     p�     p�     ���    ��3    ��?    ��?    ���   ����   ���    ��    ���     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?                                                                                              �      �e     p�     ��     ��     ��?     ���    ����   ���   ����     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?                                                                                       0     0�    ��e     s��    ��     ��     ��?     ���    ����   ���   ����     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?                                                                               �     0      0         �      �e    �     ��?    ����    ����   ����   ����     ��?     ��?     ��>     �?     ��     ��;     W_9     \s     �s     ��     �s9     ��?    ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������           $ ( ,   $(,  $(,      
             " $ & ( * , . ������������������������@� �� @� �� ������@� � ���� ���� ��   �� ��� �� ��� �������� � 00�� ���� ��   ,�����,�����������,��� pp�� ���� ��   M�����M�����������M��� ��� ������ �   ��� m��� ��   �   �  � � �   ��09 �   � ������ ���? ��? ������ �   �� �   � �����   � ���: ��: ������ �   ��� �   ������   � ���: ��: ������ � � ��� �   �������� ���? ��? ������ � ��� �   ���� m��� m�   �   �l� � � �m�: �   ��������������   ��� ��� ����� ���� ��������������   ���� �0�� ���� ����� ���� �� ��� ����   �� � �p�� �� � ����� ��� @� �� ����   @� � ���� @� � ����                                                                                                �� �� @� �� @� �� @� ���� �� �� �� ���� ��� �� ��� �� ��� �� ���� �� 0� 0��������,��K��,��K��,������ �� p� p��믫���M�����M�����M������ �� �������묯� ���� ���� ��� � � �� ��L���� 묷� ���� m��� m��  � � �� �뜳��: 묳� �� ���� ������  � � �� �묳 � 묳� �� ����� ����� � � �� �묳 � 묳� ������ �4��� @�� � � �� �뭳��: 묳� ��m�� ���: � m � � l��� ���0�� ���� ����   �~���� G� � ���: ������ �� �����   ��� ���� � ����� ����� �� ��� �   �� ���  � ��� �� ���� �� �@� �   @��� �@�  � �� ��  @��� �                                                                                                � ����@�  � �� @�  �� ���@� ���@� @� � 0�����  � L�� ��  �� ����� ����� �� � p���,���� ���,����� ���,�����,��,�������M��p� ������0�� ���M�����M��M���m �� ����   ����:� �   �    ��l���� p: �<�� @��}���� �� ��  �� �������� � �O� � � ���� ��� ���  �8 ��������  � 듿 � ,�� ����������� p9 ����@� ��  �� � M��<����������� 0 ���@�� � 09  ��l � �  � m���  m�m l �l  m � ������� ������������ � ���� � ������0�� ������  � ������ � ������ � ����� p�� �����   � �� ��  � �� ��  � ���@� ��� ���@�   � @� @�  � @� @�                                                                                                 �����?�?�?<��??<? ?0�������??<?<?0?<?<?<?<?<? ? ?0?<�?<??? �<?<?<?<?<?<?<�?<?<?0?<?<?<? ?<? ? ? ?<� <�? �??<?<?<?<?<? �?<?<?0?<?<�? ?<��??�?� <�? ?3?<?<?<?0���?<?<?0��??<? ?<? ? ?<?<� <�? ?0?<?<�??? <�?<???3?<?<?<?0?<? ? ?<?<�?<???<?0?<?<? ?????<�?<��??<?<����?? �?<��?<�??0?<�? �<??�����<?<                                                ?<�?����?<�?�?�?��        ��UU  UU  UU  ?<???<�?<?<?<? ?  <?<?<    ���<?�UU  UU  UU  ?<�?<� < <?<�� ??<?<    ��� ?�UU  UU  UU  ��?<���?< <?< �?<    �??��UU  UU  UU  �� ?<�?  <�? <?<�?<�?        ��UU  UU  UU  �?<?<�? ?< <?<?<�?< <� �        UU  UU  UU  ��?���?� <������ �    ��UU  UU  UU                            �         UU  UU  UU    UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UUUU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU    UU                                          UU  UU                                          UU  UU                                          UU  UU                                          UU  UU                                          UU  UU                                          UUUU                                              UU                                              UU                                              UU                                              UU                                              UU                                                                                            UU                                              UU                                              UU                                              UU                                              UU                                              UU                                              UU                                              UUUU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU  UU                                                UU                                              UUUU                                              UU                                              UU                                              UU                                              UU                                              UU                                              UU                                              UU                                                                                            UU                                              UU                                              UU                                              UU                                              UU                                              UU         UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU       UU         UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU       UUUU                   @         P   P         UU                   @         P   P         UU                              P   P         UU      @                       P   @        UU      @                       P   @        UU      @                       P   @        UU      @                       P   @        UU      @                       P   @                @                       P   @      UU        @                       P   @      UU        @                       P   @      UU        @                       P   @      UU        @  @                    @  @      UU        @  @                    @  @      UU        P   @                    @         UU        P   @                    @         UUUU      P   @                    @           UU      P   @                    @           UU      P   @                    @           UU      P   @                    @           UU      P   @                    @           UU      P   @                    @           UU      P   @UUUUUUUUUUUUUUUUUUUUUU           UU      P   @UUUUUUUUUUUUUUUUUUUUUU                      @         @         @         UU           @         @         @         UU           @         @         @         UU           P          @                   UU           P          @                   UU           P          @                   UU           P          @                   UU           P          @                   UUUU         P          @                     UU         P          @                     UU         P          @                     UU         P          @             P        UU         P          @             P        UU         P          @             P        UU         P          @             P        UU         P          @             P                   P          @             P      UU           P          @             P      UU                     @             P      UU                     @             P      UU       <             @             P<     UU       ����������������������������������     UU       �                               @�     UU       �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��     UUUU     �������������������������������       UU     �1�0�0�0�0�p�0�0�0�4�0L�       UU     ����������������������������������       UU     �1�0�0�0�0�p�0�0�0�4�0L�       UU     ����������������������������������       UU     �1�0�0�0�0�p�0�0�0�4�0L�       UU     ����������������������������������       UU     �1�0�0�0�0�p�0�0�0�4�0L�              ����������������������������������     UU       |              @          P    =     UU       P              @          P         UU       P              @          P         UU       P              @          P         UU       P              @          P         UU       P              @          P         UU       P              @          P         UUUU     P              @          P           UU     P              @          P           UU     P              @          P           UU                   @          P           UU                   @          P           UU                   @          P           UU                   @          P           UU        @          @          @                    @          @          @        UU          @          @          @        UU          @          @          @        UU          @          @          @        UU          @          @          @        UU          @          @          @   P     UU          @          @          @   P     UU          @          @          @   P     UUUU        @          @          @   P       UU        @          @          @   P       UU        @          @          @   P       UU        @          @          @   P       UU        @          @          @   P       UU        @          @          @   P       UU        P           @              P       UU        PUUUUUUUUUUUUUUUUUUUUUUUU   P             @   PUUUUUUUUUUUUUUUUUUUUUUUU   @    UU      @   P                           @    UU      @   P                           @    UU      @   P                           @    UU      @   P                           @    UU      @   P                           @    UU      @   P                           @    UU      @   P                           @    UUUU    @   P                           @      UU    @   P                           @      UU    @   P                           @      UU    P    P                                  UU    P                                      UU    P                                      UU    P                                      UU    P                                            P                                    UU      P                                    UU      P                                    UU      P                                    UU      P                                    UU                                          UU                                          UU                     @                   UUUU                   @                     UU    TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU      UU    TUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU      UU                                              UU                                              UU                                              UU                                              UU                                                                                            UU                                              UU                                              UU                                              UU                                              UU                                              UU                                              UU                                              UUUU                                              UU                                                �    W9   ���   �~�    ��    [9    l   ��   �]�  py�  l��  ��>  ܗ�;  \[�9  ��9  ���5  �W�5  ח�9  ���:  <�??  ��5�  חו����}����u 7�9� ����  |�  ���   �   �V9   ���    w�    ��    W9    \   ��>   ��  ���  ��  ��  ܫ�  \�~9  ���5  ���5  ׫�5  ��6  ���6  <�?  ���5  ��u�  �5w��9�w��=��������  s�  ���      �  |5 ���  ��  ��  \:  �  �9  p9  \��������~��������|����|w�����W����� ;� 7p 7p ;� ��  ��  ��  �0  0     �  \=  k� �7  ��  �5  �  l  l ��5 p��?pk[�pk�7p����o�Z���o=���װZ�=���ְj�?��� p7� �7� �� �; �7  77  7;  ;  �� @(�P@X��@���@���@�A�@AH�pAx��A���Aؒ B�0B8�`Bh��B���Bȓ�B�� C(�PCX��C���C���C��i� ����� `��8�� ��� `��i� ������;��� ��_���� � @���#8�

����������������������/� ������� `��8�� ����Bd��
&
&
&
&���
&e��e��i ���i@���i����i����/� ������� ` �é����腼�D��� ����� ������� � �� p� L������� `��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������              �?                |�               ��              pP�              U�              <L�              �L��             �^_9             �7��           �\w��          �W�0ޑ_�         | �s]���         �F�xU�         G��u�A�         L�py�T�        �\�x��>       �W�0��s�       | �s9 �]�?        �F�8 �7        <G��� �w       ��M�py� \�       |�]�x��       ��7���       |P�w9 �] �?      U��8 �w |�     <G�_�� ����   ��L��z� \�pP�   |�^y�� �J  ��3��_�� L�  |P�s��] �?L�09  U��T_�w |�p8  GU�������79��  LJ9 ���|P�w8��  �� GB� UF�� � �0� LT� G����  p�\�>�?L�0y��  ��p�|�0yGA�  ���>��790]T�    S�|P�w8]]�>    G9  �F��G���    L:  G��QP��?     �  L�0ySeP: �    �  pxG���       09��L� @       p4|�: �A       ���09 �>9       �QP:p G�w8        S�� S~��        G�  ��W��        L  _9�W}�        9 ����G:        09 T�U}�        p�A�WG�         �p�>�ב          0�L�� �9        09 \�� �       �8p8�Wy��A�       9��|�x��>       ����G��MA�        � ����>         � W� �s�         � � ��>          0 � ��              �              �A�               �>              �A�               �>                �                <      ����������������  OO���O��3��T3�<�  �t=5]�5]s]����L�  �}��U_��s������? �u��_���s]���5��4 __���_}Us��U�u]�5 ����������������?                          �?                      0       �?      �          �?  �  �  �      �     �A� �?  �  \�  [: �9  C4      D �  �� l� �A4  ׯ��� ��� � �      3w 4  ��  �����  �}���  w� ���      �����  L�  �� w�  ��w�  �� �w�     �M��|�  �  �� ��  � ��  G�  ��  �� �� ��  �  O��G�  w��G��]��G��A��ty��G�������\�����\��?�p\������[z���]�t�~�?��p�e�_��t���_�9��������0CC4��t�~�QZ��ח9��A�t{�ꩪtT���f�0D� ��]D�T�U�����������������w���?Q���C3w�TDW��w�}ߥUwߩ�ww��|ߩ���U�?��w�EW���U3wW�w�OU��U��j��y����GyU�?�v��^N�]���WUӔWUG�f�G�j�G���G���_�V����5GyG��u�O�V�G����k�\�k�]����{�_�[�A��5]^�q����[�]�o����?���w��z�}p�^y����_{_}��}t�n�?w��g�ytë{�Ѯ�f�_�P�?���t���ҝ4��t]���v������@T�����?�ѩ�A�ה�TS>�ҭ[:ў��W�������Q�9�o����O����ۥǟ��z}dӦ�U�N�[�ww�w� ���U�Ou��}���ݚ��}���OY���U��^��yT�� �}߹ֺNy�N뫪N�j�����NZ�w�U�z��G�UG�AT������y�嫪�j���������U��~�]�G�]��G���A�{�sy��q���q�{�A���G�W��]�_��_�������������nz��Ѥ��\�^DSDs���u�[��䩪���MDC��9��D��C�_�^]�3w��y���e�A�����@S3wQ����3w����s�^�m����������������@S��P�UV�ݫ�޽�P{w��N�٩w��w�UU�ݪ�w�P�M�[T�OUYN窪N�ו����妦��v���VUN窪��D��]T�NUY媪喧�������G�z�G�W�媪G�U�tym���՚����Z�������]���^�[�q���]������A�w��������A�Dӝ��?���_�_u��_���]o餪�ҭ�ѝ[z��3w�S��w�yp�o��]Dw�A�WS����DW�DGצ�M��WG�������@o9S3w����W����3wW�3wW����M�����}���UW����ݖ[�ݫ���W���W�w����m:M痛��DC�OU�M�A�O�^N竪N�V�M�[�����ty�:�V�G�QS�NU����奞媪�U�坮Gy��������UG��f�ty���������V�ty��_���ҭ���k����A����M�ݫ�ݫ��[���_��ud���֭��e��u��n�ҭ��]���]��ҭ��ҭ�zp׮9���~e��{�V�5��n}d�~9 C�> C�zd��wd���P�����������������������������������������UUU9mUUUUUU9mUUUUU�q|^UUUUU9mUUUUUU9mUUU���~�������~��������8������~�������~����������������������������������������~�������~������?�������~�������~�������{�������;߷������׿����~�������{�������~��������p�����>y�����?��������~�������{��������Q�������������{�������{������z������zG�����SUU������z������z����z��������_��������������{�������z�������z�����窪����绪���y}����z����z�������ݔ����z������{Ծ������z�������z�����U����:�����������z����z�������4Q����:�G������������z�������z�����������������<@��������z�������������u����NC���4D�������������������������O=������_���?��O���������UUUUUUUWUU���w}UUUu��{UU5=MW��UUWUUUUUUUTU  ��@5}UUUq_�;U5=MCU �WUUDDEDDD�����u^UUEt_�{DEu= M�����UTDDDDT1U��s�^UU�]��TQ5�L��j�yUDD @D �������_U���UT�3������?D D  @ wU��t�yU �U�T4MNWUpGA   @@   �|���t�  �C� 0N^G]U �      @      �] p��4�  w�?�Cp�y �              ��9y�   �5�S �3}�~                  ��t��   w1� �s��          @          ���y?   wL� ��~�                      9�    ��@ 0C9                       ��?     � P ��                               � T                                    �                                     3@                                    �P                                   ��T                                   ��U                                   ��OU                                   03_                 ������������������?���������������������������������������?���������������������                  p3OU                                    ��E                                    ��SD                                    ��S                                    ��G                                    3�T                                    3�U                                    7�T                                   ��<E                                   ��<U                                   03U                  ���������������������������������������                 ��OQ                                   3�OQ                                   7�WU                                  ���CQ                  ����������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@ P TP PP UUT@@PPP PUUUU
� B��ZB BB)TU���jB B BUUUUP ��T� 
�U�ZP�� �T� � 
�UUUUj ���Pj �UY��Vi�� �ZB � �UUUU@ � hV �U` TUh�(P�
� �UUUU���i����Z�ViZjUUj�ZU�Z��Z��j�j���i�jUU�����������U���������U�����U�����U�����U�����������T���������T�����T�����T�����T������T��γ�Ļ�T���T���T���T����������Ϩ��������飯���Ϩ����Ϩ����Ϩ�����������T���������T�����T�����T�����T��޷޷޷޷�T��޷���T��޷�T��޷�T��޷�T�����������T���������T�����T�����T�����T����������� ��������� ����� ����� ����� ������T���ĳ��T���T���T���T�����������T���������T�����T�����T�����TU          TU        TU    TU    TU    TU����]����WUU�]�����_UU����UU����UU�}��UU����]uu�uUUU�]��]��UUU]]u]UU]��]UU��u]UU����]����WUU�]��}}�_UU�}u�UU]��}UU��u�UU����]Uw�UWUU]]�u]�U]UU�]u�UU���]UU]�u�UU���_W����WUU]��u���_UU��u�UU����UU]�u�U�����������U���������U�����U�����U�����U�����������T���������T�����T�����T�����T������T�ĳ�Ļ�T���T���T���T����������Ϩ��������飯���Ϩ����Ϩ����Ϩ�����������T���������T�����T�����T�����T��޷޷޷޷�T�з�Կ�T��޷�T��޷�T��޷�T�����������T���������T�����T�����T�����T����������� ��������� ����� ����� ����� ������T��ĳ��T���T���T���T�����������T���������T�����T�����T�����TU          TU        TU    TU    TU    T������������������������������������������������������������Ļ��ĳ���������������������������������������������Ϸ޿�����Я�������������������������������������������Ļ��Ļ��Ļ����������ĳ������������Ϸ�Է������������������������������w��ej�dftw�̫��"Fyt 8��Bk��R6��S4W��Eh��f��ʇ���eUVxvfx��y������wwwfgwwwxwwx�www�wx�����������������wwww�wwwwwwwwwww�x�������������������������������wwwwwww���w���wvwvwy�����wwx�w���������vfx��vx������wgwwwwgx��wx��������x���wwx�wwwxw�����wxx�������������wwwwx���������x���wx�������x��wwx��wx���x��wwwwwx�������x��vw��wgx��ww���fx��wx������wx���wx��www����������wx���x���w���ww���w���w����w���������������x���www��wx���ww����������������������������wx����w����ww���wx���x���w���wx����w���wx�������wx��w����wx��ww����w����x�����������w����x��������������ww������������x����w���������wwx���x������w���w���wx��ww������ww���������x���x���x�������w�������������������wx�������ww��x����x��w�������ww������������������x����w����������������w���wx�������wx���x���w���wx�����������������������������x���w���wwx�������x���wx���������������������������                �w��ej�dftw�̫��"Fyt 8��Bk��R6��S4W��Eh��f��ʇ���eUVxvfx��y������wwwfgwwwxwwx�www�wx�����������������wwww�wwwwwwwwwww�x�������������������������������wwwwwww���w���wvwvwy�����wwx�w���������vfx��vx������wgwwwwgx��wx��������x���wwx�wwwxw�����wxx�������������wwwwx���������x���wx�������x��wwx��wx���x��wwwwwx�������x��vw��wgx��ww���fx��wx������wx���wx��www����������wx���x���w���ww���w���w����w���������������x���www��wx���ww����������������������������wx����w����ww���wx���x���w���wx����w���wx�������wx��w����wx��ww����w����x�����������w����x��������������ww������������x����w���������wwx���x������w���w���wx��ww������ww���������x���x���x�������w�������������������wx�������ww��x����x��w�������ww������������������x����w����������������w���wx�������wx���x���w���wx�����������������������������x���w���wwx�������x���wx���������������������������                �w��Uy���1 $h�����ʆS   5i�����S!#Ex���˻���fffwx���������wfwww��x�������ww��wx�������w�������wwwwx���������������x�x��������w��w����������x������������w�������ww������������x�����������ww�������������wwww��������x����������x��������������������wwwx���������������������������������������������������������                ��������i����!� 	� \ 'q 2!"4VDEh��h�ۻ��������������������������쇾�Ez�Fu  Q                            #42#VeVf��w����˽���������������˪��ۘ�������������������������������������������������������������̻��������˻�̻�����������ffvUDC332                          "#324D3DUUUVfgffwwgxwwwx�ww�ww��wwwwwwwwvgwfgvffffgvgwwwwwwx����������������������������˻�������������wwffeUUTDD3333""""""""""""#333DDDDUUVffwwwx���������������������������������������������������������������˻�������������������wwwwwvfffffffUUUUUUUUUUUUUUTEUUTDDDDDDDDDDDDDDDDDEUUUUUUUUUUUUUUUUUUUUUUUUUeVfffffffffffffffffffgwwwwwwwwwwwwwx��������������������������������������������������������������������������������������������������������wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww��                �����������������������������������������������������������������������������������������������������������g�@�KV�������o���  �   `    ���(���������������@�0���P���������             �PJm�~���������������������ٶ�
p\_��I�P                       ?o�������������������o�u� b        # @(� @          8��������������������������W�B�a       ��<P�R����)"�?��Tf����������������������&�@              $ %Sl������̞��)�50F��X��������������������o�d��Q                @�n��������������������{猃z��4sWRfGA aEf����W�h���v�6Tc�8TFr$&eVTVGC�k���������������������eW2 0            E8GU>���������������z��G��X6=U4q6G�S�xF������G��5K�1b Q3B#5F�$�3xuh�W�EGu�������ܬ��������������ʗ�cU       4!��e�����x���ݚ���������}ּ��ic{e~�3f�uId�X�x�y{v~ۅz�gxw�y����W���ggGde#Ev%dGSTFggtifkhf����������������ۻ���8CfT3$1tTSTGBx%TJe�eewsw�V�xdytxY��������������������tFC3   10SWf����̻�쬺�ʌ����ewFg4r$"%2V2eGdh��z����̽�������ܺ����wVvT%TDER2D32UcU6cxww��y��������w�j��g�w��v������̬����������˪�v�44#       !DdXx�������������껩�v�WwfvdvFvVwgwy��y�j���xvvFwDfWuwV�v�x������̫�˻����G�WeT5DVDFefV�v�����۫�ܼ�ܺ�����xwvfVfwgewffwhvw�f�wx������g�wvh�x���������v�wehdVVeF�Wxv�y��˹���������ۛ��efD3       35Txx��������������ʺ���eeEcED5ETFvfvy����������xx�fuWUeUFfWfWww�y������ܽ��̺������gugeUFeFTTFffxw�x�����˼˻�����wuUUDD3B"""4CUUvx��������������̺���xeUUDB4"31#3DDTVUWvVwvgx��������������˻������x�wudUTDTDDUEfwhh�x���������������xxwgwgfgWgww���������������������������x�x��wfwfUVTTETEDUVffy���������̻�̻�����wvuVdUDDUUCUVVgx��������������y�wvwufefVeffgww�������������������wwfvgfffVfvfVfvww�wx���������������wvwwgwvwwwwxw�w�����������whvfEVUVeeVfwww���������˼������ufUTCDC3DDDDVff����������̻��������wffTeVEEUUUffw�����������������wwvffVeUeUUVUWgxx�����������������wvfeEDUDDDTUEUfvwx������̼�̼�����wfeTD332"#333DEffx�������������̻�����fUTD4333C4DEUVfgw�����������������wwwwvfffffgwww����������������wwwfffUUUUUUVVfffwx�����������������������wwfffffffffffffgwwwx���������������������                �� ���  ��� � ��� � ��� ��" ���! ��d-��/��.� �&���'�'�%�&�$ ���'�r� ��'��d�(���)�'�'�%�&�$d-��. ���)�)�)�%�(�$��.��- ���)�D� �Lܮ � 鯥'�%��.�&�$� �- ۯ�&i�&�$ ���(�$��- ۯ�(8��(�$ ���(�T� �L ���/��.��-�L�$�J�% �� �� � ���2 鯈� ��� `H�Z�-
����� �����.�*�/�+�%�,�%� Յ0��Յ1�$JJ�� %!�0� ���+�Ȁ��*�
�,�/�+�L��z�h`H� �! �����!h`H�Z�/���� ���� ��z�h`� �3�4 �� ��� � � � � � � � d^d_`�3���D�4���(�?� ���8�9� �  ���L� ���E�F� �  ��?�?�:� ���L�L�G� O��4���(�Y� �� ���R�S� � � �  8��Y�Y�T� ��`�5�6�8ȱ6�9ȱ6�:ȱ6�;ȱ6�<)
���=��>Ȅ5d?d@�:� �"�A�鲅6�鲅7� �
�6� �dA���Ad5��`�O�P�RȱP�SȱP�TȱP�UȱP�V)
���W��XȄOdYdZ�T� �� �4 �� ���8�9� � �E�F� � `�B�C�EȱC�FȱC�GȱC�HȱC�I)
���J��KȄBdLdM�G� �"�N�벅C�벅D� �
�C� �dN���NdB��`H�Z�;)?	@�\�;*��%\�\�@�=��<)@��J��\�\Ȅ@�=����@�<d@�\�^�� �^z�h`H�Z�H)?	@�\�H*��%\�\�M�J��I)@��J��\�\ȄM�J����M�IdM�\�_�� �_z�h`H�Z�U)?	@�\�U*��%\�\�Z�W��V)@��J��\�\ȄZ�W����Z�VdZ�\� � �^�_z�h`� d^`� d_`��P�QdO��[ �� 8����4` �� /2�   �

		�
	�    ��  ����޲���� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                    ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������dxآ � �� �� �é�X� � �dxآ � �� �� �� =���X ��4 ���q �� �� �L�H�Z�' J� k��$ �	J��%  q�z�h@���# `�`H�Z��f� � ���\�����d��  I�����,) ��)��)��*��)���+����� H�H�H�H�H �h�h�h�h�h� � #�z�h@� ��  (�`�EH� b¥ w¢dd &&&8������������ ���h b¦� `�EH� b¥ w¢d�d��&� &��e����e�����榁��h ���`��I��ݥ�I���8���ޥ���`� � ����`� ��`
� ��e � �i ��� �� �� �` ��l  � Z� �� � ���� ��0	��z��L��`Z� ��������������0	��z��L��`	 I�i`H� �h`H�I���I�����h`�e � �`�`�e��`�`�e����`�`e����`�`e����`�`H� I�� �I��� ��h`H�I���I�����h`ڢ �JJJM
j.
....����` ���
�L�H �8�����8��������h �`� I�� �I��� ��`�� H�H��H��H�� d �ũ  h�h��h��h�h� ``���H��)��h




����& `H�Z� ��  	 � �� � ȱ � ȱ � ��� z�h`d�����`x ;é�X` �Ü � � � `� � � � `H�Z� H�H�@�� � � �  ��h�h� z�h`���ڊJJy Յ����i ���)�����ʅ������%������`�{�G�a��a`�[�<�A��A`�:��0��`�.��$`�,��%`�'��&`�"��'`�?��(`�!��)`�`��H�֠� ����h�	i


������,�� ��� ��Z ��z��m����L[�H�m�h�`lH �é �h �â��  ���i����i�����
i̅��	����	� ���� � ����� �����������i0���扥�i0����Ɔ��`H �é �h �â��H ���i����i�����
i̅��H��	����	� ���� � ����� �����������i0���扥�i0����Ɔ��h��`�� �������ȱ�����i/��������`��)H����H��������h`� ����Z �â�
� ������i0�������z������HZ�.*.*.*.*)������ ��hzi�h��Ɔ��`��)�����)���`���
I|�I5�	�I�` �å���`��H��H�e�iJJ�
�
ڦ����I��he�)����I��	��� ��%��� �
�ȑ�����%	����i0�������h��h��`�Z��H��H�	�e�iJJ��ʆ
����t��� ����ȥ���ȥ
��ȥ	��� W¦	�
��������i0���扥 W����h��h��z�`�t���u���v�
��w�	����x���	�
��������i0���扥 A����`��H��H������I��	���%	�����i0�������h��h��`��e�JJ�	�����I�2��������=������ ������	�����	���e�)����I�1���ڦ�����=�����`����������� cǭ�m�8���� �î�� cǮ��� �ì� 3Ǭ���m�8�� �ì�L3ǩ `��`�چ�
����-�I�����A��i��� � ���0����-�&�������0���,�����)�ɠ ���Ѐm)����
I

��@�  �ɀTH��	��h}���I

�ڹ˝ �O˝ ��i� ��ڦ�)� �Ȋ������	@�� ��	@� ��0L�`H� � ��� �  ��he � ��)�Ff Ff Ff ��)���� `0�0�1���A�lɉɳ��ɣ�`��
i� ��L������I�-��� � ���� }��� ���( `�)������ zÜ �( �`��i�ڦ�)� �Ȋ�����`���������`��i� H ��� � ���  �����h`hL;í8�


e瘝�Yޙ� �Zޙ� ��`���� zÜ �( �* ��Ll�


�� �Qޙ� ���������t�������������`1 Player 2 Player Beginner Intermediate Pro Select Level Fault Out C  Game P  Game C  Set P  Set C  Match P  Match 0123456789ABCDEF �  �  �  �     ����     U��0�����?� @��v
�F�F��o/�R"�ʢ|X7�����zdP=+����Ǽ������}voic]XSNJFB>:741.+)&$"                                       �������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������                                                                  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������                																















 @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @��    				



    !!!!""""####$$$$%%%%&&&&''''(((())))****++++,,,,----....////0000111122223333444455556666777788889999::::;;;;<<<<====>>>>???? 0333<???<???<???0333<???<???<???0333<???<???<???������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^_____`````aaaaaabbbbbccccc�ď�4��T�� �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �  ��  ��  ��  ��  `�  @�   �   �  �  ��  ��  ��  `�  @�   �   �  �  ��  ��  ��  `�  @�   �   �  �   �HF �H j��d P����� x� ް   ޱ   ޲   ޳   ޴   ޵   ޶   ޷   �������   
����   ��   ��2��������   ��(���   ������   �����   �� �&�   ��������   ��������   ,�28�>�D�J�   2�   P�(V��   \�b�h�   ��������   ��������   h�n�t�z�   ��������     �ք�  y
         �֊�  �
         �x.�?�?�/�    �<?�?�?�?�  �
�*�
��?�5b�5���1_��o��	$   �$   �$   ���                        �                        �                        ��  �0   �0   �	  ��  �0   �0   �	  ��΂< 0 0< _ < 0 0< _ H 0 0< _ F 0 0H _ : 0 0: _ : 0 0: _ : 0 09 _ : 0 0; _ < 0 0< _ < 0 0< _ H 0 0< _ F 0 0H _ ? 0 0? _ ? 0 0? _ A 0 0F _ E 0 0A ^ �� lن �� pن `� lن `� lن �� pن �� lن �� pن `� lن `� lن `� lن `� pن �� lن �� pن `� lن `� lن �� pن �� lن �� pن `� lن `� lن `� lن `� pن `� pن `����H U H D F K H > "K G �F � F O E D F 2 .K O J M H K J O H U H T F Q H G K K �M � M \ K 9 �H S H D F @ �H ^ H N F V 
H R K E �F � 0F M E N F / 1K N J N H J J Q H O H M F U H I K P �M � 	M P K < �H F H _ F G yT � R X Q S O [ �M � M [ O V 
Q ^ R Z Q U O _ H B T � R U Q O O a �W � W R V [ eT \ T \ R W iT � R Y Q Y O [ �M � M \ O ] Q Z R Z Q ^ O ] H P T � "R ] Q [ O \ �W � W T V N rT \ T F R Z f��΂7 ^ 2C ; U7 - 39 - 9 - 3E > R9 ( 8; - ; - 3? ( hB ) 7G + 5; ( ; ) ; , ���; - > 4 ,; ? Q7 7 )= * @ 9 '= < T9 1 /? ) B ; %? B ;  ? " B & 
G 6 �� lن �� pن �� lن `� lن �� pن �� lن `� lن �� pن �� lن `� lن `� pن 0� pن 0� pن 0��ي�    (��    t�t�    Eڌ���  ]ݭ���          ���������	�������� ������� ����ɪ�e�ɿ����`���� ��iJJ���iJJe����	� ����ȥ���ȥ��8��
ȥ	��Șe����橦	�
��������i0���扥�e������ޥ�� �������L1��� �� 0`�� ��ȱ ��� ��ȅ���ȅ���ȅ8��
��Ȫ� A¤
��������i0���扥�e�������`�����Hȱ����h�������`���)�-��)@���	@��� ���L�ߠ��8�������芑� ��`���� ȱ����
e�� �ȱ �ȱ �������) ���	��`� ��� L�ߠ������`Z�� �� ��z �å�
i̅i��Ԡ �� ����0 å�iJJ�	�08�	�
������ɪ�Xe�ɿ�Q���L�	� ��I�������� ��� I���ȱ�I�I���֑���i0���扥�e	����Ɔд`ZH����� ��hz`ZH����� ��hz`����������)�����`��� �w
�� � � �� �� �� ��u
���� �ƀ� U� �� �� � � ���0& K���w
����
)� � ��L� |�Lး�����w
�٠h�  ;�d�dŜ�d�dϭw
��Y�t
�% ���; ��ʠ� �� � ���x
�x
�� |�L� ��� ��ʠ� �� � �� |�L�8�0� E�� |�L�w
��	 �� �L�̅ �ͅ�ȅ�Ʌ ����8� �̥���ͥЅ �х�ʅ�˅ ����8� �Х���Ѧͤ� ̈́�L-���d�d�d�d�d�d�d�d�d�d�d�dխ��	���ǩ���`dǩ��`���dũ�ĩ��ǩ��ƥ�¥��d�d�dͩȅ�d�d�d�d�d�d�d�d�d˩��dɩ��`���dũ��dǩK�ƥ�¥��d�d�dͩȅ�d�d�d�d�d�d�d�d�d˩��dɩ��`��t
���w
�٠`�  ;é؍V�a�U�_)�	 �_���d�d�dͩ��d�d�dѩ���d�d�d�d�d˩��dɩ��`��t
���w
�٠`�  ;é؍g�ʍf�p)�	 �p���d�d�dͩ��d�dө��ѩ��d�d�d�d�d˩��dɩ��`��t
���w
�٠d�  ;æ�� � Ff �iF��i ��e �Њe�ѥ iP�̥i ��d�d�d�d�d�d�d�d�d˩��dɩ��`��t
���w
�٠d�  ;æ��� Ff �iK��i ��e ��e� фХ iv�̥i ��d�d�d�d�d�d�d�d�d˩��dɩ��`�ä� 8�/��� ��Ѕ �х 8��� �Ǥ� 8�K��� � ���Մ�`�/8�� �Å�Ѕ �х 8��� �Ǥ� 8�K��� � ���Մ�`�/8�� �Å�Ѕ �х 8��� �K8�ƅ� �ǅ ���Մ�`��Å� �¥8�/��� ��Ѕ �х 8��� �K8�ƅ� �ǅ ���Մ�`�t
dѩn��dͩ҅�d�d�d�d�d�d�d�d�d˩ ��dɩ��`�t
���ѩ���dͩ҅�d�d�d�d�d�d�d�d�d˩ ��dɩ��`�t
���ѩ��Щ�ͩ"��d�d�d�d�d�d�d�d�d˩��dɩ
��`�t
dѩ���dͩ���d�d�d�d�d�d�d�d�d˩��dɩ
��`�ƅ �ǅ�ä� {�� d�S� 8��i@��i��ƅ �ǅ�Ť� ��� d�>� 8��p8倍�偍�����ƅ �ǅ� �  ��� d�>� 8��p8倍�偍�� ���S�� � ������ ���>�� � ������ ���S�� � ������ ���>�� � ���i��i ��H�J�7�9�I�K�8�:��H��I��7��8�����������	��
���`�Z�� 8��� ��� � ��h8� �h��`�Z�H� Hd�d� 8��� ����� ��h8� � h��he �he�`���� �� {�� d�S� 8��i@�p�i�q� � �� �� ��� d�>� 8��p8倅r�偅s�p� �q��S�� � ���8��p�� �q�r� �s��>�� � ���8��r�� �s���� �� {�� d�S� 8��i@�t�i�u� � �� �� ��� d�>� 8��p8倅v�偅w�t� �u��S�� � ���8��t�� �u�tɯ�dtdu�v� �w��>�� � ���8� �v�� �w``O->��H��O �ߢ�` �ߢ�- 6ߢ�> 6ߢ�` i�� 6ߢ�O i�� 6ߢ�O i�� �ޢ�` i�� �ޢ�> �ޢ�- ��h���� hå���`�����)��/������%�������
�������������� `����`�p�j�l�r�k�m�t�Y�[�v�Z�\`��i��̥�i�����eԅ֥�eՅ���e̅Υ�eͅ���eЅҥ�eхӥ΅ �υ�7�� � ���eąĊeŅť҅ �Ӆ�-�� � ���eƅƊeǅǥօ �ׅ�-�� � ���eeÅæפ�d�-� �֦ׄϤ�d�7� �τΦӤ�d�-� �ӄ�`�Ʈ��I�i�:��® �I�i�7�i0�`� `�ƅܥǅ�dߩK�� z��M�ƅܥǅݩ��ߩ��� z��8��i� ��i �� �ܥ��dߩ/�� z��� �ܥ�ݩ��ߩх� z���`� `����%�Ǥ� �� ����ąܥŅ�dߩ�� z�� T�`��i�����-i���%��i������ƅܥǅ�dߩZ�� z��� `��`�؍g���f�p)��p�؍V�@�U�_)��_L��5�6���L@�"� �2 �id� � �d�K��d�����驵�����م�d�K����������驵��d�)��dǩK�Ʃ؍g���f�p)��p�2�؍V�@�U�_)��_�n� ����驵��d���d�K����������驵��������d�K��d�����ǩ��Ʃ؍V�F�U�_)��_�؍g���f�p)��p�2 �� ����dũ�Ģ����Ä�dǩK��d�d�d�d�d�d�`���L����8�¨��ê ݄�dߩ�� z���2�.�0�؍g���f�p)��p`��ܥ�ݥޥÅ� z��� �}��� �(�+�*�������0���؎+�*��0I�w
�D��ܥ�ݥƅޥǅ� z��
�-�n�,�%��ܥ��dߩ
�� z�����-���,�d�
���$m*�$�%m+�%�&m,�&�'m-�'�&� �'��(��)� ���e��e��$� �%��(��)� ���e��e��%�$�(��)� �%�$�'�&�(��)� �'�&��ܥ��dߩA�� z��d�@���ܥ�ݩ��ߩ��� z�����㩿���ܥ��dߩP�� z��d�O��+*�Q�+0i�0�.�A�.�0�2�5�؍g�֍f�p)��p��2`�2��؍g��f�p)��p��2`�2`�2`2#�$�%�&�'�qʽ��#���(�)�*�+�,�-`���W�2�^�,�-��� �� ���$���+�P�*��0�3���+���*���0�"�.�؍g���f�p)��p�2`�#��#`L���2`ü��u������j�l�k�m�Y�[�Z�\��� �� ��p�j�r�k�t�Y�v�Z`�����Ä����ǩ��ƭ��(� ��؍g���f�p)��p�2L��4� �Lu�`�4� ��!��؍V�X�U�_)��_�3L��)-*�!��)0��)�*�؍V�X�U�_)��_L��L����E�4� � u��ąܥŅ�dߩ*�� z��' b�2� � �ix�� �I�i�ԩ���`��d�`�4� �;�ąܥŅ�dߩ*�� z��' 
�3� � �ix�� �I�i�ԩ���`��d�`�ąܥŅ�dߩ�� z��.������é��©؍V�F�U�_)��_��- 6ߢ�> 6�`�ąܥŅ�dߩ*�� z��^�)-*�V��)0�P�)�* 
�  � � (� �� �ť�




���0�eԅԊeՅե�I�i



���0�eЅЊeх�`��Æ� ,���L��Lu� �­
)i���������ąܥŅ�dߩ*�� z��ӥ�8�¨���ê �� �������8�ƨ���Ǫ� Ю�����ܥ�ݥޥÅ� z���؍g��f�p)�	 �p��ٍg��f�p)�	 �p��2�.�*�+�,�-  ��ܥ�ݩ��ߩ��� z����ܥ��dߩ%�� z��
�
)� ���ܥ�ݩ��ߩ�� z�� �� ���� 9���� ��Lu��5�F��)0�7�L���5��8�¥����؍V���U�_)�	 �_��؍V���U�_)�	 �_��8�¨���ê �� б����ƅܥǅݥ�ޥ�� z�����8�訥����1�
�-��)�ąܥŅ�dߩ*�� z��������� ��  � �� �� u�`��ܥ�ݩ��ߩ�� z��� `��ܥ��dߩ�� z���`�`��ܥ�ݩ��ߩ�� z��� `��ܥ��dߩ�� z���`�` �ť�����0�e��e���� �0��ܥ��dߩ�� z��� ���ܥ��dߩ*�� z��� �)�2��ܥ�ݩ��ߩم� z�����٥�ܥ�ݩ��ߩ��� z���������`�_)0� �`�0��؍V�@�U�_)��_�5�:�;` �Ŏ8�9�8�խ9
I�i���0�e��e���ܥ�ݩ��ߩ��� z����������ܥ�ݩ��ߩ��� z�����驡�襶
���0�e��e���ܥ�ݩ��ߩ��� z�����穷���ܥ��dߩK�� z��d�J��8��9�;�>�9�;��8�:�.�:�8�؍V�m�U�_)��_��؍V�|�U�_)��_`����)�t
� ��ʠ� �� � ���x
�x
�� |�hhhhL�` ��Ѥ� �� �,��(�դ� �� ����ąܥŅ�dߩ�� z�����`��i������i�����i������i����`�����(����L��I�i��L��4� ��8�� ���1L�� �­
)�����L(�I�i��L��
)���5L���7) �U����0����0�eЅЊeхѦ��
 (� ���I�iJ��28����I�i���0�eԅԊeՅ�`���
 (� �䥷��L��Lf� �� �Ü � �ׅ�ȅ �$� 1�ׅ�΅ �.�� 1�I���ʅ��0�l�  4ĩ  �d���l�"� ����������)����)@��ߥ�)������Ӧ��� ��ƩH� ��h` @�@�A�G@H U�U�V�\@]� �  � � � �  � � ��U����U�� �Ü � �	ڽ��H�
����� �����������h ����ߩ[���ʅ��(�@�  4ĩd���ʅ��(�P�  4ĩq���ʅ��(�`�  4ĩu���ʅ�� ���  4ĩׅ��� � �
 1�ׅ�څ �h�
 1�  �d���@�� ����������)��8��)@��i��� �� �ɀͥ�)������e������Ņ� �ɀ���H� ��h`���<� ڦ�� �â���hH�<����Ά��� kť�i�������` ��G�;�ؠ"���ؠ1�V�U�_)�	 �_�؍g���f�p)��p� � � ������ �Ü � �ׅ�ԅ � �< 1�  � t� %� ����������)��������)����+�G�L�`�4�0 �é����"�����������0 L �������0 L© A����`�|� �í% ���|�0 �í& ���F�W��E������|� �� ��� hí% ���# h�Ɔ���E������|�0 �� ��� hí& ��� h�Ɔ��`��Lhâd� �í' ���d�0 �í( ���F��s�&�=�%�@�s�&�%� �s�.ڊ


i��	� ���ڽ@ ���	�0 ���ڽ= �����s��`
i�����i ����L���������R����H��H�� �����0��������1��� A©` L����h��h��`�נ�r��נ�� ��r����@L1� é����
���@��� ���@��0��#�'���������i(������i`�����i`������`Pause �+���)��`� �ɜ+��i(���i@� �âP� �Ʃ����O����� 4ĥ�)�����)����+L�Ɔ���� �������



����8�Jm�H8����i8�Z �å�i�ڠ  �� 9Ʃ����  ��hi���L4�		 ��* ��* ���( ���) �C��D` �­D�`�C��D�( `�CJJJJ��
)}�����	��( `�E�F�G`�$���$`����$`���(�$`�(��#�(��)�$`�L���(�#`L���#���#`����#`���(�#`�(��$�(��)�#`�L���(�$`L���#�$��E�&�&�	���
�%��L#�`�#�$��E�%�%�	���
�&��L8�`��F�(�(����G`��F�'�'����G`Deuce �$�(��#�(����M �� �L�Ƣ8�@ �à@�O 9Ʃ���@�O �Ǣ@�H�C �Ģ@�h�P �ĭ$�	�p�H <��.��	�`�H A��!��	�`�H K���(�	�`�H U���p�H _��#�	�p�h <��.��	�`�h A��!��	�`�h K���(�	�`�h U���p�h _�L��Z���,����,���,��������,�)�*�+`�0L�ĩ1��5�	��3��0�	��4��0�	��AL���Z�	H� ��h�zhi��L�� U���� _�L�� ��L�� U���� _�� �� �� *��x
��� ��E�a ��G�� �ɢʠ��G��(�ʠ��"�F��ʠ����ʠ���ʠ��E���ʠ� �� � �� 3��F�
�&m%J�	 ��L!�LS�`�rI�r`� I� `�8��`����ٙ-�#ٙ>��)�*�+�
�i���h��X���W�֍R���Q�׍c�h�b�Ía��`�ÍP��O�؍V�F�U�؍g���f�2�������r��`���  � ���#  zé����& ��`��� � ��  ��� t ���`��u� �M�