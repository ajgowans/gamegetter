                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �???�? ? �?0��?�  ��?� ��         <0??�? ? ?0?0<<?0??  0??���         ? ??�? ? ? �0?0? ??   ?�����         ? ??�? ? ? �0? ? ??   ?�����          ? ??�? ? ?0�3? ?0?   ?���?�?          ? �?�?? ? �?�3? �?�   ?��3?��          ? ???? ? ?0�????0?   ?0�3���         ? ???? ? ? �??<? ??   ?0�3���         ? ????0?0? �??<? ??   ?0�3���         <0????<?<?0?<<?0??   ?0�3���         �????�?�?�?<��???   ?0�3���                                                PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                                                                                                                                                                                                                                                                                                                                                    �����                                 �W�����                               |��VU���                             ���jUUU����                             ��kU@UU�U�                            |�ZU@UU�W�>  �                        _�VU P@U�^U�  �?                       �{�UU PU�_U� ��                      �U@TU�~UU ��                      ��U@UU��UU? ��?                     �W��UPUU��UU? ���                    �U�UPAUU��UP= ���                �   |�W�UUUUUU�~T�?����                0  �zU�UUUUUU��~5����               0  �U�UUUUUU�WA�_=����               ��   _U��UUUU��P�����               �   [U��_UUU���^�����               � ��[U��UUU��A�� ����              ���Z�
�UU��WQ�V:   ���            �  ?��/���U���W��n>    ���               �?�����U���    ���            0   ���߯���UPi��       ��            0� ? 0?�U���_PZP�       ��            � < ?�~U��W U�?       ��             0 ?��WUUU P�V�        �               ?�|UUUUUU���        �             �  ?� WU   UU��?         �             <  ?� kUUUUUU���          <            � �� ��UUUUU��          ?           �  �� ���������         �           ?   �����������          �          �����  �< �������           �               �� �  �����                           0���  ���                            ��                                     � ?                                 � �   �                �               0��   �               �               ��              ���               �                ��               �  �             ��                �   �                                    0                                     0                                    �            ��                       �                                                                                                            �����������������������������������?    ����UUUUUUUUUUUU��UUUUUUUUUUUU���?    PUUUUUU��_�uu���������U�_U�UUUUU    PUU���WUUUUU��_������_U��UUUUU���UU    PUUUUUUUUUU�U�_����_�_UU�UUUUUUUU    ��_UUUUUU��UU�_�}]��U�WUU��_UUUU��?    �����������������������������������?    PUUUU�������U�}��]]�UU������UUUU    PUUU������_UUU_����}_UUU������_UU    �����������������������������������?    ��WUUUUUU����_�_���W�_����UUUUUU�?    PUUUUUUU���������_��_�������_UUUUUU    PUUUUUU�����_���_U�_��_�����_UUUUU    PUUUUU������U�_��WU�U�������WUUUU    PUUUU������_��W��WU��U��W������WUUU    PUUUU������U��U��UU��W��_�������UUU    �����������������������������������?    ����UUUUU��U�U���U��_U��WUUUUU��?    ���WUUUUU��W��U���U��U��_UUUUU��?    ��WUUUUU���U��_U����U���U���UUUUUU�?    �_UUUUUU��_U��WU����UU��_U��_UUUUUU5    PUUUUUU���UU��UU����UU��U���UUUUUU    PUUUUUU��U��UU����WU���UU��_UUUUU    �����������������������������������?    ������_U���WU���WUUU���UU���WU�����?    ������UU���UU���WUUU���WU���U�����?    �����_U���U����UUUU���_U����UU����?    �����UU���_U����UUUU���UU���_U����?    ����_UU���WU����UUUU����UU����UU���?    ����UU����UU���UUUU����UU����WU���?    �����������������������������������?    PU����UUU���UUU������UUU���UU����U    PU���UU���UUU������WUU����UUU���_    P����WUU���_UUU������WUU����WUU����    P����UUU���WUUU������WUUU���_UUU���    ����_UUU���WUUU������_UUU����UUU���?    ����UUU����UUUU������_UUU����WUU���?    ���UUU����UUU�������_UUU����_UUU��?    ���WUUU���_UUU�������UUU����UUU��?    ���UUU����_UUU�������UUUU����UUUU�?    ��_UUU����UUUU��������UUUU����WUUU�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ����?� ��?��� �?                 300    300  �0                  300    300  30                  �����  � �0  ��                  0 0   �30  30 0                  0 0   30  �0 0                  00���  � 300  �?0                                                                                                                                                                                                                                                                                                                                                                                                                             ����|U=\�5��6��6��6\�5pU��      �? ����>�U>�U>��>���� 0 0 ��?������?����?�? � ����?��? � ����?��?0� ��� ?� ?0� ����<<� <��? ����<0�  ��? ����? �  ��? �����? ��?��� ����? ����� ����<0��<���?��<<��<��?�� ?��< �<?���?�?�< �<<���?�?� ���?��?���                �?� �?�?������ �?�����?��������?����?�?�� ?����?�?��<<����?�?��<0����?��� �? ����?��� ��? ��� ��?��3 �? ����? �3 �<0����? � �<<����? � � ?���� � ��?���?� � ��?��?�?�  � ����?�                                              �        ��  <0��0   �?<   <��0����<   ����+?���?  ��Z��� �WW�?   ?� � ? ��   ��.<��<���  � 0��� ��  p��� :�@v  p���}��@�  pg[@U@���  p��p ��  �{�     @�  �z��
 �3p�  ���? �p�3  �L �� 3? 1�3  �< �� 0<�3  ��3��   ��3  ���� �  �3  ��� �����0  0?03��"���   �    
��   ���� �b
��  ��0�� � J�?  �0�! �H��  �̴ � �3@�  o 0�   N �  � <0 " �< � �  � �   3�0���0� �� �� 01
 ��L0  k��* �����  o3Á���B���  ����   �@O�  ��p   �pg?  �kq<�(<0M�  ��|� ��0=�   ��3���0��   ��>�� ���  ����� �0��   �?0,� *8��   �Ͽ       ��   3� ��T� ?�    ���/��0��   ��0 �� ��  � �+<<<� �  �[�?<�?���  ��0   �p�   ��  < 0 ��    �0>   ���   ��Z�� ��Z��   ����< <3��3   0����������  �  �   00?   � �� 0 0       �             �                                                                            �                            0   �     3        � �  0        � 0 0��     ��3��:    0���<�?��    ����� ���     _AU<UA�0      l� �9�      �|t �=�     0�0 @A     0?<�   3<�    �|� �4=    <U  �<3  U<    ����0��    �4����?��    3 ��(�� �    � �� �    ? ���
�� �     ,
 �8 40    �O������    �|͋� "�s=     s� � �O�      ��   �3      0� ��@     �?0�  �      � �   0  ��0�    ��   1�� �L4      ���  ��      ��" �"     �� �(�(� �    � ���� �    � ��(�� �    � �� �� �    ���33����    ��� ��    ��<� ?<�    �0 A 0�3    ̜ A� 63    0� A�A� >    �� �0    ��PW��c��     <<�>��<<       ��?���       <3� ���<     ���  ��      0  0        ��   0   3        0    0    �    0                 0         0                                        0    ���0  �   �   3   ? �    ���    0   0  0   �00< 0   ���   �  "� 0�  �         �      0 � �   � 0  �  �  � < <   3 0      ��    0        0            �  0 �   �� 0�  �   3      0 �         �   �        �  0 0  �         �    �3      �              0 � 0�     � 0      �        0            � �0 # ��  �         0 �  0�       0  0     0  �  0� 0    3     � 0   �      � 0     �  0     �          �       ��     �   0  �     �  0   �     �   �  < <�    �   0�   �  �           ̀     �  3  0     0          0     � � �0  0  ��    0          �0�    � 300� � 00 0�    �  0      �  0   0 0�   �      ��        0� �                 0   �� 0 0     � � �� �   3   �0 � ����  � � �   0       �     �  �0 0   � � 0     �0         � 3     �H�Z��)�J �K �@��l ��L ��H ��I � �� ���� �� �\ �� �[  ��� �r� V��� ���� ���� �� �� �\ �� �[ ��L ��I  ���� �� �� �\ �� �[ ��I ��L  ��� �D� V逹 V� V�� �\ ��I �� �[ ��L  l�� i�� �[  ��� �[ ��L  l�� 8��� �[  ��� �� V逺 ]� �� t�2 V�� ��z�hL� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         U�WU�j�������W���W���_���_��5\�����p���s��=|���_��UU�몪��UU�UUUU몪�����U������������ |��\��0\��_���W��UU��UU�몪��UU�UUUU몪�몪��UU��UU���U�����������������U��UU��UU��UU�몪��UU�UUUU몪�몪��UU��UU���W��_��0\��\�� |�������������U������UU�UUUU몪�몪���_��=|���s��p�����5\���_���_���W���W���W��j����W�UUUU몪�몪��UU��UU����������5��50��= �����������W���U�{����UU�UUUU몪�몪��UU��UU��U�������?3��?3������U���UU��UU��UU�몪��UU�UUUU۪�������sU���W����������= ��50��5����������UU��UU�몪��UU����W���^���z�UUzoUU�oUU�o�j�m��ym��ym��ym��yo���o���o�j��UUz���_ � �p����=Wss5[ss9[9�{�5�v�5���9�U�9ץ�5�V�5�[�9[�9Wp5��?���\��l���lo��\[��\�Z�lWU�l�_�\۝�\���l���l���\���|�����? �   �?�*�	�	�*�?    �\>�:���   ����:�����:������?��������\�\�\�\��?��o���n���n���������𬪪?���?� ����������>������������� ��� ��� 𬪪?���?��p������_3����������  ����5\��:���?���0󬪪?�����p�����0���ϟ��������0�����p��𬪪?���*
  �  �  ��P�����P��:��:��
���  �
  ����*������������������������������������������������������������������������������������������������� ����=��5�z�5���5W_}5�W�7w�u7���7WWu5�_�5���5�z�5��5���=� ����<�U<0 ( �+������ pD�@2 �� ��' ڧ   � �� ��� @2�p�����+ �0 ( <�U<���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                                                                jUUUjUUUjUUUjUUUjEUUjEUUjEUUjEUUjUUUjUUUjUUUjUUUjEUUjEUUjEUUjEUUUUU�UUU�UUU�UUU�UUQ�UUQ�UUQ�UUQ�UUU�UUU�UUU�UUU�UUQ�UUQ�UUQ�UUQ�UBUR��URZ��RYZ���R�% R�%U�@&U)J�Vi%�R�% V%%UV
)UjRI��R��VRURV�h	��)���* �

*Z)�&���)���
�����  �	��X�%�X�%���*� � (�� Z���V�  TP @ U     PPP@    @     @ UP @A  P     P@% �P	 ��P�  T%  �
P  T  � % (T% T%T �
T%  T%  T	P	�U	  �   UU  UUU  UU  UU  UU  UUU  UU    UU  UU UU  UU  UU  UU U  U  TU PU @U @UU@UU PU @U  UU  U @U PU@UU@U @U PU  TUP� d� T�  �    @  d� T�*����� ��
 �� **  �* U  @Y �@��"����������ڿ�oY����U��U���Z���V������VU��U��V��jUU�V�U���i�Z�f������������j��������i������U���VU��jUU�������V�jU��U�Z����������������U����������V����j���j�j�j�j���������������������������������������e��j�j�Z�j�U�������U���j������ߪ����������������������� �� ��  ����V
��e
 �Y�@j�� �fU@��� ��Z @�f�f��J ����j��ffU   �  �
@�)  �&  �* ��** ��  �  �  �   �A  � �� j�
��U����ffUZV���jjeY����UVZe�iefZ���������F������ �*  @ @         Y���Y�ZVee�iYVeYi�Z�Vf�iZUf�jf���������
���B ��  �            UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUUUQUUUQUUUQ�UUQ�UUU��������������UUU�UUU�UUU� U�EUU�UUU�UUU�UUU�UUU�EUU�EUU�EUU�EUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU U UUUUUUUUUUUU������������������������UUUUUUUUUUUUU U UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQ�UUQ�UUQ�UUQ�UUU�UUU�UUU�UUU�UUQ�U P�UUU�UUU�UUU�������������jUUUjEUUjEUUUEUUUEUUUEUUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�����UUU�UUU����|UUU|UUU����|UUU|UUU����|UUU�UUUê���UUU�UUU��������UUU�UUUê���UUU=UUU=���>UUU=UUU=���>UUU=UUU�����UUU�UUU����>�fff�����fff�����fff����י���fffי�������fff�����fff�����fffי��fff>����fff����>fffי�������fff����י���fffי��>fff�����fff>���� � �U��_u]�U���U�UU��Uu� U�� _�5 ��/ U�������  �������  𪪪���  �몮���?  �������: ���������?������߯��������߫����ww�ݫ�����ww�ݫ����z����^UUUU��>��WUUUUժ:��U���ZU�:�����������U^UU�U����WUU������U�_UW����UUUUW����wU�Uݪ:��_UmyU��:��Wmy�ժ:��WUmyUժ>������ת����p�ת�����_�׺>����UU�ת�����UU�ת����UUת���WUU�պ��gUUUU٪���WUUUU��? k�������  kf������  kffUU���  offUU��9  lff�j��9  lff�o��9  ���:���:  ���?����U             �� �g�pկlU�>lU�>�U�>�U�>���?���?���?����� ��  �  0      �� �g�pկlU�>lU�>�U�>�U�>���?���?���?����� ��                                                                                                                                                                                                       ��      �     ��      �>     ��    ��?     <�    �<     �    �0   ��    ��� ���      �> ��5      \��� ���      ��� ��      �>� �      p�� �_      ��� ��?      �V_� _���      �o5 ��?�������   �������V�     W�������j�     ���������     ������{��    �zU��VU��U�   �����VU����   �����VU����6   �����VU�����   �����VU�����  ����U�VU�V��V p�����Z�����V�_eU���j�j��UV�WYUe�Y����gUY=�VVU�UV�jUVYUY=��U`U�UUUU��Pe��fXUUU�ZUUUBe��ZVUUU�hUUU	�������_P�������V����B���Z�ꫪ������
���������������������_UUUUUUUUUUUUU�ך�隮隮隮��7������������*����������������7?���?���?<�7SL1�SL1�SL1��SL1�SL1�SL���?���?���?��|�������������=�UUUUUUUUUUUUU��������������                                                                                    �             �        �     �        �     �        �   ��        l   �9        l9   l9        ��   [:        �� �Z>        �� �V        �V: ��        �Z� k�        �Z��Z�        �Z��Z�        ����W�        ��U�U�        ������        ��_U��    ���/�UT�����W����UUUUU���V�\���/EUUUQ���V5pU���UTUU���U�U��/0UT��jU W��o@UT��Z�  W��/  U  ��V�  \U�/�  ���U5  pU�+�����U  �W��������   _��������    _���� �����    ����������?    ����������?   �������W����*  �����������*  [���?�����[� ����?�����������_���
������������������w����������������������������_���� ��ϳ���������  �����������?      �����          ����          ����:          ��ÿ          ��ë          0���          ���           ���            ��            ��             �              <                                                          ��            ��            ��            �}?          ��U��        ��|U=W        _���W�        W�_U�_�       �U����_U      �U��U3_U      �U��U3_U      �U��U3_U      �U��}3WU      �U����WU      �U��U3WU      �W��U�W�      �WUUUUU�      �WUUUUU�       WUUUUU�       �_UUUUU�   ����UUUUU����?����UUUUU����:����{UUUUU��ꫪ���WUUU�竪�ꫪ��[_UUU�嫪�ꫪ����UUU﫪�ꫪ����_U�_�������������?����?LDD�������_1�ַ���ޗGDD4LDD�Z�   n�1�k�����GDD4������   �����>�UUU�������UUU �UU������zUU�  �_U��   �zU�  p�������/�j  |U�X�����%�U=  \UX����_%pU5  \U�Z����W�~U5  \�UU��ZUU�_5  \��UU% XUU��5  ܾ�WU��ZUի�7  ���_UUUUU���>  ��:������?��:  ��ʣ�����ʣ�>  ��ʣz�<�ʣ�?  ��:�~���:��   �^��z���    ���W�����     ���������      ���?��?�?                                                                              � �T  i歎 �[ �� �\  ����T `Z�
��W��e ȹW��f ���G i7�ez L�`H�Z�
��W��e ȹW��f ���e�d�8�7�G z�h L�`H�Z8�7�N �G �a��d��N ���G ��d�G ��A8�7�G ��a�G h`H�A8�7�N �G �a��d��N ���G ��d�G ��Z8�7�G ��a�G h`��� ��U �)��_ ��� �@�l �� �t �u �v �w �x �y �z �{ � �d�| �� �� ����$�| �� �� `�J �K �L �O �� �"�!�4�� �*�+�,�� �V ���'�� ��� i�� �� �� �� ���� 8��� �� �� �� ��� ��� �� �� �� �5�6�7�8�9�:�;�<�=�>�?�@��� �� �� �A�� �E�F�B�C�D��� ��-�/�3�1�(�0�2�C����������	��
��������������� �#��$��U ���������l ��� �� �_ �^ �� �Y �� �� ���F �j �k �� ���
� ��`H�Z J� ]� ���� ��� � ���� ���  Qܩ� �ܩ�-�3�� �%�U �#���� ��� �� �� �� �� �_ �^ �� ��` �  ��	 L� J�L����  ;� ,୮ �n �� {� o� �� ��ή ή �� �_ �^ �� �<� m� f� L�z�h`H�Z�o �{ 0N��n �z 0D��m �y 0:�o �x 0P��n �w 0F��m �v 0<�o �u 0J��n �t 0@��m �s 06��I �� � 4��d� �| ������� �- Z��d� �� ������� � �� G��d� �� ������� z�h`�m �n �o `H�  ���� V�h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<3<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���*      �?�?      ��������ȥҥܥ�������"�,�6�@�J�T�^�h�r�|�������������¦̦֦���������&�0�:�D�N�X�b�l�v���������������ƧЧڧ�������*�*�4�>�H�R�\�f�p�z���������������ʨԨި�������$�.�8�B�L�V�`�j�t�~�������������ĩΩة���� �
���(�2�<�F�P�Z�d�n�x���������������ȪҪܪ�������"�,�6�@�J�T�^�h�r�|�������������«̫֫���������&�0�:�D�N�X�b�l�v���������������ƬЬڬ������� �*�4�>�H�R�\�f�p�z���������������ʭԭޭ�������$�.�8�B�L�V�j�j�t�~�������������خخخ���� �
���(�2�<�F�P�Z�d�n�x���������������ȯүܯ�������"�,�6�@�J�T�^�h�r�|�������������°ְ̰���������&�0�:�D�N�X�b�l�v���������������Ʊбڱ������� �*�4�>�H�R�\�f�p�z���������������ʲԲ޲�������$�.�8�B�L�V�`�j�t�~�������������ĳγس���� �
���(�2�<�F�P�Z�d�n�x���������������ȴҴܴ�������"�,�6�45454545,,,,,,,,--------------------,,,,,,,,,,,,,,HIHIHIHILMLMJKJKLMLMJKJK,,,,,,,,,,LMLM---JKJK---LMLM---JKJK---LMLMJKJKLMLMJKJK---------------------------45--------45----4545BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBLMLMLMLMJKJKJKJKLMLMLMLMJKJKJKJKBBBBLMLMLMLMJKJKJKJKLMLMJKJKBBBBBBBBBBBBCCCCCCCCCCCCCCCCCCCCCCCCDDDDCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD----DDDD----DDDD----D,,,----D,,,CCCC,,,,CCCC,,,,CCCC,,,,CCCC,,,,CCCCHI,,,,HIHIHICCBBCCCBBBCCCBBBCCCBBBCCLM,,JK,,LM,,,JKLMLMJKJKCCCCLMLMCCCCJKJKCCCC----CCCC----PQPQNONONONOPQPQPQPQNONONONOPQPQPQPQNONONONOPQPQPQPQNONONO,,PQPQPQ,,NONODDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCLMJKLMJKLMRTTVJKSUUWlklklklDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDfTTe---dUUg---------------,,,,,,CCCBBBBBCCCBBBBBCCCBBBBBCCCBBBBBCCCBBBBBBBBBBLMLMLMJKJKJKLMLMJKJK,,,,,,kl,,,kRTTTV,,SUUUWl,kl,-----,kl,-----,,-----,,-----,,--BBBBBB--BBBBBB--BBBBBB--BBBBBB--LMLM--JKJKLMLMJKJK,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD-----------BBBBBBBB--BBBBBBBB--BBBBBBBB--BBBBBBBB--BBBBBBBB--BBBBBBBB--BBBBBBBB--BBBBBBBB-----------,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,kl,,,,,,,,kl,,,,,,,,,,,,,,,,,,,,,,,,,,,,LMCCCCCCJKCCCCCCLMLMCCCCJKJKCCCCDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD----DDDD--------CCCCCCCCCCCCCCCCCCCCBBBBCCCCBBBBCCCCBBBBCCCCBBBBCCCCBBLM,,,,JK,,,,LM,,,,JKLMLMJKJKCCCCLMLMCCCCJKJKCCCC----CCCC----NONOPQPQNONONONOPQPQPQPQNONODDDDPQPQDDDDNONODDDDPQPQDDDDNO,,DDPQ,,DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDklklklklklDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD...LM.JK.LMLM.JKJK..RTTV....SUUW..k.lk.lDDDDDDk.lDDDDDDD.lDDDDDDD.lDDDDDDD.D...----.----.----.----.----.----.-.-.-CCCCCCk.lCCCCCCCk.lCCCCCCCk.lCCCCCC.lCCCCCC.lCCCCk.lCLMLMk.lJKJKk.lLMLM.JKJK..,,,,,.,,,,,.,,,,,.,,.--,---,,---,,--,-,---B---B--BB--BBB--LMLM-JKJKk.lLMLMk.lJKJKk.lk.l,,,,,DD.l-,,,,,DD.l-,,,,,,.-,,,,,,.-,,,,,,.-DDDDDD.DDDDDD.DDDDDDk.lDDDDDDk.lDDDDDDk.lk.lk.lCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC����뺮�뺮�����iUUeiU�ei��g�?3g�?3gi��giU�eiUUe����뺮�뺮���������뺮�뺮�����YUUiY�Ui��i����������iY�UiYUUi����뺮�뺮���������ۺ�����������\U%8�U%��%h?�%h�%h�%h�%h=�%����뺮�뺮���������뺮�뺮�����X|)X�p)X3p)X�)X�)X��+XU?,XU5/�������뺮���������뺮�뺮�����h=�%h�%h�%h�%h?�%��%8�U%�\U%��������ۺ����������뺮�뺮�����XU5/XU?,X��+X�)X�)X3p)X�p)X|)����뺮�뺮����������z����������h�W%h�_%h�_%h5\%h�%hp%h�s%h=|%����뺮�뺮���������뺮�뺮�����X=|)X�s)Xp)X�)X5\)X�_)X�_)X�W)����뺯��z������UUU�UUU�UUU�UUUUUUQUUUQUUU@UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@UUUEUUUEUUUUUUjUUUjUUUjUUUjUUUjUUUjUUUjUUUjEUUjEUUjEUUjEUUjEUUjU jUUUjUUUjUUU������������������������UUU�UUU�UUU� UP�UUQ�UUQ�UUQ�UUQ�UUQ�UUU�UUU�UUU�UUU�oUUUoUUUoUUUoUUUoEUUoEUUoEUUoEUUoUUUoUUUoUUUoUUUoEUUoEUUoEUUoEUUUUU�UUU�UUU�UUU�UUQ�UUQ�UUQ�UUQ�UUU�UUU�UUU�UUQ�UUQ�UUQ�UUQ�UUQ������������VUUUUUUUUU�VUUUUUUUUU�VUUUUUUUUU�VU�W]]��_�VU]��]�U]U�VU]��]�U]U�VU���]]�W�VU]��]]�]U�VU]��]]�]U�VU]�����_�VUUUUUUUUU�VUUUUUUUUU�VUUUUUUUUU�VUUUUUUUUU������������                    ����          �����         ������        ���U���       ��UUU��      �UUUUU��      �_UUUUU��    ��UUUUUUU�� ���UU��_UU�����UU= |UU�����UU��UU���?���WUU]�uUU��>l��WUUW��UU��W9l��W��U�U�W��W9|��W�oUUU�_�W_=��U�jUUU�U��;o��U�VUUU��U�
���կVUUU��W������oUUUUU�_�_�o�w�oUUUUU�_�_�o���oUUUUU�_�[�o���oUUUUU��[�o���kUUUUU��[�o���[UUUUU��[�o���[UUUUU��_���[UUUUU�����w�[UUUUU�����u�[UUUUU�]+���w�[UUUUU�_���_�w�kUUUUU�_��[�կU���U�W��[�տ֪ת��W�{�[�U�ڂׂ��U�{�[�U��ת�U�{�[=|U�����_U=|��U������WU����>|UU�����UU=�����UU��ז�UU��>�ϿUU��זUU��?��VUՖזWU������[UՖזWU� ��[UՖזWU�  ��kUՖזWU�  ��kUՖזWU�  ��kUՖזWU�  �Z�U����WU��  �k�U����WU��   o�VՖזW�~�    ��ZՖזW�_�    ��k����W�>    �Z�UUUUU��    �k�ZUUU�~�     ���UUU�_�      �V�UUU��>      �j����^�      ��������       ��?����        ��   �         ����     �v �y �w �z �x �{ � �� �� ����`�s �v �t �w �u �x � �| �� ����`�m �s �n �t �o �u `�m �v �n �w �o �x `�m �y �n �z �o �{ `H���T ��� �d�� �u )�G  ��t  ��s  ���� �n�� �x )�G  ��w  ��v  ���� �x�� �{ )�G  ��z  ��y  ��h`H���T ��� �d�� � ���� �n�� � ���� �x�� � ��h`H�Z�� � �L�� ؽ m���b��� � �d�G  L��]���  8� V� V� V� �� ��  ������� �� U������ ՙ U����� U��8��� L�� ���� u���� L�����  u���Е U�����  u�L.�z�h`���?�;l9�:,8    �?�5�6�:�>     ��>`�`��>�     �>�:�6�5�?    ,8�:l9�;�?��  � ���:\>�  ������=WUU5��_=�V��U9 p���p�U�p����U9 �V���_=WUU5���=���        ����|ZZ�\UU�|����� lU��gwUg��g lU��|���\UU�|ZZ������W�U���_���z[UU���W��%[���[��Z��Z���[��%[���W�[UUꫪ�z���_�W�U�?�������������? ��?�;�;�����?��pp��>�?0   ���ة��  ��� � �P � � �Q � �ߍ& � t ����< ��= �� � �<����= ��� J�XL �H�Z�W �X � ��X �/ ��/ � �� ��(z�h@H�' )�	�W �Z �# �$ �% hX@                                                                                                                      ���T  � J� X�  ��Lԥ� �� u�@�l �  �� J� z� ���  �� u���	��#�l ���F  ݛ u� L� b� B� X�  �� J� Y� j� J��� ��� � ���� ���  Q� �� ;圹 ��U  o�ή ή ή ή �� �_ �^ �� �x֜� �_ �^ �  �� L� f� m� �@�l �  ��L(� -� �� �٭4��� 4� �� .� ,� X� �� U� �� t� {� !� �� �� R� �� %� Q�L��H�� ɑ� �� �魼 � ����  �� �魼 � ��� h`Hک�� �P�� �� ������,��9��F�V�
 ���`  �©�B� ���`  �©�1� ���`  �©� � ���`  �©�� ���`  �©	 ���h`�
�� �<�� `HZڭ  	����2 V� V��� �� �� �A�B�C�D�E�F�#�� �� �  	���� �ȭ  	���� bĭ  	���� �í  	���� Cŭ  	���� ƭ  ��� �� ���zh`H�Z t歭 �[ �� �\ �J �K �#���$�L �&�%�	�U �L �% ��z�h`HZ�#���# �í� ɐ� �� �魼 ���� �� �� ��zh`Hڮ$����U �K����U �@����U �5����U �*����U �����U �� ���U �	�!���U �U �%�� �� �A�B�C�D�E�F��� �h`HZ�#���# �ĭ� �0=� �� �魼 ���� L��ή �� �孮 �P  �� �魼 ���� ��� �F��� ��� zh`Hڮ$����U �K����U �@����U �5����U �*����U �����U �� ���U �	�!���U �U �%�� �� �A�B�C�D�E�F��� �h`H�#� ���# nŭ� �0 �� �ꭼ ���έ h`HڮU ��� �$��&L�����!�$��&L������$��&L������$��&L����� �$��&�.���!�$��&�����$��&���
��$��&�� �� �A�B�C�D�E�F��� �h`H�#� ���# @ƭ� �$ �� =ꭼ ���� h`HڮU ����$��&L������$��&L������$��&L������$��&L������$��&L������$��&�����$��&���
��$��&�� �� �A�B�C�D�E�F��� �h`H�Z�%��.�� � �	 �� ��L���� J�L���� ��L���� �L����.�� � �	 � H�L���� ]�L���� ��L���� !�L����.�� � �	 1� ��L���� p�L���� ��L���� .�L����+�� � �	 P� "�L���� ��L���� ���� ;�L����.�� � �	 o� ��L���� ��L���� ��L���� �L����.�� � �	 �� ��L���� ��L���� ��L���� !�L����.�� � �	 �� m�L���� ��L���� ��L���� .�L����-�� � �	 �� ��L���� ��L���� ��L���� ;ˀ�	�L��z�h`H�Z�� �� ���  ���� �� �A�B�C�D�E�F�� z�h`H�� i�� ��� �� i�� ��� �� i	�� ��� �� i�� ��� h`H�� iʹ ��� 8�� �Ͳ ��� h`H�� iͫ ��� 8�� �ͬ ��� h`H�� i�5��5�� i�6��6h`H�� i�7��7�� i�8��8h`H�� i�9��9�� i�:��:h`H8�� ��;��;�� i�<��<h`H�� �=��=�� i�>��>h`H�� �?��?�� �@��@h`HZ�� ��M bέ�L �� �[ �� ��� �\ ��  Eέ��# ��ί ί �� � �� ɐ��� �ѭ� � �� �� �� �� �� �zh` �� �� �� �� � H�` �� �� � H� 1� ��` � H� 1� �� P� "�` 1� �� P� "� o� ��` P� "� o� �� �� ��` o� �� �� �� �� m�` �� �� �� m� �� ��` �� m� �� �� �� ��` �� �� 1� �� o� �� �� m�` � H� P� "� �� �� �� ��` �� �� o� ��` � H� �� ��` 1� �� �� m�` P� "� �� ��`HZ�B��a bέ�L ��� �[ �� �� �\ ��  Eέ��7 ��� 8�� ��� �� � �� ɐ��� �'�� л�� �'��� ��B�� �� �� �� �zh`HZ�C��C bέ�L �� �\ �� ��� �[ ��  Eέ�� ��� �� �'��� �ۭ� �'��C�6�� �5�� �zh`HZ�D��Z bέ�L ��� �[ �� �� �\ ��  Eέ��0 ��� �� i�� �� ɜ��� �'��� �­� ɜ��� �'��D�8�� �7�� �zh`HZ�A��F bέ�L �� �[ �� ��� �\ ��  Eέ�� ��� � �� ɞ��� �ح� ɞ��A�:�� �9�� �zh`HZ�E��Z bέ�L ��� �[ �� �� �\ �� �� ɜ�3�� �0, Eέ��" ��Σ �� i�� �� �­� ɜ��� ���E�<�� �;�� �zh`HZ�� ��A bέ�L �� �\ �� ��� �[ ��  Eέ�� ��Υ �� �0
��ݭ� ��� �>�� �=�� �zh`HZ�F��a bέ�L ��� �[ �� �� �\ ��  Eέ��7 ��Χ 8�� ��� �� � �� ɐ�� �0�� л�� ��� ��F�@�� �?�� �zh`��� �� �� � K� �� �� ��`�J �K  i�`�J �K ��L  i�`H���! l� T� �� �� � D� �� �� �� �� �έ�� �ѭ�� ҭ�� 4�h`HZ�� ����!��S��+��'��5��1��H�� � T�O�� � �F�� �(0B�=�� ɠ��4�� �(00�+�� � �"�� ɠ���� �(0��� � ��� �  G�zh`��� ��� `�� ��4�� �[ �� �� �\ ��  �ޜ  !խ�� G�L���� 8�� ��� �`�� ��+�� �\ �� �� �[ ��  �ޜ  !խ�� G�L���� �`�� ��4�� �[ �� �� �\ ��  �ޜ  !խ�� G�L��� �� i�� �`�� ��1�� �[ �� �� �\ ��  �ޜ  !խ�� G�L@��� ��� �`�� ��4�� �[ �� �� �\ ��  �ޜ  !խ�� G�L��� �� i�� �`�� ��+�� �\ �� �� �[ ��  �ޜ  !խ�� G�L���� �`�� ��4�� �[ �� �� �\ ��  �ޜ  !խ�� G�L���� 8�� ��� �`�� ��1�� �[ �� �� �\ ��  �ޜ  !խ�� G�L0��� i�� �`HZ�*��L lέ� �[ �� ��� �\ ��  �ޜ  !խ���� �� ɟ��� �� ��� ɟ��	�� �
�� �zh`H lέ� �\ �� �� �[ ��  �� �ޜ  !խ��;�� ͭ ��� ��� �� ͮ �� �� �� �� ��� �� �� �� �� ���� ��� �h`HZ lέ� �[ �� ��� �\ ��  �ޜ  !խ���� �� �0�� �� ��� ���� ��� �zh`HZ�� ��^�k ̮ �@0�j ͭ �	��� �C��� �<��� �5�j ͭ �	��� �$��� ���� ��j ͭ ���� ���� zh`H���!�J �K �� �L  t�� �\ �� �[  �� ��h`HZ�� ���� i��� ����� i��� ����� i��� i����� i��� i����� i��� i����� i��� ����� ��� i����� ��� �zh`�� �� �� �� �� ���(��
��
�<�����  !�`����`����� �� �� �� ���  �� !�`������� �� �� ��V `����� �� �� �� �� �ө�  !�`������� �� ��V `����� �� �� �� ����  �� !�`������� �� ��V `����� �� �� �� ����  �� !�`������� �� ��V `�0���� �� �� �� ��  �� !�`�(���� �� �� �� ����  �� !�`����(�� �� ���V `HZ��� �� m�� �� �� m� �� �� ͸ ��� ͷ ��� mͪ �L���� m� ͖ �j� ����� r� �L�� ��� W�L������ r� �� W�L����� �L����� ��L�����  �L��� �� m�� �� �� m� �� �� ͸ �&�� ͷ ��� mͩ �L��� m� ͕ �Li��zh`H �� 2� o� �� թ�H ��I �� �[ �� �\ ��J �K �
�L  ��h`�4��L���� � r��� � �N��  �� �ש�� �� �� �� �B�C�D�E�F�� ������-�3�/�0�1�( 5ڀ�� � �T  �ܩ��T 8��� ��`��H ��I �� �[ �� �\ ��J �K �
�L  ��(`� �0�� �0�� �� `H�Z� �� �����h�i� ���� �W��� ��� ��  �܀@��V ��� �4������(�� �� ��� �� �� �B�C�D�E�F�A��V �� �� �� z�h`� �T  �ܩ��T ��H ��I �� �[ �� �\ ��J �K � r��
�L  �� u� ��`HZڭG�F�#�G�� ����	���� ���� ��2�� �� �� � 0L�؜�  ���� �� �� �� �� ��  �؜� � ��l  j� J��2�� �� �0&�$��� ��� �P�� � ��  ��� L� J�L ���V  b�La���V � r��zh`�� ��Ln٩�H ��I �� �[ �� �\ ��J �K � r� ��
�L  �� u� �� u��� i�[ �� i�\ � r� �� �� u� �� u��� i
�[ �� �\ � r� �� �� u� �� u��� i(�\ �� �[ � r� �� �� u� �� u��� i
�[ �� i(�\ � r� �� �� u� �� u��J �K �� �[ �� �\ ��H �<�I ��L �@�l �  �� r� �� u� ���L � r� �� �� ���L � r� �� u� ���L �L � r� �� j� ���� `HZ�4��D t��U �#�� �� �0�� �4��� �"���  �� o� V� l�ή ή ή ή �� ��zh`HZ�ΐ �� � 0 u�� �ܩ�� ���� ��4L`� J� m� f�  �� �� �� u� � u� J� �� uܩ8�� ���  Q� �۩��  d� tۜl �  ������� L� l�� ��
���  �ۀ]���  �ۭ  ������ L����2�� �l ��)� ��L[��  ��У L��� �����  l� �ۀ� L� l���  �ۭ  ������L�� L� J� m� f� �@�l �  ���� �)��� �2�L(��zh`�
�� �d�� �  ��`�
�� �x�� � ��`��[ �d�\ ��H �
�I ��J ��K ��L  ��`��[ �x�\ ��H �
�I ��J ��K ��L  ��`H�Z �� ]� ���[ �(�\ ��K �L ��J ��H �I �@�l �  �� ���L ��[  ��l � ��z�h`H�Z�V ��R��mm �m �n i �n �o i )�o ؜V z�h`�� �� �� �� �o )�G  ��n  ��m  ��`��� �(�� � ���� �(�� �u )�G  ��t  ��s  ��8�� ��� � ��`H�Z��[ ��\ ��I ��H �@��J �K ��L  ��%�� ��� �� �G  ��C�z�h`H�Z u� �� m� f��)��&  L���[ �F�\ ���T ��J �K ��L ��I ��H  �� o� ��  ��� L��� �ߍ&  �� ]�z�h`�� i�� �� �� i�� �� �� i�� �� �� i�� �� �� i�� �� �� �� �� i	�� �� �� i�� �� `��H �<�I ��J �K `H�Z��)�� ����(��.��4��:L>ީ
�H �(�I ��J �K ��L �& �ݩ�L � �ݩ�L � �ݩ�L � �ݩ�L �� �[ �� �\  ���)z�h`��� ��`H�2��# ���� �� �� �0Q�2���!�" `݀>� �:�!����  �ݭ� �&�!��"��"����  �ݭ� �0�"��!h`��� �� �� 8� �� ��`�� �� �� �� `H lέ� �[ �� �� �\ ��  �� �ޜ  !խ���� i�� �� �� �� ɜ��� ��� �� �� �� �h`H lέ� �[ �� �� �\ ��  �� �ޜ  !խ���� i�� �� ɜ��� �� �� �� �h`H�� ���D lέ� �[ �� �� �\ ��  �� �ޜ  !խ���� i�� �� ɜ��� �� �� �� �h`H lέ� �[ �� �� �\ ��  �� �ޜ  !խ���� i�� �� �� �� ɜ��� �'��� �� �� �� �h`H�-��= t�J �K ��L �� �[ �� �\  ���� �� �� �� �� �0O ���-��� �0� �> � �魼 ���� ɠ�
��-�� �� �� �� �� ��� �� �k �� �j  ��h`�� �j i��� �� �k i��� ���� `H�3��f t�J �K ��*�L �� �\ �� �[  �� � �魼 ���� �� �� �� �� �0#�3���� i�	�� �� i�
�� L��L��� �x � �魼 � �& =ꭼ � �c �ꭼ � �f�� �� �� i�
L���� �� �� i�	�� i�
��* ��8�� �� �07�038�� � �8�� �� ���� �#�* ���� �� �"�* ��h`H�� �LS�/��I�J �K ��L  t�� �\ �� �[  ���� �� �"5�/��8�� ���� �� i��� �� ��� �� i� �h`H�1��S t�J �K ��+�L �� �\ �� �[  ���� �� �� ɐ�#���18�� ��� ��� i�� �Ld�Lr�� �$ $� �魼 ��<�� � ɠ0ɀ0��1�Lr��� �� 8�� ���� i���+ ?�0 $� =ꭼ ���H $� �ꭼ ���I�� �� 8�� ��Lr�8�� � �0:�068�� � �8�� �� ���� �� �#�+ ?��� �� �"�+ ?�h`H�� �L
�(��L
��J �K ��L  t�� �\ �� �� �[ ��  ���L  V� �� �� �ө�� ��� ��  !թ�� ��� ���*�� ͭ ���� ��� �� ͮ ���� �� ��� �� �h`�� �� �� �� �� ��� ���  ��`H�0��$�  �� �� � !խ ���� ɠ�&��0�� ��  �� �� � !խ ����0��� ��� � h`Hڮ� � ���� �5����� �*����� ����	�� ����
�� �	����� �h`H�0��  t歽 �[ �� �\ ��J �K �� �L  ��h`H�Z�� �F0���F �� �O �� ���F �O �� �_  ;�F ɠ����F � �Y z�h`HZڭ` �J  t�F �� �\ � �[ �_ �K �^ �L �l ��) ���^ �[ i�[ �(�� �� G� oí` �J �^ �_ 8�� ��� �\ ��
а�� �zh`H�4�� �� � ?� �� ��h`�-������J �K �� �L �� �[ �� �\  ��`�3������J �K �*�L �� �\ �� �[  ��`�/������J �K ��L �� �\ �� �[  ��`�1������J �K �+�L �� �\ �� �[  ��`��H ��I `��H ��I `H��U �U ��L����L����L����L����L����L����L����L���	���U �U �%�h`H��$�$����&LG�����&LG�����&LG�����&LG�����&LG�����&LG�� ���&LG��!���&LG��"�
��&��$�h`H�Z� �< �@�= � � � �<����= ���z�h`� �T  ����T `�[ �\ ��J ��K �L �(�H ���I  �� V�[ �\ `Hڪ���




�N ��)N �& �h`H�Z�[ �a �@�b �J 
�����B ����C �K 
��B�D ȱB�E �L ��D�i �i 
��e��c �e��d �d ml �d �\ � ��a i0�a �b i �b �� �� � �b �0 �)��	�c-T �a��)��	�c-T a�a��H ���a i0�a �b i �b �c mH �c �d i �d ��I Чz�h`H�Z
�����R ����S � �R�$��a��b��c��d�8�7�G  ��Ȁ�z�h`H�Z�)�JJJJ�G  ��)�G  ��z�h`xH�Z�G �a��$��b��%��c��&��d��'�����< ����= ��M �� �Q��@ ����A �� �<-T �@�< Ȳ<-T �@�< ��M ��� � z�hX`�Z�/���� ���� ��z�`ڢ( V�����`ڢ
 V�����`ڢ V�����`ڢ V�����`H�Z�� �a �@�b �� �� �a i0�a �b i �b �� �� �a)�����a)����H �Ꜽ ���� z�h`H�Z�� �a �@�b �� mI �� �� �a i0�a �b i �b �� �� �a)����a)����H �Ꜽ ���� z�h`HZ��� i�a �@�b �� �a i0�a �b i �b ��� � �a)����!�����a i0�a �b i �b ��I �ڜ� ���� �zh`HZ�8�� ��a �@�b �� �a i0�a �b i �b ��� � �a)���a i0�a �b i �b ��I �ߜ� ���� �zh`�� �� �� ��  t�` t�� �� �� �� ` t�� �� �� �� ` t�� �� �� �� `HڮY ���-�������-�"�� �� L��� �/�������/�(�� �K�� L��� �1�������1�
�� ���� L����3�������3��� �� L��	��(����(�(�� ��� L�� ��0����0��� �� ��� �� ��F��Y �G�Y ��2��� �� �h`Hڭ� �A0LU�O �d0�O LU���0�-��&�����-�� �0��� �	�� i�� �� LU����(����(�(�� �<�� LU��� �/�������/�(�� �x�� LU��F�@�1��6���/��1�� �0� �� ��� �
��� �	�� i	�� ���� LU��H�>�3��4���-��3�� �#0��� ��� �
��� �	8�� ��� �� LU��P��0����0�� ��� ��� �� �h`� � �  f� m� � � � � � � � �: �; �ߍ& �* `H�Z� ���Q� ���.� � f� � � �  ]� � m� � � �  ��� � �	 � #�� � � � �� ���.�( � f� m�! �" � � � �  ��( �( �# � ��(z�h`� �� ȱ� ȱ�	 ȱ�
 ȱ� )
��X�� �X�� Ȍ � � �	 � �'� �6� ȱ6� � �� � �� ��Ȍ � ��`� ��! ȱ�" ȱ�# ȱ�$ ȱ�% )
��X��& �X��' Ȍ �( �) �# � �#� �  f� m� � � � � � � � `� �� ȱ� ȱ� ȱ� ȱ� )
��X�� �X�� Ȍ � � � � �'� �8� ȱ8� � �� � �� ��Ȍ � ��`H�Z�
 )?	@�+ �
 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �: �� �: z�h`H�Z� )?	@�+ � 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �; �� �; z�h`H�Z�$ )?	@�+ �$ 4��-+ �+ �) �&��% )@��J��+ �+ Ȍ) �&����) �% �) �+ � � �: �; z�h`� �: `� �; `�T�� �U��  � ��*  �� ��� `H�Z

�����6 ȹ���7 ȹ���8 ȹ���9 � �6� �8� ȱ6� �8� � � �� �  #� �� ]� ���� z�h`H�Z
��L�� �L��  � ��*  �� ��� z�h` �� � �� �� �� j� w� � �� �� �� �� �$� �� �� �� x� �� _� Y� _� j� w� � �� �� �� ��    �� �� �� �� �� �� �� �� �� �� j� w$� �� �� �� �� �� �� �� �� �� �� � j� H� j`� � w� � �� �� �<� �� �� j�    _� Y� _� w� �� �� �� �� �$� �� �� �� ���@�� �� �� �� �� ����@�h�T�� �� �� �� �� ��@�T�   }���}�@� �� Y� _$� j� w� � �� �� �� �� �� �� � j�   .�}�������:�\�:�����.�}�   ����\���\�����T��.�� ��.�T�   �.�� ��T�}�:���}�T�}����@���������   �T���}@�����������}�T������0�   �������.�T��}�}0�   �� �� :� ��    �� �� �� ��    �� \� �� \� :�    ���������f���f���������   �����������B�@�f���f�����@�   f���f���@���f����@�����@�B�B�B�B�   �@�B��@�����B���@�B����0�   f�f�f�f��f���@�f����0�    � �� �� �� �� �� �� �� �� �� �� �� ��    ����.�@�T�h�}�����������    �  _�  T�  ?�  �  ?�  �  �  �  �    }� ��  ��     �� /2�   
	 �
	�
 �
��


		�		�	�
�
��

		�
	����4�@���Y��  ��������������������������������������������  c����C��  �O�����9�  s�����0�B�  O�V�a�j�w�����������������Hڍ- �1 ���0 �h`H�Z�0 ���F�- 
�����2 ����3 �1 

��2�'�* ȱ2



�4 �5 ȱ2�/ �) ȱ24 �( �1 � ��z�h`�0 �* `���� ��
 ����.� �� ��CONTINUE$SCORE$HEIGHTa$END$YOURaSCOREa$STAGEaONE$STAGEaTWO$STAGEaTHREE$STAGEaFOUR$STAGEaFIVE$FIRSTaATTACK$FIGHTaALONG$COMEaINaSTAR$GOaFORaSUCCESS$WINaLASTaFIGHT$HIGHaSCORE$YOUaAREaVERYaLUCKY$�����+�5�?�K�V�a�n�z�����| � � ���������� ���`� ��*�:�*�:�	0123;<@A\]^_`abctu !"#
6XYZ[$%&'()*+=>?EFGhijmnopqrs  Pp�| � � 
dnxt�4�t�����t���􅀀����0�p������� �@��� �@�������;ݾ�����Ђ��Ђ��HYHZt� @$Y @ @ @ @ @ Y���4�4�ݿ� �@�t�����4�4�4�4�����ЄЄЄͿ0�4�t���4�t����4��4�t����4�t����4�t����4���0���p������� � �@�@���@����� ��f�g�h@�����H[�^Pb��,�l�M�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     J� �p�