�R�����R��ҁ����"�2�B�ҁR�b�r���������ҁ҂����"�2�B�R�b�r���������҃����"�2�B�R�b�r���������҄����"�2�B�R�b�r���������҅����"�2�B�R�b�r���������҆����"�2�B�R�b�r���������҇����"�2�B�R�b�r���������҈����"�2�B�R�b�r���������҉����"�2�B�R�b�r���������Ҋ����"�2�B�R�b�r���������ҋ����"�2�ҁB�ҁR�ҁb�r���������Ҍ����"�2�B�R�b�r���������ҍ����"�2�B�R�b�r�B�������B���B�B�ҎB�����"�"�2�B�                           � � �         � � � ���������������� � � � � � � � ��������������� � � � � � � � ����ꪪ������������ �     � � �         � � � ��o��f��gf��ff�� | � | � | � | �ff��ff��ff��f�� | � | � � � � �f��f晙ff��gf���f�� �                    ? ??��           ���ߪ����������_UUWWWUU�_�_>___||UU�U�U}UUUUUUUU||��������U]UUWWW�W�W������     ? �?������       ���ϙ?f���f��f��?    ��>?<<  � � <        <<������f��  ? ???���f����           ����                       < � �           ? < ��� � �     �� � � ?     ������ ���UU���g��g��g��gUUUUUUUU���f���f���f���g����            ���                         � �            � ����#���#���� � /�?"���?������"� � / � / � / � �����������"��#����            ����                        ? �              � ��������g��ff��ffÏ�"��>��������"��ff���g���g���g���"���"���#�������            ?��          �             ��������W�W�W�W�W�W�����������������W�W�W�W�W�W�W�W�����������������W�W�W�W�W�W�W�W����            ��?�             � � � �_�W�UU            � �            ������"���?������"�U_U_UWUWUWUW}W�����������"��"�W�_�UU_U_UU������        ? �����            �����������           ?�=�UUUUUUUUUUUU�U�=���f��}��f��U�U�UUUUUU�_����f��}f���f���o��� ?             ?�                          ���            � ���իիի���꽪���������������꿪����������������������������� �            �����U�U�V�W�o@�           ����� � � @    � ��f�}f�������f��������U�W�W�W�W�f�����������f��W�������������            ��                     � � ��o � ����k�VkUVUUU�Z�UkU[UWUWUWUWUUUUUUUUUUUUUUUU�WUWUUUUUU�WeW�We��e�������������W�UfU�UfU�UeUUZU����������ff���������       ������WU       � �"��/"��#"��#>������������>�?o#��?"��/"��?"���[�[�V��Ƽſѿ�����            ���������           �����     @@������UVU�ZkUVUUUUUUUUUUUUUUUUUU���������UUU������������������������������������������VZU��[�V�U�Uo�o���UUUUU�������UPU��S�T�T<ռ����UUU�U�������ffYU�f�UoU[UVUUUUUUUUUUUUUUUUUUUU�@��?�?�s�����U�U�U�U�T�T�SESE����������������SSSSSSSUSU    ������VUUUUU     ��?����U�U�UUUUUUUUUUUUUU�����������������U�Z�j����������������������f晙�����j�Z��������UfU��g��f���UfU��� � � � ���/UU������ff��ffU�f?�?�������ff��UUUU@�?��?���UfU�UUTUSUOU?U<U�?�����������T�T�T�R�R�S�S�S�����������������S�S�S�S�S�S�S�S            � ���?f>��e���e�             ��f���e���f��f�        ��e���?           ? ��?��f���f���ef��UfU�  ? ~ � ���UeU�UeU�UUU�UUU�������f>�>UUUUUUUUUUUUUUUUf>�>f~�~f���f���UUU�UeU�Uf��ff��                �����Ѽżż�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U�U~U~UoUoUoUoUoU     @ � � � � �oUoU_U[U[U[U[U[U � � � � � �@o�oWUVUVUUUUUUUUUUU�[�[�V�U�UUoU_U             � � � � �@��o�[�V_U��<@�_� ��_���}}}}}��}}f���f��f��f���������?A ?�QUTUTUTUPL��Ӫ���� UUUUUUUUUU�Z�V�UUUUUUUUUUUUUUUUUU�U���PU�������PUTUUU�T?UCUTUUUUUUUUUUUT�C���U�U�UUUUUUUU@U/U�U�U�UUUUUUUUUUUUUUUUUUQU �
�+�����������? � �_�z���S�S�Q�T?TUBUTU�0��3�3���0� ��     ��?<<�?�? <�?���?<<�?�? <�?���?<< �� �?�?��}U}U}U}U��}}}}}}��}}}}}}��}U�_�_}U��}}}}�}��}}}}}�_]u��w���w�}}�_f晙ff��ff��ef��UUUUTUPUPUBURUUUef��ef��ef��ef��ef��ef��ef��Uf��Uf��UfU�UfU�UfU�UfU�UfU�Uf��Uf��Uf��ef��ef��ef��UUUUUUUUUUUUUUU�ef��ef��ff��ff��UUU�UeU�UeU�Uf��ff��ff��ff��ff��WUWUUUUUUUUUUUUUUUUUUUUUUUUUUUUU"�2�B�R�b�r���������ґ����"�2�B�R�b�r���������Ғ����"�2�B�R�b�r���������ғ����"�2�B�R�b�r���������Ҕ����"�2�B�R�b�r���������ҕ����"�2�B�R�b�r���������Җ����"�2�B�R�b�r���������җ����"�2�B�R�b�r���������Ҙ����"�2�B�R�b�r���������ҙ����"�2�B�R�b�r���������Қ����"�2�B�R�b�r���������қ����"�2�B�R�b�r���������Ҝ����"�2�B�R�b�r���������ҝ����"�2�B�R�b�r���������Ҟ����"�2�B�R�b�r�����        �
 ����`�� �                                         � `  �J ���� �
                      ��        �
 ��ff��ff��ff�h��I��
��*�ff��ff��`����`����ff��  ff��ff�� �              ff�h��I��`����`�� �                                         � `  �J ��           � `  ��`��F�DD�J ����`��DDDD��DDF�DDDDDDDD�Hd!�J	 ����              �� �
                      ��        �
 ��ff��ff��ff�a��I��
`�*�ff��ff��
`����
`�*��ff��  ff��ff���ff��ff��ff��  ff��a&�)�

 ��ff��ff��ff��h&�)��
 �J@      �
 ��b�b��� ��      UU        F�DDDDDD  @	�
	 ����DDDD�Hd!�� ��F�DD�J	 ����`��DDDD��DDF�DDDDDDDD�Hd!�J	 ����              �� �
                      ��   � ` `�Z`��aIff��ff��ff��a&�)a���	 �J@      �

 ����
 �J      UU        @            UU  @PDQED          @QEDQE@      PDQEDQEDQE      UU        @                @PDQEDUU        @	QEDQE@      �
	 ���� ��        UU      F�DDDDDD  @	�
	 ��b���              b���`�� �                                 � ` `��`��V�UUUUUU�Z`����`��UUUUUU��UUUUUUUUV�UUUUUUUUUUUU��UUV�YeYe�Z	`��          @�� �J@      PDQEDQEDQE      UU        @            UU  @PDQED          @QEDQE@      PDQEDQEDQE      UU        @                @PDQEDUU        @QEDQE@      PDQEDQEDQE        UU      @                @�
 ����UUUUUUUUV�XeXe��	`��V�UUUUUU                �Z`����`��UUUUUUUU��UUUUUU �              UUV�XeXe�Z`��                   � ` `�Z`���
 ���� ��                V�UUUUUUUUUUUU��   	 	 �
	 ��UUUUUUUUUUV�YeYe��	 ��V�UUUUUU�Z	`����	`��UUUUUU��UUUUUUUUV�UUUUUUUUUUUU��UUV�YeYe�Z	`��          @�� �J@      PDQEDQEDQE      UU        @            UU  @PDQED          @QEDQE@      PDQEDQEDQE      UU        @                @PDQEDUU        @QEDQE@      PDQEDQEDQE        UU      @                @�
 ����UUUUUUUUV�YeYe��	`��V�UUUUUU�Z	`����	`��UUUUUUUU��UUUUUUV�UUUUUUUUUUUUUUUUV�Y%Y%�
	 ����`�� �      ��UUUUUUUUV�X%X%��	 �
                       �
 ���� �
                           	 	 �
	 ����	 ��                V�UUUUUUUUUUUU��   	 	 �
	 ��b�          @b��� ���      PDQEDQEDQE      UU        @            UU  @PDQED          @QEDQE@      PDQEDQEDQE      UU        @                @PDQEDUU        @QEDQE@      PDQEDQEDQE        UU      @                �`��j���b���UUUUUUUUV�Y%Y%b���	 �
       �
	 ����	 �
                                             ��        �
 ��DDDDF�!Hd��	 ���DDDD�`����`��DD��DDDD�            UUDD�H$a�`��          @�� ���      PDQEDQEDQE      UU        @                �`��j���UU        �`���`�f&��ff���j�����`�ff��ff��  ��ff��f&��ff��ff��ff��ff�bF���j	���UU              �� �
                      ��        �
 ��DDDDF�!Hd��	`���DDDD�`����`��DD��DDDD�DDDDDD��DD�I$!�
 ��DDDDDD�H$!�� �
       �
 ��b�b��� Z�                f���ff��ff��ff��   
 	 �
	 ��  ��ff��ff�bF����
 �*d���ff���j	�����
`�ff��ff��  ��ff��d&��ff��ff��ff��ff�bF���j	�����              �� �
                      ��        �
 ��DDDDDD�I$!�� �
       �
 ���� �
                                                          
 	 �
	 ����
 ��                d���ff��ff��ff��   
 	 �
	 ����              �� �
                        �.�>�N�^�n�~���������Πޠ�����.�>�N�^�n�~���������Ρޡ�����.�>�N�^�n�~���������΢ޢ�����.�>�N�^�n�~���������Σޣ�UUUUUUUUUUUUUUUUUU�U�U�W�_U�_UU�_U_U�_U_U�UU_U_U_U_U_U_U�UU�_U_U�_U_U�UU�__}_U_U_U_}�_UU��W�W�W�W�W�WUU_}��}_}_}_}UU�__}_}_}_}_}�_UU�W___}_}_}__�WUU�_U_U�_U_U�     � ����������������������ެ��������� ��UpU��    ��UU��  = � � ��UU��uUUUUW�]UW_U�UU��     � U�������=U�_�u�U=UwUU�?W���                    ����0��0�                       ������� 0 0 0    0 �������_�U�UpUlU�����ijiZ�Z����   � � �������UUUUUUUU}U��  ? � �����<� �< ���?;�>�?��?UUU5�?   �  � s s s s  ��  ��UUUUUUUU�p�p�p��� �0��� }}}}}}��    ��  ���0 � ��|UWU��      ��_5\�  ? � � � � � � 3 ?�� � �?� � �U=U���     ��D0�p0p�0�p�0p�0pG<=w�7wL<3pL0���?    ��DD� p 0<p     � ����<0<p 0�ODt�D��� ����>w�DD1DD�D<� �w�w��?�� ? ���UU_}_}_}�_}_}_}UU�_U_U�_U_U�UU�__}_U_U_U_}�_UU_}__�W�U�W___}UU�_U_U�_U_U�UU�__}_}�_�W___}UU�__}_U_U_U_}�_UU_}_}_}_}_}_}�_UU_}}�}�__}_}UU�__}U}�_U}_}�_UU�__}_U�__}_}�_UU�__}_}�U}_}�_��������ʥڥ���
��*�:�J�Z�j�z���������ʦڦ���
��*�:�J�Z�j�z���������ʧڧ���
��*�:�J�Z�j�z���������ʨڨ���
��*�:�J�Z�j�z���������ʩک���
��*�:�J�Z�j�z���������ʪڪ���
��*�:�J�Z�j�z���������ʫګ���
��*�:�J�Z�j�z���������ʬڬ���
��*�:�J�Z�j�z���������ʭڭ���
��*�:�J�Z�j�z���������ʮڮ���
��*�:�J�Z�j�z���������ʯگ���
��*�:�J�Z�j�z���������ʰڰ���
��*�:�J�Z�j�z���������ʱڱ                     � � � �󯿪�����������������������:�����������������������������������@    @ @ P Tϫ=�����Z?j=��������������      = 5 � � � � � � ? � ��          ���������� UP�T���_x�Z�j��Z������V[�������������         � � � �𯰪                  �������������  U_U�U�_<������VW��W���������������                                    ���������������   < < <�� � ��?���������ǪǪ��  �  W?�             � � �U=��    ������������ � � � � � �         � �?��1qqqq�s�s�<<��� � ���           : ��    ������������     � � � � | |��� � � � <     � ��_�|�|��Z���������j�꼪���Z���� � ��������������������� � � � � �             ��������������� � � � � �        ��??�_<����������                                           �?�ꪪ����_U_UWWUE        _ _�W�W�U|E_                 ? � ���U��y��V�����j���������������������  ��\U\U|�p5p�pU  �U5U55p55U5pUp�p5p5p5p5�  U5WWWW5\5�    ��pU\U\�\\\  �UU5_5p5p5p5\\\\�\UpU��  p5p5p5_5U5U�    �\\\\\\  �?p5p5p5p5p5p5\\\\�\UpU��  p5p5p5_5U5U�    �\\\5\�\U\]  �p5p5p5p5s5}5\}\�\\\\�  u5U5W5\5p5p5�    ��\U\U\�\\\  �UU5_5p5p5p5\\\\�\U\U��  p5p5p5_5U5U�  ����������������w��+�?���������������������������������������� �             ������������� �                  �� � ����:�         0 ���������U�D�x x ^ ^ ^�W�W��E�xEx                   � � _����|j�֯������Ww�~��W���������������������������������_T���l/�/�,�/�,�/�/ /�?0?@? ? ? � �������  ��_�|�z��������������                          ����������UUUEE ��                         ��?_��֪ڪj�j�jU������������j�j��U��������������������������������_<��
�0�0� � � � � � <         P�      @ TO��� ���]���������������������       � 0 0 �  0 � 0 0�<�    �> � ��      = � �Zj=���V    ������������]U\W��U�]�W�E� p p p p �                        = = ������������������W����_����v�ڟj�j�ڧv��_������WT�R�H�B�B�O�C�N�B�J�@u@]P�P�P�P�PUUU�UpU_��_Z�����������V���������������           0 �� � 0   <0�?    �Z�j����կj��کj�j}���U7U� 5��U  � �����������WUWWDEE  E  E  E U _                                      � ���?����_������]j�کu��j�ju�کj��]����_��������������������������������������?� ���_j���z   �?�������������������������������������������S�_���������TS�ӫ���>�C0TL�L������������������Uy� � �                                                                           ? � ��������������������������������������������������������������?   ��UpU\V�j�j�j����������������{�{�{��쩰���ৠ��������� � � � <���^STU�[�]�S�T�?0UL]L_�p��<              ^ ^ xxx�U�_�� �                                                               � ������������������������������������������������������� >        ? �UU=Z=j����֪V�Z�j�������������������������j�ij�j�j�j�j�o��� �?�����n5n[� <     @ T@UT�U_�\| � � �                            _ z��                                                < ������������������������������������*�?�?�?������ � ?                   X�h�x���������Ȳز�����(�8�H�X�h�x���������ȳس�����(�8�H�X�h�x���������ȴش�����(�8�H�X�h�x���������                �������� � �������������������쫬������������������� ? ���:�:�:�:�:�:�:�;�:�:�:�:�:�?������������ � ��������������������������������������
�/�/�
 * ���/�/�������������/�/���*������pUpUpU\U\U\U\}\}\}\}\U\W\]\up�pU�U�U W W��WU���UUUU5U5U5}5}5}5}5U5�5u5]5WUUU� � �?U�����<<<�?�?<��?<<<<�?��?�? �� �?�?<<<�?�?<<<<<?<�<�??<<��?<<<<�?���?<<�?�  ��?<<�?�<�?�? ��? <�?��?�?� � � � � � <<<<<<�?�<??<���??<  ��\U\U|�p5p�pU  �U5U55p55U5pUp�p5p5p5p5�  U5WWWW5\5�    ��pU\U\�\\\  �UU5_5p5p5p5\\\\�\UpU��  p5p5p5_5U5U�    �\\\\\\  �?p5p5p5p5p5p5\\\\�\UpU��  p5p5p5_5U5U�    �\\\5\�\U\]  �p5p5p5p5s5}5\}\�\\\\�  u5U5W5\5p5p5�    ��\U\U\�\\\  �UU5_5p5p5p5\\\\�\U\U��  p5p5p5_5U5U�              ��\U            �U5\U��            U5�            Ե޺����U� �$% �wx��� &'67GHWXghy⼊��()89IJYZijz{����*+:;KL[\kl|}��� 	,-<=MN]^mn~�� �
./>?OP_`op����� 01@AQRabqr������ !23BCSTcdst������"#45DEUVefuv������ �������� �������� �������� ���⽾��� �������� ������
 ������
 ������ �� ���� ���������� �F…���fhi�gjk�GHlm��FIJno��� 01KLpq���������	23MNrs���������
45OPtu��������� !67QRvw��������"#89STxy�������$%:;UVz{�������&'<=WX|}��������()>?YZ~��������*+@A[\�����������,-BC]^�����������./DE_`�����������abc�����de���炊��炍���� � 	
	  � !& � �"#' � �$%( � �  �  � !& �),- �"#' �*./ �$%( �+01 �),-  �*./ � 8234567A � 79:	 �; �< �= �) �s� �$ �s� �$ �t� �V#Ziz� t� �V#$ �(8[j{����U �V# $ �)9\k|���� $ �V#s�*:]l}����dV# �t�+O^m~����e �s� �,P_n����1 �t� �-Q`o�����2 s� �$ .Rap����� �t� �V!/Sbq����$ �
"0Tcr����	u �;<?@CDGHKL���v �=>ABEFIJMN���� �� ������ �� �����' �%3Wfw����7 �&4Xgx����� �65Yhy���� � � � #$'(+,/034 �!"%&)*-.1256 � �	 �#$ �	 �%& �
 �	 �#$ �		 �%& � �	 �#$ �	 �%& �    �  ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`�����������h�Ȁ؀�����(�8�H�X�h�x���������ȁ؁�����(�8�H�X�h�x���������Ȃ؂�����(�8�H�X�h�x���������ȃ؃�����(�8�H�X�h�x���������Ȅ؄�����(�8�H�X�h�x���������ȅ؅�����(�8�H�X���������������� �Ϫ��:�:�:�Ϊë��������������êΫ���������� ��Ϊ��� ��êΪ��ê��������������ΪΪΪΪΪΪ�������������������𪯪����������� : : : : ����������������������:�:�:�ꫪ����             �ê         � � �ê�����þþ����� �κ�ξ�κΪ��          ? ����            3��:�:�:�:����?������>����  �?����������������������������������+�+�+�+�+�+�+�+������������������������z�_�������������  ����������������������������  ����������������DDDD�?�??<<T=DDDD����?  OUU=U=U=�?�? <U=UADDDDUU�� �U�DDDD����? � �WU=U?UOW�_�OOPP�_U�U�U�����  OUOUOUOU?U���� DDDD?O?O � UOU�U�UUOUO?O?O@PDDDDU=U=�? <U=�?�? <U=U=U=U=UADDDD����?  _U���� _UU���� DDDD?_? � �U�?�?@OUOUO?O?O@PDDDDU=U=�<<_==�=�?�?�??U<UA�q��w���3�0�_����������UU  DDDDUUUU��  UU��+���+��
������*�*�*�*�*����]�]�]u]�]u]u]u]�?�����
�
��EEPUUA�T�T�U�U���ժ�����zD{{E}���׫W�W��  5 �?_�U��?5 �?U�Uժ^����U���                      ��z�_UU��      �_�z�굪�� � � �UUUUUUUUUUWU}U�U��|�WU�_<\�_WUWUUUTUQUTUEUP�U���UUUUUUU��U�U���^UUUUUU_Uu_�����                UUUUVUWU^UzU�U�UUUUUUUUUUUUUUUUUUUUUEUEPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUQUTUUUUUUUUUUUUUUUUUUUUUUUUU UPUQUTUUUUUUUUUUQUAQQETPTUUUPUTAUAQTPUAUUUTUUUUUUUUU@@@TTTPQ@PTUUUUUQ@AQDU@UUUUUUUUUUUUUUUQU@UAAUA@UUUUUUUUUU@AUTPU@UQUUE@UQTUQUUUUAUUUTUQUTUEUPUUUU                �W�W�W�W�U�U�U}U��
��*�:�J�Z�j�z���������ʈڈ���
��*�:�J�Z�j�z���������ʉډ���
��*�:�J�Z�j�z���������ʊڊ���
��*�:�J�Z�j�z���������ʋڋ���
��*�:�J�Z�j�z���������ʌڌ���
��*�:�J�Z�j�z���������ʍڍ���
��*�:�J�Z�j�z���������ʎڎ���
��*�:�J�Z�j�z���������ʏڏ���
��*�:�J�Z�j�z���������ʐڐ���
��*�:�J�Z�j�z���������ʑڑ���
��*�:�J�Z�j�z���������ʒڒ���
��*�:�J�Z�j�z���������ʓړ���
��*�:�J�Z�j�z�                  ��??<        ?<�?�    ��?<<<<<<<<<<�?�    <<?<?<?<�<�<�<�?�???<<    ��� � � � � � � � � � � �     � � � � � � � � � � � � � �     <<?<?<?<�<�<�?�????<<    <<<<<<<<<<<<�?�    ����    �?�?    ����    ��??<< ? ��� �   � �     <<<<<<��� � � � � �     �?�?    ��    �?�?    �?�??   ? �� ? < < ?��    <<?<?<?<�<�<�<�?�???<<    ��?<<<<<<<<<<�?�  ����U�U������������eo���_u_U_AO0?��W_U_U_U_U_U_U_U_U_U_U_U_U_U_U_U_U_U_U_U_U_U�V_Y_XX��_Y_Y_Y_�_U_U_U_U_U_U_U_U_�_=__�_U��of������of��of_U�W\ߧ_U��of���������� �f�Z���j�Z�Ue�������UQL�7w�UUUUUUUUUUUUUU�UeUeUeU�UUUUUUUUUUUUUUUUUUUUUUUUUUUU�VUXUXX�VUUUUUUU�ժU�UUUUW�|��k[�\�����Z�Z�Z��������ժ��������ff��������������k���������j�������}��sw]UUUUUUUUUUUUU��UaUaU`��eUeUe��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��V��mW�_��UUUUUUUWU����}UU_�����_�VU��UU����ff��������������������������ժV�j��ʰ*��UUUUUUUUUUUUUUUUUU�ZUeUa`�ZeUaU`UZUUUUTUPDEQT  UTQE@QEQEQTUTUU_UpU_UUUUUUUW�\� <��g����������sf��qup�]�s�]��ff�������������j������������������������U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUAPETEQQETUUUTUPUUUUUUUTUTUUUTUUUTUUUUUUUUUUUUUU�U�U�WU\UW�f����n�[�ۙ�fۛ�\[W�UUU���f��������������������������������������UUUUUUUTUQEUUQUADUUQEUUQUTUUUU��VVV��UUUUUUUU��VVV ��UUUUUUUUUUUUUUUU��UU��u]�[�VUU}���p����  �|�\U�w�VU��VU�������������j����������ꪪ����U�UUTUTTUUEPQEUUAUUEQPUUTTTUUU��VVV��UUUUUUUUUUVUVUVUUUUUUUUUUUU�U�U�UUU���U�U�W���qn���n���>�=���mŭŭ�������f�������������������������������WUUU��VVV��UVUVUV��VUVV��UUUUUUUUVUVUV@EUEDEUU@QPQQUTQUQQU��j��uW�j�ZVF2SL0�PQ\U\U�W}_]]VU��Z��ff��������������������������������������U�UU��VVV ��UVV V�UVUVUVUUUUUUUUUUUUUUUUUUUTUTUT�U5�@UUUUUUPUTUU�TfQfWfUfU�UUUUWUWU\U\U��lf������, ������ WU\U��ff������������������n�������n�����������UUUUUUVUVUVUUUUUUUUUUUUUUUU�UuUuU�U�U�U�U�U�U���j����UUUUUU�U5U�UUUU��k��յֵ���U�UUUU��ff������ ������ꪪ  }U�U��ff������������*����.���������n����������U�UUUUUUUUUUUUUUU�UU��U_������j�Z�Z�Z�Z�j���������=7�7sU\U�����U�U5�WW�   �Ze�Z����f��W���U�U��_�����  UUUU��ff����������������j��������ꯪ���UUUU�U5U� 5       =��#C-49�9��@�@�C�C��?��U0 ��|�0��035�<� � �      y �An��骾����j�z��U�U��������_UUUUUU��ff�����������j���������k����������:���5            ��      �
      
�  # # � ? � � ����0pp p\�\ W \uN�z��٬k�k�n����Wq���ƪƪZ������������UUUUUUUU��ff������������*�?��Ʀʕ*W�\:�� S C ��               
� � p p
\ \ W W�U�U�UpUpU\U\UWUWUUUUUUUU�U�U�UUUUUUUUUUUUUUWUW�W�W�]j�P�T�T]�mf����������ff��iU�UiUU�UU��ff��������������
��Ws�ݺ:�:���:_:p5���UpUpU\U\UWUWUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UURUR��PUTUTU��UUUUUUUUUUUU�j@�T�T��j�U�U�Uj�ff����������ff��UUUUZUiUUU��ff�������?��N�N�N�L���]�����L�L�N�N�N�O�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�N�M�M�M�N�N�N�N�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�N�N�N�N�N�O�N�N�z���������U���f������          ��  <<<?�������<<<�?�?<��?<�?�   <??�?�?�<�<�<�<��?<<<<�?��?�? �?�? �?�?��?<  <�?�<?<�<�<�?�??<� � � � � � � � <<<�?�?<<<�?�?�������,�<�L�\�l�|���������̖ܖ�����,�<�L�\�l�|���������̗ܗ�����,�<�L�\�l�|���������̘ܘ�����,�<�L�\�l�|���������̙ܙ�����,�<�L�\�l�|���������̚ܚ�����,�<�L�\�l�|���������̛ܛ�����,�<�L�\�l�|���������̜ܜ�����,�<�L�\�l�|���������̝ܝ�����,�<�L�\�l�|���������̞ܞ�����,�<�L�\�l�|���������̟ܟ�����,�<�L�\�l�|���������̠ܠ�����,�<�L�\�l�|���������̡ܡ�����,�<�L�\�l�|�����UUUUUUUUUUUUUUUUUU�_�}_U_U_U_U_U_U_U_U}��_UUUU�_�_}_}_}_}_}_}_}_}_}_}��_UUUU_}_}}}}�}�}�}��___}_}UUUU�_�_�U�U�U�U�U�U�U�U�U�U�U�UUUUU�U�U�U�U�U�U�U�U�U�U�U�U�U�UUUUU_}_}}}}�}�}��____}_}UUUU_}_}_}_}_}_}_}_}_}_}_}_}��_UUUU����_U_U_U_U��_U_U_U_U����UUUU�W�__}_}UU_�_�W�U�UUU�U�UUUUU_}_}_}_}_}}_�_�W�U�U�U�U�U�UUUUU��_U_U_U_U�_�__U_U_U_U��UUUU��U_U_UU�W�_UU}U}U�_�WUUUU_}_}}}}�}�}�}��___}_}UUUU�_�_}_}_}_}_}_}_}_}_}_}��_UU����U_U_UODOD    __UT U_    ���W�U�u�U�U�U�� �W?\{��ololo�o����q�ů���Z�Z�Z�j�j�j�j��������ϻϮ��_�o�o��ſ�V�Z�j������������UUUUUUDDDD        UAT @ @UU     �� �\W5�7�5W5W��  uU�u��󪱫�j���jū�jū�j��󪳫󪌫̪��1�Ÿ��Ÿ�[k������V�V�Z�k�o��Ŭűű��j��������UUUUUUDDDD           U       �?��_5u�������������? @��{�����;/����Y�V�YVYf�j����f��쮱����WkZ�Z�Z�Z�j�j�j�j�Z�[�[�\���������UUUUUUDDDD                      0@ @�   0 �         PCP    SP  2 � [nk1o1�1�1�1�1���ż����Z�[�n�k�lò̲�����+Z,ZlZlZ�Z�j�j�k���������UUUUUUDDDD                  PUUQ  U T               U U U   TT                  @   @           1 � ŀ� ƀc[�[qlq�q����������������UUUUUUDDDD                    P  U                         @                     @    P @          � XV	XV	U%V	U%U�U%U�UUUUff��ff������������UUUUUUDDDD     ��|��?<< ��UpUpU�U\�\U\�����p��W\��             @  @           @ @   TUU  QUUQU@@          �`	X%`	X%V�X%V�UUUUUUff��ff������������UUUUUUDDDD                7 5 �@uS�7M U            @TUT  UU           @   EEUU  TEUU D           �`	X%`	X%V�XeV�UUU�UUff��ff������������UUUUUUDDDD                      PTUT    T U                 @         �       @ ��@���< � | � 
�%`��%`�XUVUXUVUUUUUUUVUUUUUff��ff������������UUUUU��4  ��������� 0 � �   PUU@    UU                           5 �w��W_��UUUw���w7U5W�? �?_��?       	�`	�%`�X%`�XUVUUff��f�>�C��������UUUU��      ??� �      ��   UT U P T U                                       @@               
 % � %���U0UNUMUS���S�T�;��������UUUU��      <<?<�<�<�<�<�?��      �   0 �             �0  �<\ �0�W W � W W �� �U � � L L SS���0�0�0�0�L�L�L�L�L��3�3>3:L>L;�N�S͔Τ>�C�P��ꤺ����������UUUU��      <�?�??<<�<�<<      ��  3 <    �   � �  ? ��W�}���u�U�_�u�U����T ]U{�ꬪ��S�S����>�:�?�N�O�N�Sꓺ�ꓺ��;�>�O�N�S�S������;��C�P���������UUUU�U  p ��? < < < ?     � � 0 �     ��0s�p���03����0;쫪��������U�u5u5�7�TUUU�_�t�:�>�:�>�:e>�:e;�>e;��dӔ�TS��N�N�O�N�O�N���>�O�N�O�S�������������UUUUUUDDDD        PATUP  U               ���WW�����U�pUp��  UUUU�|��ﺻ��������>�;�>�?�3�4�4�L9M6M9MMNONPN�N�O�N�O�Ӻ3�4;5�������U�U�U��D��D�� � � � � � �P�U���� � �U� � � � ����� ��� ����u�u�]�]�]��������U�W�~�������������������������������������:�>�:�>�:�M��������������UUUUUUUUUUUU�W�W_}_}}_�_�W�W�W�W�W�_}__}_}��_}�_�_}��__U_U_U_}���}�}�}�}�_�_}_}_}_}��_��_U�_�__U���_�_}_U_U_}��__}}�}�}��__}�U�U�U�U�U�U�U�U_}_}_}��_}_}_}���W�W�W�W�W�W>�N�^�n�~���������Τޤ�����.�>�N�^�n�~���������Υޥ�����.�>�N�^�n�~���������Φަ�����.�>�N�^�n�~���������Χާ�����.�>�N�^�n�~���������Ψި�����.�>�N�^�n�~���������Ωީ�����.�>�N�^�n�~���������Ϊު�����.�>�N�^�n�~���������Ϋޫ�����.�>�N�^�n�~���������άެ�����.�>�N�^�n�~���������έޭ�����.�>�N�^�n�~���������ήޮ�����.�>�N�^�n�~���������ίޯ�����.�>�N�^�n�~���������UUUUUUUUUUUUUUUUUU�_�}_U_U_U_U_U_U_U_U}��_UUUU�_�_}_}_}_}_}_}_}_}_}_}��_UUUU_}_}}}}�}�}�}��___}_}UUUU�_�_�U�U�U�U�U�U�U�U�U�U�U�UUUUU�U�U�U�U�U�U�U�U�U�U�U�U�U�UUUUU_}_}}}}�}�}��____}_}UUUU_}_}_}_}_}_}_}_}_}_}_}_}��_UUUU����_U_U_U_U��_U_U_U_U����UUUU�W�__}_}UU_�_�W�U�UUU�U�UUUUU_}_}_}_}_}}_�_�W�U�U�U�U�U�UUUUU��_U_U_U_U�_�__U_U_U_U��UUUU��U_U_UU�W�_UU}U}U�_�WUUUU_}_}}}}�}�}�}��___}_}UUUU�_�_}_}_}_}_}_}_}_}_}_}��_UU����?   �0���            PO OP    OP   U_         @O     �?�@U_�_���_U_�_�_7_M_S�T�T?UU�U��_�U��������     0�|W�U��pupu\u\U\U\�\�\�p�p��� W |�P  U    � � � � ��@�@��� � � � � � �      @@        � @� = � S�TUSUTUUUUUUUUUU�U�����UuU]U��������    �W�UUUUUU_�u]u]u]UUUUU�������
����UUW��     �|W�U�UkV�UkV�UkV�Uk֫�k֫�k֫U�U�V�U�V�U���կ?�      �?0@�U�U�U�U�U=U�� = �?�uUu�_]U]U]Uu��������     0 �50�0��]�]]UU_zzz^� 5     � ��o��UUUU}U�U��50�3<�@�� � � pp=��_YDjQZD��        ��|��������� �   �  S S�T��0�0UOUq���W_\q}���������           @ @    @ P     ���*�If�EVUEU}U�U�U�UpUpU�UW_s�p�p>p5\�WUUUU���?��Z̚0�0�����Uͪ:�ꪪ�����? @UUUUU_�_�_�W}UUUU���_�UUUUU��������               P T           @ P         @q t1T5 5 5 5 5 5 5 5P��� � ?  � \{=���l갪ê�:�ꬪ���0�?��0UOU]U�U�UU5U5U5U5U�U5U5UMUM��������               P T          T  T           TP         U @             ��W|UW�����]�u�ץ^�y�f�����;�     �� PUUUUUUUU���� ��_�PUUUUUUUUU��������       � W | ��pu�w ��\�� � � �@q� �         P@       PP             ��UU����������������z���� � � � � � � ��� �UUUUUUUU���� �_�UUUUUUUUU��������        5 7 � � ���P� UCV?��]W �ppWp\�\�pq��U@W\ � p p \ \ � ��u�u���wV]��������U�z��_��k���
h�B�?����j���j�����������������C�T�T1U�u����������       ��Wp�p�����p�p���� ��z�^s]�UUU�_���������Z\ku����_��u�WW�    �W��V���������������uv���]^�z�y�y�xk���?8   ��UU������_�UU_}_}_}_}UUUU��������      � U?�ժj�����������������וUUUjU��U����z�_�U_UU�w�]z����upup]\]\WU���C�]jwjצ՝՝6�6�6�5��jZ� =           �V=�֪ګ?� � U]�W���������          ? �}=v�v�ڵڭo������{�^U~VY�շ��U�U�U5���  tt tt�w�wU�U��� � 5 u P @           � W W �         � 0 L S���up]p]\U\U\�תת�Z�jU���������                 @ P       C@      ��         PUU_��?    P       @U TU@   P �U�UU�U ��U�[C�TUUUUUWU]}]�����UUU��z�z�^�W��������            P@        P U           �p�\y\n�kW�W�W�]�]���y�yU啕��?          U@          P@        �U�WU�W� � UUUU5U5U5U�U�U�U�U�U�U�U���������            @P       @P        �\��� :��W}�U��_�W��� V^�5P T @  @U              @    @            ��\U��   � �P0����SU�UW_U�������� � � � � � � ������ � � � � � � � � � � � �S����S� � � � � � � � � � �� � � � � � � � � �T��T� � ���@� � � � � ���U���7���U�U���]�]�U�U���W����UUUUUUUUUUUU�W�W_}_}}�_�W�W�W�W�W�_}__}_}��_}�_�_}��__U_U_U_}���}�}�}�}�_�_}_}_}_}��_��_U�_�__U���_�_}_U_U_}��__}}}�}�___}�U�U�U�U�U�U�U�U_}_}_}��_}_}_}���W�W�W�W�W�W�������ű˲ѳ��K�GX�RQVX�SUNX�TPOX�K�X� 	X�KRQX�
X�KSUX�KTPX�K�X�K�GX�RQVX�SUN�TPOHKGWIKHKGWIKHKGABC?KRQVMJKRQVMJ34679;=>ESUNLFKSUNLFK5U8:<D@Y12�"!&(*,.02K�$# %')+-/K� �'1;EOYcmw������ �(2<FPZdnx������ �)3=GQ[eoy������ � *4>HR\fpz������ �!+5?IS]gq{������ �",6@JT^hr|������ �#-7AKU_is}������ �$.8BLV`jt~������ �%/9CMWaku������ �&0:DNXblv������� �	 	 �
  � � � � ����� ���� �����ž� � �'1;EOYcmw������ �(2<FPZdnx������ �)3=GQ[eoy������ � *4>HR\fpz������ �!+5?IS]gq{������ �",6@JT^hr|������ �#-7AKU_is}������ �$.8BLV`jt~������ �%/9CMWaku������ �&0:DNXblv������� �	 	 �
  � � � � ����� ���� �����ž� � �'1;EOYcmw������ �(2<FPZdnx������ �)3=GQ[eoy������ � *4>HR\fpz������ �!+5?IS]gq{������ �",6@JT^hr|������ �#-7AKU_is}������ �$.8BLV`jt~������ �%/9CMWaku������ �&0:DNXblv������� �	 	 �
  � � � � ����� ���� �����ž� �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`Ҁ�����,�>�P�b�t���������΁�����(�:�L�^�p�����������<�~����D���Ȅ
�L���0���Đ6���ڑ,�~�В"�t�Ɠ�j����`����V�������0�B�T�f�x���������җ�� �>�\�z�����Ԙ��R���֙h������`�
�D���0�T��x�
���.���R���<<<�?�?<����?<�?���?<  <�?���?<<<<�?��?�? �� �?�?�?�? ��   �?�? ��?<�?�<<<�?�?<<<�?�?�����?�?�?�?������ <�?�? ? ��?<      �?�?<??�?�<�<�<�<�<<<?<�<�??<<��?�?<<<�?���?<<�?�  ��?<<<�?�<��?<<�?�<�?�? ��? <�?���� � � � � � <<<<<<�?�<<<<<<���<�<�<�<�<�???<<??<���??<<??<��� � � �?�? ��� �?�?                    ���pUU\UU5\�_5\p5\p5\p5\p5\p5\p5\�_5\UU5pUU���         �  \5  W5  W5  W5  5  p5  p5  p5  p5  p5  p5  p5  �         ��? pU�\UU\�W\W���  p5  \  W ��  ���pUU5pUU5���        ���pUU\UU5\�5�p5 �5 WU WU �5�p5\�5\UU5pUU���          �  �W |U WU�UUp�Wp5W\W\�W\UU5\UU5��W  W  �         ���\UU\UU\��\  \��\UU\UU5��5  p5��5\UU5\UU���        ���pUU\UU\��\  \��\UU\UU5\�5\p5\�5\UU5pUU���        ���\UU\UU5\�5\p5�\  \  W  W ��  ��  p5  p5  �         ���pUU\UU5\�5\p5\�5pUUpUU\�5\p5\�5\UU5pUU���        ���pUU\UU5\�5\p5\�5\UU5pUU5��5  p5��5\UU5\UU���    (      ���             �      ��*          h)   ���VU�    ���  V�      ��*    pUU �AA   �*  (     ��� �!H  �� � �
�
 p  `!H	     �U�
  �  `!H	     `U	��
��W `AA	���*  `U	 �* pUU `UU	VUU�  XU% � pU `�j	���*� XU% �* \<T5 `V�	 `	 � � 
�\<T5 `UU	 �* � ����  \< 5 `UU	�V�� ���    \<�4 `UU	`UU	  ���    W � `UU	XUU%� �    W������XUU%"VT�    W]UU\UU5XUU%� ���?   W]UU����UU�����ꨨ W]UU�j�
Vj骪:���?   W]UUX�W%VUժ�:V��    W]UU�~�*VUժ�:V�� �*�uQQ W� VUժ�:V�� *�r�uL�UUX�֦�:V��  "\UwLpUU���U�:֪�# "\UwLpAA���]�:֪�#  |�L\05���]�:���.�
�u�Q� \05�W�]���UU.  \U�U� \05\]妩���.  \U�U� \05G�ꪪ:�Z����^U�U� \AA53sժ�:���  �� �? \UU533���:���    W5 \UU5G4 ���   �0 \ \�5�7 �� 
  �����?\�_5w= ���  \UWUU�\�W5w7���?�D  \U����\UU5wݰ����  ��   ���?��������?  WU   WUU�W5    �*��  ��   �����?    ����        (      ���             �      ��*          h)   ���VU�    ���  V�      ��*    pUU �UU   �*  (     ��� �EQ  �� � �
�
 p  `!H	     �U�
  �  `!H	     `U	��
��W `!H	���*  `U	 �* pUU `EQ	VUU�  XU% � pAU `UU	����  XU% �* \<U5 `UU	 `	�  � 
�\<@5 `��	 �*�  ����  \<<5 `�Z	�V��  ���    \<<5 `UU	`UU	  ���    WAA� `UU	XUU%* �    W������XUU�� VT�    W]UU\UU5Xii%* ���?   W]UU���Vii�����ꨨ W]UU�j�
Vi骪:���?   W]UUX�W%VUժ�:V��   �]UU�~�*VUժ�:V�� �*p�uQQ W� VUժ�:V�� *�^UwL�UUX�֦�:V��  "\UwLpUU���U�:֪�# "|�wLpAA���U�:֪�# "�uL\05�U�ߟ:���.  \U�Q� \05�W�U���UU.�
\U�U� \05\]妩���.  \U�U� \05W�ꪪ:�Z�������U� \AA5Gtժ�:���    �? \UU533���:���  �0 W5 \UU5G4 ���   �0 \ \�5�7 ���*  �����?\�_5w� ����  \UWUU�\UU5wW���?�D  \U����\UU5w������  ��   ���?�7������?  WU   WUU�W5    �*��  ��   �����?    ����        (      ���             �      ��*          h)   ���VU�    ���  V�      ��*    pUU �UU   �*  (     ��� �EQ  �� � �
�
 p  `!H	     �U�
  �  `!H	     `U	��
��W `!H	���*  `U	 �* pUU `EQ	VUU�  XU% � pAA `UU	���� XU% �* \<<5 `UU	 `	  � 
�\<<5 `��	 �*   ��  \<<5 `�Z	�V�" ���    \<<5 `UU	`UU	   �    WAA� `UU	XUU�
 �    W������XUU%  VU� � W]UU\UU5Xii�
 ���?� W]UU���Vii������ W]UU�j�
Vi骪:���?  �]UUX�W%VUժ�:V��   p�]QQ�~�*VUժ�:V�� �*\UwL W� VUժ�:V�� *�^UwL�UUXU�*�:V��  "|�wLpUU����0:֪�#  �uwLpAA�_��0:֪�#  \UQQ\  5�U��0:���.�
\U�U� \  5�W�*���u].  \U�U� \<<5\]媪��u].  ���U� \  5W�ꪯ:���������� \AA5Gt��:���  �0 w7 \UU533��:���  �0 �5 \UU5G4 ���   �0 \ \�5W5 ����*  �����?\�_5�� ����  \UWUU�\UU5w����?�D  \U����\UU5w7�����  ��   ���?w=������?  WU   WUU��7    �*��  ��   �����?    ����                   0   �     ?� 0 � ;  ��� ����  ��>�3����3�������  ����������  ������������������������������������������  ����������������������������������������  ��������������������  ���������� �������������������������ꪪ����:��:����:;�:� �������  0    <�������������0 ��<<<<�  �?�?<<<<�? 0 <<<<<<�<<< � �?<<<<�?<< � ��?�?<?�? 00 <<��<<� ���������������������� �  �? ������������:���:���:���:���:쪪;���:���:���:������:���?��������� �  �? ������������:캮;캮;���:���:���:���:���:���:������:���?��������� �  �? ������������:���:���:���:���:���:���:���:���:������:���?��������� �  �? ������������:���:���:���:���:���:���:���;���:������:���?��������� �  �? ������������:쪪;���:���:���:��:��:��:���:������:���?��������� �  �? ���������쪪;���:���:���:���:���:���:���:���:������:���?@UU���@UU �  UU P����������_}��}���������_��_���@��TUU�������@UU���@UU �  UU P����������_}��}�������UU�UU�W���@��TUU�������@UU���@UU �  UU P�����t��������������W���A������@��TUU�������@UU���@UU �  UU P�����t��������������W���������@��TUU�������@UU���@UU �  UU P�����������w}�_}�������_��W��_����@��TUU�������@UU���@UU �  UU P�����������w}�W}���������������@��TUU����������pUUpUUpUU\UU5\}U5\}U5\}U5\}�5\UU5\UU5\UU5pUUp]upu]��W�UU���?WUU��������pUUpUUpUU\UU5\}}5\}}5\}}5\}}5\UU5\UU5\UU5pUUp�p�_��W�UU���?WUU��������pUUpUUpUU\UU5\]u5\}}5\}}5\}}5\UU5\UU5\UU5p�p]�pU��UU�UU���?WUU��������pUUpUUpUU\UU5\UU5\UU5\UU5\�5\UU5\UU5\UU5p�Wp�_p�_��W�UU���?WUU��������pUUpUUpUU\UU5\]u5\}}5\}}5\}}5\UU5\UU5\UU5p�_p�p}}�UU�UU���?WUU��������pUUpUUpUU\UU5\UU5\UU5\UU5\�5\UU5\UU5\UU5p�_p�p��UU�UU���?WUU�����          ��      ���?��    ��?<<<<�?�<?<�<�<�?�??<��?<<�?�  ��� � � � ���?�?��������?<  <�?�<??�?�<�<�<�<�<����������?�� < �?�?<<<�����<<<<<<�?���?<<<<<<<<<<�?�����������������? ��� � < <   �?�?��?< < < <�� < < <<�?� ���<<<�?�?  ��    ��? < < <<�?���?<   ��?<<<<�?���?<   ���� � � < < ��?<<<<��<<<<�?���?<<<<�?�? < < < <�?�������:���:��� �: ������������:쪪;���:���:���:���?�����������
���/���/���
 � ���
���/~����׿~�����_��_�/���
���*�����������pUUpUU\UU5\}}5\}}5\}}5�UU7�W�7\}}5p�W�UU W� ���?WUU�����  �  <0�<��;����;�<0p<��\5;3��W��0��UU;0�zUU����z^y�z^y�zy^��y^���W���� ?��u]�����W<0��ZU ������z�W<�޵^3ܼ��W<�������������������� ����   �:   ���  |UU=  ��Z�  ���� ����Z����Z����Z����Z����Z����Z����Z����Z����[���Z����Z����U��������UU5�����?��������_����U ����   �'   ���  ��) ���������	�_��'�����'����W��U�WU����WW��������W��՟�W�_�'�_UU�'��UU�	��_�_ ���� �����*�������������UU �UUU�UUU�U_��U_�pU_�UpU_�UpU_�UpUUUUpUUUUpUUUUp}UU_p�U�UpUWuUpU]]U�U�W�UUU WUU�  \UU0  �U   _�  �����\UUU0�����?<�<  <�?<  <<<  �<<  �<<  �<<  ��?�?  ���  �<� <<�?��<� <<�?�?�<� ?<?< <�<� ?<?< <�<� ?<?< <�<� �<�< <�<� �<�<��?�<� �<�<���<� �?�? ��<� ?? ��?� ?? �?� ?? ??� <<�?<<� <<�?<� �?� �?� ? �  �  � ? � �� ��  ?�  <�  <�  ?� �� �<�<<�?<<<<<<<<<<<<<�<<�<<� <<� <<� <<� <<� �?�?� ����<�?�???<<�? <�? <�< <�< <�< <�< <�< <�< <�<<<�<�?�?�<���< �  W �U wU�?wU]�w]]�w]�?w�� wu� w�? wu� wu� w�? �u5 75 � �����? �� �������w?��������3���?0 ���?  ��������?����  ��?�����03��  p��  p�_  ��x�-�x�C-�p�B��@�����������������?�����? �� �������w?��������3���?0 ���? ���������? ��� ���?0����00��  p��  p�_  ��x -�x�@-�p@��@�����������������?�����?�W����w����������������<���������?����?�����������������������������?����00���������?���  <�������?��3� ������?�����?�W����w����������������<���������?����?��������������������������00����?������� ����������0�0���?������3��?������?�����?�?�����?�������_�_�����}��������������??�����?���������� 3� ���3���<<���3���0����� 0��0�<  <��?��+�3��?0������?�����?�?�����?�������_�_�����}��������������??�����?���������� 0 ���3���<<���3���0�������0��0�<�<�<�?<���3��?0������?�����?���/����������������?<��?��?  ��?  ��<���3��0�3 2����:�#�� �,�8�� � ����*�� �� 0��� �� ?�� �������?�����?���/����������������?<��?��?  ��?���<����3 2�3<�0����:�#�
#�,��� � ����*�� ������?� �� ?�� �������?�����?������_?������������?���������<���� 0��Ï
����/���L?0���<�1���<�1��� ��,  ��0����� ���@��������_���S�������?�����?������_?������������?���������<���� 0��Ï
����/  ���  0���?�0��<0�  �� ��,���0���������L��������W���S�������?���L����`���̦�"�F������3�M�o�����ߩ?�����_�����߬?�����_�����?�O�_�*��}�    ������������ �:  �  �� ���������������������:���:���:���:���:���:���:������:���?                ������������ �:  �  �� ���������������:���:���:���:���:���:������:���?������������ �/  �* ���������/8�?,��Ͽ�������������?������/�?�/������*������������        ������������ �/  �* ���������/���/�?���Ͽ���������/��/�����說+�������� �� �UU�UUpUUpUUp�Wp�Wp�Wp�Wp�WpUUpUUpUUp�WpUU�UU�UU W�  �?  \5 ���\UU5���?         �� �UU�UUpUUpUUp�Wp�Wp�Wp�WpUUpUUpU]p�W�UU�UU W�  �?  \5 ���\UU5���?��6�ի���:��?  p�  s��?\�U�\�U�\��?\}5 \W5 \� \W5 \W5 \� |W5 �W5  � �l6�?��p��9l6�9��9�?�?g������4l2�9�?��gƛ�gƛ�g��?g��� �� ����� �  �?  ��  g�  ��  g�  �� ��I�f&���f&����ff��� �� �����������?�?�?�?���?�? � � � � � �; �;������������ �; �; � ������� �  �?  �?  �  �?  �� ��������������������������� ��  �?  � ��������:l9l9l9l9l9l9���l9�?�?��[�[�[�[�[�[�[�[�[�l9l9�.�?W��� �� ����V��V��V��V��V��V��V��V��V��V��V� [�  [�  l9  �.  �� �V�������
XUU%XUU%���
 `	  �* �V�`UU	XUU%XUU%XeU%Xei%XeU%XeU%XUU%XUU%XUU%�Z�&h�Z)XUU%XUU%���*VUU�����        ���
XUU%XUU%���
 `	  �* �V�`UU	XeY%XeY%XeY%XeY%XUU%XUU%XUU%�Z�&h�j*hff&hff&���*VUU�����    ���\UU5��� p  �  |=  W� �UU�UUpu]pu]pu]pu]pUU���p]wp]up�_pUUpUU���?WUU�����        ���\UU��� p  �  |=  W� �UU�UUpUUpu]pu]pUUpUU���p]wp]wp]up�_���?WUU��������*VUU�VUU����*`UU
`U�	`Yj	`�e	`�e	`�e	`�Z	`eU	`YU	�VU�UU��Z�ie�UU V�  V�  X% ���*  �����    ���*VUU�VUU����*`UU
`U�	`Yj	`�e	`�e	`�e	`�Z	`eU	`YU	�VU��Z��j��Z ��  V�  X% ���*VUU�����                 �  �� ������������:���:���:���:���?���լ�~լ��լ��?���:�ww;�ww;���?��������         �  �� ������������:���:���:���;��>���:��_;���:���:���:���;���:���:���:���?�������������������� �:  �:  ��  �� ������������������������:���:���:������������?�������������������� �:  �:  ��  �� ������������������������:��:��:����������?�����������?\UU5���? p  \5  W� �UUpUU\UU5�_�7ww��wu]�ww���]u�\UU5\�5p��p���W�UU W� ���?WUU��������?\UU5���? p  \5  W� �UUpUU\UU5�_�7wu]�ww��ww���_��\UU5��7p��p}}��W�UU W� ���?WUU��������*VUU�VUU����* `	  �* �V�`UU	`UU	`Z�	`eY	XUU%�j�&���*���
�j�
�Z�`UU	`ii	`��	�UU���*VUU�����    ���*VUU�VUU����* d  �* �V�`UU	`Ze	`eY	XUU%�j�&���*���
�j�
�Z�`�V	`�Z	`ii	�UU���*VUU��������`UU	��� `	  �* �V�`UU	`eY	XeY%XUU%Xii%X��%XV�%XUU%XUU%XUU%XUU%XUU%���*VUU�����                        ���`UU	��� `	  �* �V�`UU	`UU	XUU%XeY%XeY%XeY%XUU%�UU&X��%XUU%XUU%XUU%���*VUU�������? pU� ��?  \  W  W �u7 �u7 �U5 ��7 �]= ��? ��� �u� �U5 �� ��? pU� ��?  \  W  W �U5 �}? �U5 ��� ��� ��? �]= ��7 �U5 ��?     �����?��  ��?���������?�    �         �    ��    �    �    �0   �W�    pUU   \_}   �u�   w�U7   w}_7  �u}_�  �u}_�  �u�U�  �����  p�_�U \�U�V \uuW[ WUUUU5 W���_5 W���_5 \���W �ի��  _�_=   �U�    _=     �    � �      ��    �0    �<    �    �W�    pUU   \UU   \UU   W_}5   �u�5  �u�U�  �uUU�  �u}_�  �u}_�  pu}_W p���U \�_�U W�U�V5 WyuW[5 WUUUU5 \U�WU �U�_�  _�W=   �U�    _=     �    � �      ��    �0    �<    �    �W�    pUU   \UU   \UU   W_}5   �u�5  �u�U�  �uUU�  �����  �u}_�  pu}_W p���U \�_�U W�U�V5 WyuW[5 WUUUU5 \U�WU �U�_�  _�W=   �U�    _=     �      �         �    ��    �    �    �0   �W�    pUU   \UU   \   ���5   wUU7  �uUU�  �u�U�  �u�U�  �����  p�^�U \�U�V \uuW[ WUUUU5 W���_5 W���_5 \���W �ի��  _�_=   �U�    _=     �   �  W �U wU�?wU]�w]]�w]�?w�� wu� w�? wu� wu� w�? �u5 75 � ����� �(�1�=�J�U�b�i�w�����������
T  <P@>A?B0C>DF04C>DF0LC>DFP H(	H8 HP 	H`<<`x 
H�	<	<
H( 
H8<<HPH` Hx	H� ������������������������������������������������������� � � �1���Q�@�@�@�� � � �p�p�p�@�@�@���� � �p�p�p�p�@�@������d�p�p�p�p�p�b������D�D�p�p�p�p�"�"����D�D�D�p�p�p�"�"�"��D�D�D�T���2�"�"�"��������������������������������������������������Ĵȵ̶          
                                   0 2 4        = ? A C E G I K M O  R T V X Z \ ^ ` b    g i k m o q s u �    | ~ � � � � �      � � � � � � � �    � � � � � � � � �  � � � � � � � � � �        � � �                � �                  �                   �                  � �                � � �        O b u � � � � � � �  M ` s � � � � � �    K ^ q � � � � �      I \ o � � � �      4 G Z m � � � �     2 E X k ~ � � �  
  0 C V i | � � �        A T g                ? R                  =                   �                  � �                � � �        = R g | � � � � � �  ? T i ~ � � � � �    A V k � � � � �      C X m � � � �      0 E Z o � � � �     2 G \ q � � � �  
  4 I ^ s � � � �        K ` u                M b                  O         ���������� ������������������ � ���������������� � � �������� � � �2� � �7� � � �� � ����� � � ���� � ������ ������,������6������ ������� ���� � ������ � �� � � �5� � �4� � � �������� � � ���������������� � ������������������ ���������
024CEGIǲŝ�È���������|�������������=R?gTA|iVCObMu`K�s^I��������������&�*F�V�f�v���������ƹֹ������������ ���������� � ���
������� ����
���� ���  
��� 
��������� ���
������� � ���������� �������� 
���  
��� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�������l �'������ �����a ���` 1� �� ��`�	)�`��!�T�"�\�#�$ �` 8�� ��.���q��- ��恥�)���	 ��怩 �-` ��
�? "���`�a�
���4�5`�	)�惥���� �������!��"�`�# m�`%&''%&&' �� ��������`� �4�4�5`��
���������l ������@��������A�J�h������������v������� �`� ���p����a�P���p����b�~���p���@� ��
� �!�"�(� �6���� ?� C��6�6���怩 �P�Q������` 
 !"( �� �� �� ��`�)�=�
�E� � E�)�
Ƃ����
悥���� ���������@� � � ?� C�`h��)�M��E���� Eू�t��8���
ƅ����
慥���� �����������@�(�(� ?� C�`���
�Q�Q��
�Q�Q��� �Q�����x���@�
�
� ?� C�`���
�P�P��
�P�P��� �P��������@��� ?� C�`8h@hPPHH
(�	)�%�Qi � EॄI���Q�
e��`�@�  ?� C�`�= ?�P
ePeQ� 
e �� �<ÙS �V ����񦅽9Åg� �8� �]�^�_�`�4�5`	      ��
��qÅ�rÅl u��å8i�(� �'�(�
�� �(��'�'i�!�(�"�x�# mߥ(i�!�8�"�x�# mߩ���-�. �� �V�S���� ���`���� �Y�Z�[�4�5`�������������������������������
��ą�ąl �?ę� Ʃ ����@� �x���S���%�@ ?� C� ���` F� ~�`�	)�%� � E�恥���� ����rč@�@�  ?� C�`%&%&%&%&%'('���� \ũ�-�.�� �������� ��>Ņ!�GŅ"�PŅ# m����	�� ��Q���Z�!�0�"�YŅ# m������ ��Q���E�!�H�"�YŅ# m�L�����ߠ �� �/�0�1�^ �d��d�^ �/�^ �
�	�
�^ �0���1 p������ ���`JKLSTUIIIppp1I0H0H4L��!��"�x�#�X�$ �`� ��/iI�!��Ņ"���Ņ# m������`X`h0H F� ��`���M \Ţ ���Ņ!��Ņ"��Ņ# m������f��Ņ!�8�"�(�# mߩ]�!�\��!�`�"�D�# m� ���`V[\8HDDWXY Fĥ��� �^�_�`�\i�4�5`��
��,ƅ�-ƅl 0�QƩ ���)�@�@� ����x�� ?� C��`�0))�$��E��I��� � Eং��ƍ��@�  ?� C�`����`��4�5`T������������������������������������������������������������������������������������
���ƅ��ƅl �Ɠ� '� �� g� � �ߥ]�R� �����������ą��ͩ����������`� �� ����P)��Q��ǅ���ǅ�Ը� ��Ǚ���Ǚ���Ǚ@�@� �� ?�Lp� C���������Ы`  
PHX@P`8HXh�����x�xph ( (08&&&&nbnVbnJVbnnbnVbnJVbn� ���� ����S������`�
�!�ȅ"��˪�Ը�� %"� ��!��`���)�!�h�"���# mߥ8i�(� �'�(�
�� �(��'�'i�!�p�"���# mߥ(i�!���"���# m�`� ���������`����#�� )@�� E����3��` � 3ʦR�S
���ȅ��ȅl �ȴ�rэԥ�
���ȅ��ȅl ��z� �D� �� 8�`�	)�)�` � E�� �  j�` �� ɦ�@�  C�`�R���e��` � _� ��`�	)?�)�` �ɦR�S����WɅ!��"�# m�` �ɦR�S����[Ʌ!��"�# m�`*,,.+--/�	)?�)�` ʦR�T�����Ʌ!��"��# m�` ʦR�T�����Ʌ!��"��# m�`20243135�	)?�)�` ʦR�U�����Ʌ!�(�"��# m�` ʦR�U�����Ʌ!�(�"��# m�`8869::7;��!�"��#� �$ �`��!��"�'�#� �$ �`�(�!��"�7�#� �$ �`�	)����`��!��"�1�#�%�$ �`�=�!�R�gʅ"��# m�`,��� ���D� )@�=����!i�#���"i�$�@� ���/i����0i� M� ��� C����$��`��� ���F� )@�?����!i�#���"i�$���/i����0i� M� ��� E��@� �����`� �� )@� C������ @�`�)��)
��) �%`��E ��悥��
�� ��`��E ��Ƃ�	��`��E ɦ� ���� �˥��.����� �� � E����掦�䄐� �� � �� � j��` �ȩ(�!�p�"��# m� �ߩ���E` 
� ���ĭ���`� ���ĥ���R�q̅/�t̅ ���1��0�/��e������ % �� )������愩���/�0�ө�0�R�q̅/�/��
e����&�� )���e������ )������愩���/�0��`  @ �ȥ)��)
�<�) �H�)��0`L��LSͥ��掦�䄐� �������"� E� ��`��F`����Ǝ��ᦄʆ�L�̥��w��E���R�w� � �"� E� � Eআ�$�c�@�#���������i#� ?� C� � C�憦����� �� �˥������掦�䄐� �� � �ͩ ��``���1���� � �R�t�% �� ���ƅǩ"� E� �� ɦ�@� �`L�˩	�E vȩ"� E� �ϩ ���������� g�` �ͩ#�b�@�"���������"� ?� C�`��� � �/� ���� �/�� 


���/�!��" �#i��`���8��� � ��� �	����� ����`��
��1΅�2΅l 5��Υ�'����"� ���ǥ�ņ�������R�S���L`��` � E��� jʥR�E�ǽ���� ��8��"������
��.���/���R���e���Ʊ}���ȱ}���Ȅ!�R


� ��Je ��R���e����Ν@�@� �!�� � ?� C�`	



	 � E� v� � �� ɦ�@�  ?� � 4� C� �� �� g� � "�`�R���e����� `�R��ˆ� ��� �  �֤�!���"������
�� � ���!�"��0�!�&����!���"�����
���������
�� ��`���"��Ӭ�� )� ���R�w� � `�R��ˆ � � �����
��� ����� � � ��
��`� Ⱦ�� )� Ć��`� ��������������������`LyЦR�w̄ ��˩
�!�� % ����!��R��S� ��R�͕��͢ � �S���������� �S������͕��4�5`� �����R�R��� �R�R�S ���`�
��R��˪� �!��" &�$


���#�!��" �#i�����ԦR��˅�
�� �%��& �� � �/�% �� ����'������R��˅� ��R���e� �� �%��&������%i'�%��&��� �%�/��'�����
��`����p�!��"���#�$�$ �L��`�G���	)���dI��d` �ۥ�
���х��хl �ѣ�\�m�q֩ �ȅ�Ʌʅ˅����`��
���х��хl ���ӎ��-�@��2� ����` � �� ��`� ���R���e��� �� �ԭ
�	 +� �� $�悥��
��` �֩ ���R���e��� �� (�悥��
�� w���`� ���R�t̅ �q̅/��0�/��e������ % �� )����m�e�������/�0��` $*06 g� �Ҧ����"��� ��



e"�� �����"􅪢 ��`� ����ʤ���



��ù �  �֥!�#��e¨� �  �֥#�!��#8�!�����ʥ�����
��`�P)���J����� `���	���� `�� ` �ҥ�� ��`��`���� �֩ ������`L�ӦR�w̅ ���<�e�����膯�R���e��� ����� � )� ���  �  �� wҥ��ː9�7���  �֥!�#�"�$���  �֥#�!�� � L�ө�� � 0�ʅ˥���������� )� �R�w̅ ���  � �R���e����� 櫥���� ��欥��
����`L@ӥ�0"�� gȤR���e��� ������������` ����`��� H��` $*06� ���/��������/��
e����"�� )���e������ )��������/�/���`�R�R��`� �R` E� P֥���� ���� �Ԥ��� � ��y� ��
��� �Ԥ��� 8��� L��槤����` FԤ����� �/�ե��
� ���
�Ƅ��� ������� �������`ƨ` %+17=CIOU�R�t̅� �#�$����
�� %��  �֥!�#��
�#�"�$�����U�հ�"�$���$�����
�!`� �!�"����"�!��`� �#�$����$�#��`��� ����/��



��!� �! �ե"��!������



e/��!� �/��`� �"���������#���ս
�$�
�!��#��樥����`�$�"`� � � �ࠐ�`���
���R�B�9 � ���[��`���� �������`� ��
��U��`� ��� ���ƅ��` 5�`���� �Ω ��`� � �R��˽ �" �դ �"���!���� � �
��`� �����
��`� ���p���������������̥ʅ˥���`� �p���������������̅�`� �����<��`� �/�0�R
����������/�;�e0��� ��/�!�0�"L:��0�0��ީ �0�/�/���` (<Pdx������ �!�"�!�<�e"�����"�"��� �"�!�!�
��`��������R���e!�� ���!��`��
���ׅ��ׅl ��n�t�w؟إاة �������R��˽ ���w̅�� ��e��� %����`���ꭠ���`�R
���؅�ȹ�؅��R�t̅���e����� %��� )�����泥�e����� %��	� )�泥����`�����������L�إ���L�ؤ�� )� ��� �� �R��˥�� ��` ����`��` wҥʅˤ�� )� ��� �� �R��˥�� ��` ����`�� wҤ�� �� ��� )� �R��˥�� ���ː��������� gȤR��˽ ������������ �������`��`��������*�& ک ���R�� �	���� )� J٥ � e٥ � �����`� � �R

�� ���ſ������� `� � �R��˽ �!��٠ ����!������� ` ���Xk~\q�����CVi|I^s�� ��ſ������� ���R��˽ �����������`� ��R��ˆ�� �� Fԥ��� ��ſ���������
��`��������������`�R��˽w̅!�
� � ���� %!�
�R���� ��`��L0ڥ�
��Lڅ�Mڅl P�/��]�]��� �]�8i�(� �'�(�
�� �(��'�'i�!�p�"��# mߥ(i�!���"��# mߢ ��0
���u^�^�Y���� ���` (Hh� �� �/�0�1�Y �d��d�Y �/�Y �
�	�
�Y �0���1 �������`� ��/i�!�ۅ"��ۅ# m������`HXh(Hh��!�X�" m�`� �! m�`�. b� ���8�5�8�g��P���`� �8�]��4 ��`��4 ��`�Q� �^�^ �
����� �\`� �^�^ �
������\`� � ���\`�Q�^�_��`��^�^��f`� �f`�_�`����f`�Q���f`��f`�P��
���4�5`���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �!�"���#�$ �` Iߥ!JJ

�!�#JJ

�#�#8�!JJ�%�%�$8�"�&�&� ����%�� a��&��`�!JJ��@��"�	�0 a��0��`�i0���`��!� �"� �#� �` I� �ߥ7
�� ��/���0� �/�!�# �߱/�" �߱/�% ���#�� a� �ߥ!�#�"��`��%��&`�/��0`�%��&`���`���<�� ���a`� ��`�  I����I�%��`� �#�!��"��#e"�#�!��`� �#�$�!��"��"�!�#���$`� � ��� )@�� � �� �`��@�䣅
�'���(����!���" Iߥ�%��& �� � ��/�%L��%�/ �� ���'� aߥ�%��&�
�'�(��`�
�����/����0` � 	�	 
�
 � � � � � � � � � � � � x x  @`����  @`����  @`����  @`������!)
� �$���" Iߥ�%��&��@�䣅
�!����"�@
��8��/�-�9��0�.� )�� �1���$�_ ?� �'�(� �/�# ��#
&(�$��'�# �#�%�1�(�'� �(� �$ ,� ���!�˥'�# �#�%�1 aߥ�%��&�
�!�"Т` ?� �/�# �� �#�% ,� ���1�!�� a��1��%��&�
�!�"��`�� ��`�/�/����0`�� )
�� �W�+�X�,l+ ��_���-�/�.�0�8�"�)��
��L�� ��*��e
��0e/�/��0`�-�/�.�0�"8��) ��*L��-�/�.�0�"�) ��*��L�� �*�)��*e
�*��0�)��`�� )�,� ��#jjj)���#

)0��#JJ)��#***)�#� `�H�
�����2����3� �1�2=E�)����� �#=E���#)�#���� h�`�0?���� � �%�/�#���#�%`��!���"��0�$�����%`� `�!8��%`� � � �* �G�H��� ���E�F`�
���������� ��(�)ȱ�*ȱ�+� ȱ�,ȱ�!�+�"�,�# mߥ+e-�+�)��(�)� �+�,e.�,�*��`�	����� �`������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�������l ����l�u�~�����-�. ������� ���` ���� ��`�`�	)�)�&` D� ��!� �"�%�# m�����`_ac`bd(Px D� �"�!� �"�%�# m�����`� �!�(�"�7�#���$ �`�H�!�(�"���#���$ �` �� D��` �� X��` �����-�. ������� ���` ���� ��`�`�	)�)�` D� ���!� �"�%�# m�����` D� ���!� �"�%�# m�����`eg_fh`��L��`���� � xآ�����&  O穠�  � � � � � ���5�� ��ԥ���5� o�LJ� �� �� �� ���L,��� ��� ��������������`�5�� �5 ��4���? "�  � �� �� ��`� �� ��@��` 	��%� �6�6� �7� �!� �"�6 �������`�4�1�& �4
�������� � �/�*���@�0�0�) �߱�# �� ;��)�0����)�) �߱�# ;��)� ��L��ɍ& `�����������/H�0H�4
��������#)�
���%ȱ�&� � �� �%�/ �����
� �� ��Lf�h�0h�/�/i�/��0�*�*��� �*�0�/iX�/��0� `�/i.�/��0`�4
�������l  �����`���;� �����R�����R�������h�Ե޺����U��ű˲ѳH�H�H�� ��� 6� |��h�h�h@ m��9�=�>ȱ9�e� �@����0���@�eJ��?� �@�@��� �* ���`��� ��� �  �ޥ?
��7�9�8�:`� �@�@� �@�@����>�
�=�>��`
��7�9�8�:�
��9�;ȱ9�<��� ��G�� 5�L�� ��L�� �� 0]��;�eJJJ���� ��G�Bȱ;�3�

��3� �e)�6� �� �!JJJJ�$�)pJJJJ	�0 h� �e u�`�@�-�>�����k�L���*��$8�'�$���)�* h� ��`� �-�$ h� ��`�*���'}$�$����)�* h� ��`�-�e�e u� h� ��`�*�Ž$8�'�$��!)�$L��!)�$���ǽ)�* h� ��`�*� h� ��`�@���)��e�0��)pJJJJ	�0�

��)�%�38�e�3��6� �3�6�3� �6� `�3ee�3���6�6��ީ�6���3��~i�@�

��f� `�e���@�-`
eee@����e��@)�*�JJJJ�'�e�-`��;���e`���ȱ;������.�@���*��� ��� �  `��ý	��	��L����ȱ;��	�L����ȱ;�L��
q;e@�e����eȱ;��@�L��E05

����E�� � �b��d)� � �c�� � �� � �G�G�c�d�S)x�OJJ�e�b��c�C��?�d0&�b8�e�b�
�c� �b�c�b� � �c� � L��eeb�b���c�c��ܩ �b�G�� � � �F0

����F�/�( �0�) �H�1�* �H�	�H�� �* `Dj!=)m!Q|#3� 8(
� X P)
�8ʈ) o	 X M�����]���_�����q���S���#�	.	.T@	.������  	.	.T@	.@T@T}!�	0� 	�	}	T	@	���������  ��� � �   ������ �� � � � � � � � ����  ր   ��#X�
<	� 	� <�#X�
<	� 	� <�#X�
<	� 	� <�#X�
<	� 	� <�"�@	�	h 	} ��#X�
<	� 	� <�#X�
<	� 	� <�"<	}	@ 	T }�"�@	�	h 	} ��#X�
<	� 	� <�"<	}	@ 	T }Ā   ����e#�� �� � �  _���e#�� �� ��� �  _�����e#�@� �� ��� �  _���e#����  ������      ��X<�<�<�<X<�<�<�<X<�<�<�<X<�<�<�<��}�h�}�<}T}@}T}X<�<�<�<X<�<�<�<  ���e#�� � � � ��� ��� � � � ����    @ @T@  @ @T@}  �}T@��� ���@�  ��� � � � ���B< � � � � ���A� � � � � � � � � X < X < X < X <   ����2�X
�
�
�
<	�	�	�	}	T	@	����e#�AAT!@!}A�!}!T!@!!T!}A�	 	 	 	 � � � � ���@� � � � � � � � � ! � ���@�  � �  ��        X�X�X�X� � � � �x<x<x<x<X�X�X�X�X�X�X�X� � � � �x<x<x<x<X�X�X�X�X�X�X�� �  c��� �   �����������������������������������������������0�   �   <��T}��}<<�}��<�}�T}��}��<<�}��<T}�}<�T}��}���<2<  I���	��		T	@	}	�	T	�	}	@�	@	}	@�	@	}	�	T	�		T	�		T		T	@	}	�	T	�	}	@�	@	}	@�	@	}	�	T	�		T	�		T	���		@	T	}	�	}	T	@		@	}�	@	}		T	�	T	��	@�  ��	T	�	}	�
<	�	T		�	}	@	}	�	}	@	}	�
<	�	T		T	�
<	T	�	T	�	}	�
<	�	T		�	}	@	}	�	}	@	}	�
<	�	T		T	�
<	T	�	T	@			T	}	�	�
<	�	�	}	T	}	�	@	}	�	T	�
<	�	T		@	}<  ��3��� ��� �������@� ��� �����@�T�} ��� �������@����������@�T�} ��� �������@������� ����� 2��!�!�!�!�!!!!!@!@!@!@@@TT}}!�!�!�!�!!!!!@!@!@!@@@TT}}!�!�!�!�!!!!!@!@!@!@������<< ��� �2   ��� ��� ��� ��� ��� ��� ��� ��������� ��� ��� ���@�   �    d  <�}<�}}���<�}�T��}��T�����  <�}<�}}���<�}  ��c���T@!T@!!@T�!}"<T@!T@!!@T�A}T@	 T@!!@T}!�!T��!���	� �!�!�B<}T	@ @}T!@!T!A�}T!@}T!@T}�TA}��!���!���!}"<!T@T!}.T!}1�@T  �}� @  �@#X"�"<"�"�#X#�"�#X"�"<"�"�#X"<"�#X"�"<"�"�#X"�#X"�!�"�!�"�#XC�"<!�"<!�#X"�#�#X"�"�"�!�#X"�#�"<"�!�"�!�"<!�#�#X"�  2�X  �"�"<A� "�"<A�  ����2�����!!}T	.TA}��������! � �  �������� ����AT	.T} ���� �  ���!!}T	.TA}��������! � �  �������� ����AT	.T} ����.!    �@A���<�CX<�<�2< "<"�A�\�\�2\ "\!�1� �<�<CX��<�B�\�\�!�"<!�"<#X"�#�"<"<!�"<!}!�"<"\"�"�!�"\!�!�"<"�"<#X"�!�"<"�"\!�    e����@T	}�TA����A@�@AT@	T  6}�!}"< }TA��	�}�B<�	}T}A�}	T@@�����A@	@TA}T	@TA��	���@ !@T	}�TA}  �@#X"<"�"<"�!�!�"<"�#�#X"�  ,"�!�"<#� "�"<B�"<"�"�#�"�#X"�"<"�"�"�!�"<"�"�"<"�!�"<!�#X"<!�"�"�� � � "<"�"<"�  w�����1}.}.0����`� ��2\�\�2\<\<b\ ������@@� .h@.A ����.}.�.�@�   ���& ��� �E�F� � � �* �G�H� � �< ����I�[�J� �K�L��M��& ��M���M A� ���K����L����i<���`�I��I`�I�K�>�]�:��8�K ���i0�N�i �O�K�����N����N�i0�N�O�i �O���K���  ���K�a�.�]�*�D ������ȑ���� ��i0��i �����I� �K�_��a�Ș ��K�a����K`�K`�J��J`�L�K�]�G��8�L ���i��i ��i0�N�i �O�L�����N����N�i0�N�O�i �O���L��� ���L�a�0�]�,�D ����ȱ����'��� ��i0��i ���ߩ�J�L�a����L`�L`



}/��N�0�i �O�J��� ���3�e��i ���N���`� � ��@�� ��������`H)�����hJJJJ�
ei@}��` 0`��� P���@p��      

�� �'�� � �����`� �/ �5�5� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ � �