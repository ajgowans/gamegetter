                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                H�Z��Y ��Z ��[ � �U ���W �W �T �U �S  pԬW �r� $��W ���V ���X  $��W �W �T �U �S ��Y ��[  p��X �X �X �T �V �S ��[ ��Y  pԬX �D� $ـ� $� $٭W �T ��[ �U �S ��Y  5��U �U �S  pԭV �S ��Y  5��V �V �S  pԭV �� $ـ�z�hL� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              �����������������������������������������������������������������[UUU����������������������������������_UUUU���������������������������_����W�VUUe����������������������������i����_UUUUUY��������������������������������UUUUUUU��������������������������_Z�f��W�UUUUUU���������������������������jU��_UjUUUUUU���������������������W�������UUUUUUUe����������������������UV������WUUUUUUUi�����������������������h��YU�UUUUUUUUi�����������������������`�����_UUUUUUUUY����������������������d������U�VUUUUUUU�����������������������j�����|U�UUUUUUUU�����������������������������\UjUUUUUUUU�����������������������������WUUUUUUUUUU�������?T�������������������|WUUUUUUUUUU�������j�������������g�����\WUUUUUUUUeU��������U�������������g����?WWUUUUUUUUeU�������d��������������g����?UkUUUUUUUUiU�������T
T������������g�����UnUUUUUUUUiU�������S@U������������g�����^UUUUUUUUiU�������?���������W���g����w�^UUUUUUUUYU�������uU������������g���uU]UUUUUUUUUU��������]U�������  ���gU��UU]UUUUUUUUUU��������UU������_�*jU�gUUZj�U]UUUUUUUUUU�������VU������e����U��UUUUUUUUUUUUU�������?�������������WZYiUU�UUUUUUUUUU���������Z�������W���i��V��j�WUUUUUUU�U����}���Si�������e����ZeUU��j�WUUUUUU�U�������������������AUUU�YUU���YUUUUUU�V������������������_@UUVUUU�ZfUUUUUU�V������������������iUUU�UUUUUV��UUUUUU�V�������@U���������UUU�UUUUUY��WUUUUUUU��������?TU��������_VUUeUUUUU����UUUUUUUU����������������YUUeUUU�VUU��WUUUUUUU�������C�U]��������eUUXUUUY�UU��UUUUUUU�������@_Ue���������U�VUUVUVUV��_UUUUUU�������XUUe����������?XVU�UUYUV���UUUUUU��������U�Z���������?XVU�UUVUYj��_UUUUUU�����c�Zf����������V���UUVUVV���UUUUjU�������V��������������UUiUUVUVVU��WUUUjU������?�j����������?`iUUUUUYU�UU��_UUU��W������TV����������PVUUUUU�UUUUU�UUU����������������������UUUUUUUZUUUU��UUU� �������������������gUUUUUUU�jUUUU��UU= �_������������������XU�UUUUUU�ZUUU���U=T������������������?��UjUUUUUU�ZUU����?Ta�����������������?VU��ZUjUUUY�jU����?T�������������������V�UjU�UUUU�j�VeU���T��U����������������SeUU�Zj�jUUeU���VU��T�W���������������UYUUUeUY��V��VYUUUU�S�WU��������������UV��V��VUUY�U�Z�UUUUYU�_U�������������_�UYU��eUUUe��ZU���UUUU�UU������������_eU��ZZVUUUe��UU����UUUZUU�������������_Y�	 �YZUU��U�U������UZUUU�����������_Y�	 �ZZUUU�V�U�������UYUUU������������WYU  ZZUUU�V���������UY�UUUU�����������WYU  ZZ�jU�V���U����WY�UUUU�����������WYU  �ZV�V�V���_UUUU�_U�UUUUU����������WeU) �����Y�����UUUUU���UUUUUU��������UeU% ���	 �����UUUUU����UUUUUU�������UeU% ��e h����_UUUUUU��_�VUUUUU�������UeY% ��i Xee��UUUUUUU��_�jUUUUU�������_UZj	��UY �ie�UUUUUUUUUU�jUUUUU�������W��U	��Ue �Ze�WUUUUUUUUUUUUUUUUU�������T�e�`i�� �V��UUUUUUUUUUUUUUUUUU������?PeY�X�Y� �U�UUUUUUUUUUUUUUUUUU������Te�� j�Y� jU�UUUUUUUUUUUUUUUUUU�������g�
 j�Y��iU�UUUUUUUUUUUUUUUUUU������P�o� �h�Y��Y��_UUUUUUUUUUUUUUUUUU�����;��_� $h�e��V��_UUUUUUUUUUUUUUUUUU���� ���%h�Y��Uj�WUUUUUUUUUUUUUUUUUU���� H����HiiY�d�U�UUUUUUUUUUUUUUU��UU��� R���?BijY) ���UUUUUUUUUUUUUUUU�VU��������?@Z�Vi ���UUUUUUUUUUUUUUUU�jU���  e�����VUe ���_UUUUUUUUUUUUUUUU��U��? HY�������O ���WUUUUUUUUUUUUUUUU��V�� PV�U��U�� �UUUUUUUUUUUUUUUUUUU�Z�� �U��@������_UUUUUUUUUUUUUUUUUUUUU�� UU�P�W����WUUUUUUUUUUUUUUUUUUUUU�� @U�_�? �������WUUUUUUUUUUUUUUUUUUUUU�� @U�W�? ������UUUUUUUUUUUUUUUU��UUU�� @U�w� ��UU��UUUUUUUUUUUUUUU����UUU���PU��� �wU�� ��UUUUUUUUUUUUUUU����WUU���V�����_U�� �UUUUUUUUUUUUUU�����_UU��V�_�� ��UU�?�_UUUUUUUUUUUUU������_UU��OV�_�@��WU� �_UUUUUUUUUUUU���� �_UU����W�?@�UU�?D�WUUUUUUUUUUU����  �UU�����W�P��UU�O@�_UUUUUUUUUU����   ��UU�����W�_�_U���WUUUUUUUUU����   ��UU�����u���_Uu���_UUUUUUUU����    ��UU��������UU����WUUUUUUU����?     ��UU�����?��WUU���WUUUUUU����?      ��UU���_�P�UU}�G��UUUUUUU���0   0  ���UU������P�UU���WUUUUU�����   0  ��jUU����W���_UU��G��UUUUU������   0  ��VUU����W���WUU���_UUUU���?��   T��VUU������P��UUU���UUU����  �  ��U��VUU������T��WUU����UU����  � ���UU�ZUU����?T�wUUU���U����?   � ����UU�kUU����?��UUU��������0     0����UU��UU���_���WUUU���w��� �     pU�_�WU��VU�����C�_UUUU�������  �    @�U}U�_U��ZU����S�WUU��������   � CU�UUU�_U��kU���u�S�WUUUU�����?   �? WUUWUU�U��oU�������]UUUU�_��?�?   �?UWUUWUU�U��U�����UUUUU��? �? �� �UWuU]UU�� ��V��_�_�UUUUU��? �? �� �UWuU]U���  ��V��_���UUUU���  �? ��T�_UW}UuU��� ��V������_UUU���    ? ��UUU�U�Uu��� ��Z��W}��WUUU��   0 0 ? ��UUU�U�U� ��� ��k��W�UU���0   0 0 �P��UUU�UU� ���?  ����W�_U���0   0 0 �U��WUUUW   ���?  ����U�wU��� 0   0 �@�U��WUUU   ����  �����?�_��� �    �U�U��WU    ����  ������W� � �  � UW�U��W? 0   ������������U  � �  �UUW�W�� ? 0�? 0 �����������U  �  � �_UUW�WU� � ��� 0 ���������}WU  �  � �_�U]�_ ���  �� � ����������]U  �  �W�_�U]?  ?0� �� ����������UU  �  �W�_�U5 �   �� ����������U���WU �� P�W�_�0 ��  � ���������������UU ��PU�_�_�0 �?  �? ��������ZUUU�_�WUU? �_WU�_U�� � 0  �?����������ZUU���WUU= UWW�_ 0 �   0  ���������VUUUUU���UUU=@UUWW�?      �  ����������ZUUUU��wUUU}UUUW�?      ��������jUUUUUUUU��_UUU}UUU� ?      �����������UUUUUUU��]UUU}UU� � �   �������VUUUUUUUUUU�_WUUU}U  � � �?  ���������ZUUUUUUUUU��UUUU=  �� � 0�� �������VUUUUUUUUUUUU�UUUU=     �0�� ���������VUUUUUUUUUUU�WUUUU� �   ����������VUUUUUUUUUUUUUUU�WUUUU� �   �����������ZUUUUUUUUUUUUUU�WUUUU� � � ��������VUUUUUUUUUUUUUUUUU�WUUUU� ��� ����������UUUUUUUUUUUUUUUUU�WUUUU� ��� ������jUUUUUUUUUUUUUUUUUUUU�WUUUU� �����������ZUUUUUUUUUUUUUUUUUUU�WUUUU� ��������UUUUUUUUUUUUUUUUUUUUUUU�WUUUU� ����������UUUUUUUUUUUUUUUUUUUUUU�WUUUU� ������ZUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUU���������ZUUUUUUUUUUUUUUUUUUUUUUUU�WUUUU������UUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUU������jUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUW]U��_WWU��_��_�wu��UU]��_�UUU�WUUUUUU��uUWwuWWUuuuWuuWuuWwUUU_WwuWWUU�WUUUUUU�]uUWwu_WUuuuWuuWuuWwUUU]WwuUWUU�WUUUUUU�]uU�uuwWUu�_�uu�uu��_UU]���UUU�WUUUUUU��uUWwu�WUuuWW�UwuwuUUU]UWuuUUU�WUUUUUUUW]UWwuWWUuu]WuuUwu�uUUU]�U]]UUU�WUUUUUUU�WU��_WWUuuu�wu��_W�UU}�W�WUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<3<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                        ��      �*V�V�V�V�V���*      �?�?      ��*�i��
����8����
� L�� V��`�X�*8����
����i��
� L�� V��X`�Y�*�i��
����i��
� L�� V��Y`�Z�*�i��
����i��
� L�� V��Z`8���`�i�`�l ��i�8��� ƃ`�l � � �� �� ƃ` �� �� � �`��S ��T ��] �� ���������5 ��`�� ��	�'0�'��S �� ����	ɀ�����T ��Z ��[ �^���Y  p��^�^���^`��Z �
�[ ��S ��T  5�`���(=�����03� ���0.� ���201� ���<0� ���������(0 '�`��`������`������(=�����03� ���0.� ���201� ���<0� ���������(0 '�`��`������`������������� '�`�����Z ��[ ���Y ` +,* �!� ���� ����� ��`�!� ���� 8���� ��`����ɯ�C��%���0����� z��i��+��������
0�� ���������� '�`�
� Q�����S �A�T  ����T ���8�T ��ɀ��`����ɿ�C�
�%���0����� z��i��+��������0�� 8��������� '�`�� Q�����S �@�T  ����T ���T `�	�#������P�i����� �d�	`�
�&��i����P�i����� �d�
`�����0� ���0� ��� ��������������0������` '�` �� č���
���� c�`�� '��� c�`8��� � ��`������3�^���B��iɀ�����T ���S �
� �����T ��� ������<�i�8�����������( ����� ��`��0 ���������T ��i�S  ����T  ��`�� '�`�������� c�`�i��0%��i�6����P��U����i��0����������8��������
����`�!���`��� '�`�����(0π���0� ��������3����������`���0��`��i�Z���`��� `���0��`8������`���� `� ��}���������� �����`"���	� ����`�� č`�����0	� ����`���(0��`�����
0"�0!�0!�0 �(0 �-0�70�<0� ��`����`����`����`����`������"� ����`�����
������ ���'� ��`���`��� '�`����8���`i��������&��$� ��i����������� �������`�!�`  ����,��*�`�����.��.�`�1������`�������8���`� �����������.��v�� ����ک �`�y���
����ɀ�8������`���`������� ���4� ��`�� '�`�����$� ��y늍�������� �������`��0��i�d���`�L�� ������ 0�L�� ������ 0۩	L�� ���LЋ ����� ���i�7�;�2���8��_��t��������������� �8����7�� ���7��` �������0#��2�
�P�
���`�������������<���ߩ�����8�������`��ĭ	�*� ��}����������� ����ݩ2�	`"��������������
� Z�� ��`�����(0��������
�� ���ܠ ���}�����P�i������ �����`i����&� ��}�����P�y��������� �����`y���䌍�쌍� ���к`

 �������9�` <����(��8�` ������
�d���;�` <����(�
����:�`�����EڭR �?�0;�����0� ���R �����i�������� �2��`ڭR ��ˀ������� 1�`
��Z�� ȹZ�� � �}��(0 '�`���S ��}�� ��ɀ����T  ����`8����� ��`��`�����i���� ��� Ȍ���: L� ��`����
i
����?8����� ��0`��+� ����� L� ��`��A�`��A���A��� ��%��<��B��i��i����� �`��i���A�i�i
��ٽ�i����i����Z� �{�������� 1� �z�`�{��S��g�����������`�i�] �i���] ��(���� 6�` ��` Ï`���� 3�` ��`���� ��` ��` ��`8�] �

�8�������`i����`8����`�`8��] 

�8�������`i����`8����`�`�`8�] �

�8�������
`i����	`8����`�`8��] 

�8�������`i����`8����`� �{�#��� � � ������{� ������������ѭm ��n ��n ��m  �π �Ҁ` � L��ýS�S �g�T ������Z ����[ ����Y  p�`�S�S �g�T ������Z ����[  5�`�� �` R�`�{
��Z�� ȹZ��	 � �}S0 �&�S�S ��}gɀ�� ��g�T `� �{`�S0�`�i�T �m8��T �
�(�T �� ��S �m�S ����S �] ����� `��������\�$ -�L!��������]�����L!��$���9����9��A������P�b ���N���0�$���0�a  � g� '����
� -���� [����
 `� �`���S ���T ��Z ��[  5թ��� � �ݩ����`�N��� ݒ`���S ���T ��Z ��[ ��Y  pԩ��� � �ݠ �������������S ���T ��`� ���޽� Ò����`���S ���T ��Z ��[  5�`�V��Y ����  �ߠ p�Z� ��z���� � ��`� U��R 
���� ȹ��	 ����c����$��� 3�`�R 
���� ȹ��	 ��
��� ȱ� ������c����` q��` ���!�F
 ���"�$` ŀ�Z�R 
���� ȹ��	 �"�z`Z�R 
���� ȹ��	 �$�z`� �� ݓ�!����%� �9`����`�!�� k�`�� k�`�� �`�� 4�`�� ��`���!� ��`�#� �`�$� k�`�(� 4�`�)� b�`�,� 4�`�-� b�`�/� 4�`�0� b�` �����'��� ���!�`��� ���������� �9���!�������`����]`��\` #-39? �����(���!� ����`ڢ ��"�i���i
��� ���9��������`�!� ��������i�0�(�$��`����!� ����� ��` ��� �!��i	�'0��� ���A�� 8������` ����!�8����� ���A�� 8������`ڢ ���%� g� ���� Ӽ����%�����`��� 8�`�� 8�`�� 8�`�� ��`�� ��`�� ��`�� �`�� L�`�	� L�`�
� L�`�� L�`�� L�`�� Յ`�� Յ`�� Յ`�� Յ`�� �`�� �`�� ��`�� ��`�� !�`�� !�`�� ��`�� ��`�� ��`�� �`�� �`�� �`�� Y�`�� �`�� �`� � �`�!� �`�"� ��`�#� �`�$� �`�%� h�`�&� ~�`�'� ��`�(� ��`�)� ��`�*� �`�+� �`�,� �`�-� �`�.� 0�`�/� �`�0� �`�1� |�`�2� �`�3� ��`�4� ��`�5� J�`�6� �`�7� <�`�8� �`�9�  �`�:� 0�`�;� E�`ccccccccccccccccccccccccccccccccccccccccccccccccc�ccccpcccccccccccccc|cuctct,ctctctctctct`ctctctlctectdctdctdPctdctdctdctdctdctectlctctctctctct`ctctccc&#&#c'%'%ccccc&#&#c'%'%ccccc&#&&#c'%''%cccc&#c'%ccc&&&&-$c''''/$cccccc&&#$c*)%c)%c,&&#c++(#c*$,c'''%c,cc$c(&#&#c**$+,c)'%c,+,cc(&#+$c++,%c)c+**-,c)'/c+,$c(#c+,*$c+(#c+,*$c)'%c+,,cc+,,cc+,(&#c+*$c)%)%c%)%c%c�pcc p`c p`cccpcc p`c p`cccpcc p`Pc p`Pccpcc pc cpccp`P@0 cp`P@0 ccpccpccp`P cp`Pcp`cp 0c 0@`c0@pc 0@`cpc`cpcp`P cp`P cp`Pcp ccp`P cp`P ccp`P@c`P@cp`c Pcp` c 0cp` 0c 0Pcp`cP cp`cPcp` 0c 0cp` 0cp `0cp cpc0c04c0c05c0c04c0c05cc14c1c16c1c15c4c1c17cc15c1c24c7c2cc5cc24cc27cc3c35c3c5cc3c36c3c34cc7c3c25cc2c6cc7c3c34c3c37cc5c3c36c3c15cc16c1c7c1c15c1c6c1c14c15cc05cc0c0�qcq cqcq
cqcqcqcqcpcpcpcpcpcpcp cpcpcpcpcpcbccbcclccbccbccbcb
cbclccbcb
cbcbclccbcbccbcclccbcbcbcbclccbcbcbcpcpcpcpcpcpcpcpcpcpcpcpcpcqcpcqcq������WUUUէ���ڧ���ڧ���ڧ���ڧ���ڧ����WUUU������������j���[�UU�[�UU�[UU�[U�U�[U�U�[�U嫪���������������թ�[��U�[��U�[��U�[��U�[��U�[��U嫪���������������_��[�uU�[��U�[��U�[��U�[�uU�[�_U嫪���������������U��[�UU�[�UU�[�UU�[�UU�[�UU�[��U嫪��������������Z��[��U�[��U�[��U�[��U�[��U�[UU嫪������������������[�UU�[�UU�[�U�[�UU�[�UU�[�UU嫪����������:�����������������������
��
�������������������������� �  < ���?  �����3�?3�? ��?� ���?<�� �0�< �������0�? ��P]������WU5]UyUyU]U]��|U   �  �� ��  _ �i� ���?\��֬��?�i� _ ��  �� �          P
 �*Pꯤ��P� �* P
 �
 Z/��X��� Z/ �
����3�3 � � � � ΀3�3���     �? ��0�
0 �0��2�02�02��2�00 0�
�� �?                 �0 �z �c� ʣ  ��  ��  ʣ �c� �z �0            � 0� 0�������:�c��Z���>����Z��c���:0����� 0    �3 �� 0 �0�  0  �0    �  �0  �  �  300 0 �� �3 <���<����������[UUU�   �   �   �   �[UUU嫪�������� �*�
  j�j� �VUUU*hUUUU�VUUUU�VUUUU�VUUUUUZUUU���UUU�
�jU�
  ���      <   �   �  �� ��� ���|�����l�������  �  �? �U� �� �   �  �  �  � ��� ����\�����l�������  �  �? �U� ��         �  � ����� �����W�l��l�������  l  �? �U� ����  ��O}U=  |U}��?  ��{��;  �v��?  ��{��:  ��w���  ��{��~����v���UU��{�꺪���w�������      p]�Z�Z�Zu���������z��w���my��{���my��v����z��{������w������{ �  Z	 �U� `UU
`UU%`UU�XUU%XUU
h�� �*  ������������^�^�z�_��}_�^�^^_�^W�^{W�^�������������^�^�_�^�}_���^���^{�^{{�^������������������z���ﭪ������^��^����� �* �j� `UU
XUU�XUU�XUU%hU�
�V�  �        �?    �;    ��    ��   ���  �n�  �?  |���  l��� [����W���������?|����?|�����_�����W�����  <   �  �� \� g����p��>p��;����W�������������j������=���f=����Z��������j���V� ��~Z9  ��Z=  ��V  �k�  ���   ��    �?    �    �    �   �������7����z�Zz�k� ��5 �[  �   <   TW  �m@�@��UU@WU@^�@^�@WU@�_@�z _�@uP���j�W\U�tUu�Um�UmtUut�ut�w�U= � @y[ �z��_�pUU�U��W��W��U����Э��W�  �ʲ�<2������.��²0�2�ú���.��²��2�����.�²��2�Ϻ�������. ?��� �2�������?X��j�����  ��*L5(������� ���Z�W�Z�W�n����������?  B ��  � � X����?(  �TP�ZUQ�n����������?.�²��2�Ϻ�������.����� �2��RA�+ P�P�ZZ��j���nUj�������������� P� U� T� T� U� E�@@� �W  �[P�[U�kUe�j��������������� P� U� T� T� U� E�@@� �W  �[P�[U�kUe�j����������.�²�<2������.��²0�2�ú�����? T�BU� @�PU�kUeꯪ������/�²��2�Ϻ���.��²��*��
����� ���Z�W�Z�W�n����������?*   �   
  .:  ��  2�  ���.�²��2Ϻ���.��²��2�Ͽ���   �   �  ��  ��  ��  ?̀�����>�����00�²����>�>���0>�����.   �  2  �� .� ²� 2�����   �  ��  0� ��� �>� ���0>�����/�²��2�Ϻ���.��²��2�Ϻ�������. ?��� �2�������?X��j��������?(  �TP�ZUQ�n����������? ����. ?��� �2�������?X��j�����²��2Ϻ���.��²��2�Ͽ�����������   OUUUO���O���O���O�U�O�U�O�U�O�U�O���O���O���O~��O~����������    UUUU������������o�W�_�W�_�W�g�W������������W���W����� ���  �U�?�>���?���?��_=��_=��W=��W>��>���?���?���?���?��O~�_O~�_O~�_O~�oO���O���O���O�U�O~U�O~U�O~U�O~��O���O���O~��O~��U>��>��e?���?���?��f>��>��U>��U>��U>���?���?���>��>��U>��U>��O~�_O~�_@~�_U~�o������������o�W�_�W�_�W�g�W������������W���W���?���?���?  �UU������������o�W�_�W�_�W�g�W������������W���W���_�_�_�_�_�_�_�o������������o�W�_�W�_�W�g�W������������W���W���_�_�_�_�_�_�_�_�_�_�_�_�_�o�_�o������������������������o�W�o�W�_�W�_�W�_�W�_�W�g�W�g�W�����������������������W���W���W���W������������������        UUUUUUUU������������������������o�W�o�W�_�W�_�W�_�W�_�W�g�W�g�W�����������������������W���W���W���W��O���O��_O~��O~��O~��O~�gO~�WO~�WO��_O���O���O���OUUU   ���������V�k�Z���W����������kի�[�[�k�[�Z�W�������������UUUU    ���������?���?���?���?��>��W>��W=��_=��_=���?���?��>��U�?  �������   �
   �Z��* �jU�U�`YUUV�
`UUUUU*hUUUUU�VUUUUU�VUUUUU�VUUUUV�VUUU�V)�UUU��
��ZU��   ���    ��  � �03�� � �  � �����:��;��:�U � � �  �  �  �  �  � �����:��;��:�V �? ?��0?��  3 �� �� ������\wpU��  ;  �  �� �03�� � �  � �����:��;p�5�U���  ;     �  p:  L�  C��P��������������� ���?�� �  �5  ��  �P�
@�������������� � ��  <�  �  p0  \�  W
��*�������������� � ��  �  � � � ������������� � � � ��� �� �?  � ������������ � �? �� �� �������������������{U��@��+)�.)�.)�+)�@�{U�������\U�: �:���⫪�����«������� ��\U�:���:������������: �> ��?� � ���?���������: �> ��?� � ��?�> ��? ���?������: �> ��?�®
�®
��?�> ��: �������?�� pU���������� ��  3 �� 0?��? ?�� ������������ ��  3  ?  ?  3  3 ��   ;  �  ���Up�5��;��:�� � � �  ���03� � ?  ;  ; �� pU\w�������� ��  3 �� 0?��? ?  �  �  ;��pU\w�������� ��  3 �� 0?��? ? �� �W� �������0���_U0������ s]� ��� �� �� �W� ����������� s]� ̭� �� < 3�����|U=����������>��:� �����^_�u~���
��   � ��x}-�U/�i/��+��
� ?? �<<��[����������    �           �         ��S��       ����� ��?  0����������  0������: �����������   ����_����    �U�կ����    �Uk������  ��?�h�j���9�   h�����:����j��������~�����������W>�ꯪ�< \UUUU������? �]�e��j��  ���j���ZU�  ���j���VP�   ��Z���@�   ��Z���@�  ���j���VP�  ���j���ZU� �]�e��j�� \UUUU������?�����W>�ꯪ�<�����~����������j����   h�����: ��?�h�j���9   �Uk������    �U�կ����   ����_����  �����������  0������: 0����������  ����� ��?   ��S��          �           �            0  <<         <  <0          0  <  <         <<  0     � �� � ����?������?�� � ��� 0��\5���Wի��\5��  ��?  ����  �� ��  �*  *<� ���0 ��������� ���� �����? ���   ���   ����? ��� ���� ��������� ���� ���0�*  *<�   �� � ����   ��?   ��?  ����  �� ��  �*  *<� ���0���������� ����� 쫮�� ����� ���� ���� ����� ����� ����������< ���� ���0�*  *<�   �� � ����   ��? 8        ��        �      �9�>      |���    � w~5Ͽ
��  \����+��  p���9�|>  ����9��  ����9֧  ����9V�   ���9V=  �?��~V-   ���oX�0  |U9���,  ��� �  p� ��� ���
�X�  ��`%�X�  �8`%�h�  �8`%
��  ��`%�� ���
`	�  p� `%�  ���c%�  |U9�c%�,  ���o�
�0 �?��~�.   ���9X=   ����9X�   ����9ا  ����9��  p���9�|>  \����+��  w~5Ͽ
�� ���    ��>      |�      �9�        �8        �,V�0WU������,V�0WU���0 �,V�,��������/V�,WU���0 ���,WU�� �����,WU���� >  ,_U����>  ,_U�����?�� ,{U-����� ,�������� ,  ���0��,30����0��,30�������  ��������  �T��  ���  �T��  ��   �T��  ��  ��T�?  � �3��T�?  �U�3��T�?  �U� ��T�  ��� ����?  ��� �Ϩ�  ��? �Ϩ�      ����     �?���     ��>��     ,�>  �     �?>         ��>         ,�>          >         ��?         ��         ��         ��         0�         0�         ��          �            �          �         �         �         �         �         �         �         � 0         �8         ��>         ��3     ��  �8     �����>     ���ÿ�3     ��?ÿ 0     ��*�/ 0��  ��*�/ 0��  ��*�+ �  �N�+ �U  �N�+��U  �N�+��?   �N�*  0?  �N   03  �N  �??  �N  �?3����?  �??����0���83>���?���8?>���0  �8 �?���?���8 �����0xU�8 �����?^U�8  ����0^U�8  �� �?�WU�8����� �WU�8���/ ?�WU�8[����3����8[�8/ 3�WU�[�8��?�WU�[�8�    ?       ��   ���� �ﯪ�9��0����9�?����������������Z�����������������V���������    ?       ��   ���� ��믪�9�?���9���������������Z����������������V�������������������������������꟮�Z��:�������:�������l�����l����� ����   �?��       �    �����������������������>�Z���:�������:��?�l������l����� ����   �?��       �     �  ��fx�=\�=��=W�>W��g�����pz>�� �  3  3  �  � �UU��jp��XY�9�V��U��[���[���W���\���3� 08  08  08    0     0    0   0�  ���  ���<   < � � ��� �  �� �� <p��� <p� � �p� � ps> ;��� ;�6���:����� l�� p��  ���9  �6W�:   �W�   lW�   ��    �    ��     �     �     �     �     �   ��  {� ��S����E�DU�T�,��;ke?���/\i�.F�.�nU<L�B�hU����T�~��?Tu��W��Zѿ�U��Y�/�go�)��;>  ,     0  0  �� ��������> ���������>��� �� ��  �������>���������?��� ��  \U ���pp�zp�p5p�z5���?���:���? ��    ��  ?��� ��������:�����;������������<�����<���������  ����  ����  ��������<�����<���:���������� ? ����3 ��0   ��?   �    �   �    ��   ���  ��  ���: 𪪿;����쫪����������������������������������<��������������:� ���� �� ?  ���3    0   ��?   �    �   �  ��   ���� ����� �����?�������������������<�����<����0��  ���  ���  ����0����<����<���?� �������� ���? ��   � ?   ���    ��    ��   ���  ���>  ����  ���� ���:����;����>�ê��:������몪?�﫯�����?�������<���?������ � �� ���  �    ��   � ?   ���    ��   �|_=5_=|�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ���ة��  ��� � �� � �� �ߍ& ��"  :٢ t ���� �� �� � ����� ��� �XL �H�Z� �
��
�	��	������������������������� �%��%���� ���ޣ����� ��� � �� x�z�(h@H�Z�' )��� �# �$ �% (z�hX@                                                                                                                                                                                                                                                                   ���  :٩��& L �����  �ߩ �˜c �d �e  ֩ �S �T �(�Z ���[ ��Y  pԜ�  }߭  ���� �˩ߍ&  h� �©��& ��`��Q �R �^ �_ �` �a �b �f �g �h �i �j �k �l �m � � � ��F���R �ȩ����[��P���` � �� � �� �� �˩��  }� Ví��  ��i � {� .ϭh ����� �˭R �
�I���  �� �����6�M��з���  }ߜM�Q � �� �ȭS�H���Q  � �ˀ� 8ր�` ��`�� 5� E� %Ω� �� k� |� �� $� n�`�[� �ǜ[��% �ǩ��[� � g� �� � ��� ��`ڭ��a�.� �U�R 
��H� ȹH� ����c������� gĀ,��8������ ���(���^� N� � �Ā��:С�`ڭR ��B��>�:� �2�R 
��H� ȹH� ����� ����(���^� Nŀ��F���`� ���i(� ���i � � ������`��!��$�	�`�R ��������
0u���0l� � �`���R ������	�	�
���������ɘ���>�c��`� �(��� ���R ��	��
�,���W�������  N����.Ж`� � �$�(��� ���S�% ���8�!�F��  N�`��.��`Zڹ������`�����z`� � ��.0	�:0
 �ŀ �ŀ �� m���F�ޭ� �í� �`�^�݁�	 �����`�^�݁�	 �����`�^�݁���A�� �4 �ƀ ����` .Ƚ �0\��!��!��������������` �` G�`��A�$���S�S������� Ô� �S`��ڭ��i
��0 h�`8����� ��`�S�$�����A�i����� ��S`�S`�S����i���A�i����� ��S` 5Ǽ���i(� ���i � ���� Z�� i)� � i � ��` 5��m�����i(� ���i � ���� Z�8� �)� � � � ��`�^�������
��A�}�� ȹA�i � `� m� � i � `��8����݁�� �  ��`ڢ � �`������ � ��������`��Ȁ���F���`� �`� ������`� �`� �������`��֍ ��׍ �N׍ ��؍ � ���
ȱ��(0�`ȱ��(0�`��׍ ��؍ �(�j����(�j���`� �F �ȹ|ȍ�� �����/�Y �^�Z ���[ ��T ��0�S  Fխ�Y  Tխ� ` �i��0��`�`�`�T ��׍ ��؍ �S �`� �� �� � ����� ���` � AʩH�S +� �ɩ �˭  ��	����  ��`��������  �߀���������  �� �թ �� �ɭ����V��H�S �ɀ���S ��T � ,�ڢʽc  ��� ����S ��T � ,Ԣʽ^  ��� �����S �F�T � ,ԩ�S �T�T � ,�`�
�S �S�T ��Z ��[ ��Y  p�`�
�S �S�T ��Z ��[  5�` ֩�S �(�T � ,ԩ�S �<�T � ,ԩ ��`�
�S �B�T �R �
�(i
 ,ԩ��X� Y̩�S �\�T �Q  �ө ��`��^ ma �^ �_ mb �_ �` i �` ؜a �b `�` �e 0��_ �d 0��^ �c 0 a�`�^ �c �_ �d �` �e `H�Z �� �ݩ �o  =ީ�)��&  �� �ʩ�S ���T �	 ,ԭ  ��� $� $� $٩ߍ&  �� �� 	� =� �ܩ��o z�h`� �S ���T �(�Z ��[  5� ��`��g � �`����`� � � � � � � � � � � �( �) �* `�����.����'��`� �R �Zˍ!�d� W���!����%� �9`685:685:<d7
<d7
��������Q�Q�F����N���`�N���� �� ��R �R �
� �˜N` �ɩ �� ֭N��� p �©��P� `� �� �˩��P� Y�` �� �����`� �Y  �����` �f �g ����Y ����Z �
�[ ���T �̍S  p�`��Y �ߠ ��Z �
�[ ���T �̍S  5�����`��Z ��[ ��Y ��S ��T  p�` � V�`�R ���  ���3��� tʀ*�� ω� ω� #ω� ω � �̉� ��`H�a� ������ �  �� � V� �� �ͩ�h`H 9� �ˬf �� �ݹg ����g �� `��	����n �f h`H��"1� �b����%���k �����b�i�n�i�z U�h`H�l �+��b�������k �����b�i�n��zh`H�j ���!��b���b�i�n�i
�z ��h`�l ��b���b�i�n�i�z`H�i ���!�
�b���b�i�n�i�z �h`�l ��b���b�i�n�i�z`� �b� U�����`� �b� ������`� �b� ������`�n�S �z�T �b��΍Z ��΍[ ��΍Y  �Э
 ���	� �b�
 ` p�`   	
�n�S �z�T �b��΍Z ��΍[  5�`�n�n�(0� �b`�b��	����`8�z�0���z`�n�n�(�`�ziɂ�ǝz`H��W�Zh`H��U�Xh`H��Y�Vh`H���h`�a�/ j� )� Y� ������m ��n ��n ��m  �π ��` b�` ��` ��`��Z ��[ ��S ��T  5�`��Z ��[ �_�S �`�T  5�`�n �B��Z �] ��[ ���Y �_�S �`�T  p� ��������.���5 ���n ��m  �π ���� � L��� 5�����`� IМ�U IМU�V IМV�W IМW`� Эm � ���i�_��` ���`Z��|�m���"0�"������mɀ�������z`���� �� �����'��#�f �f ���f  g� '� �� 	̩���  �ߩ `��S �i�T ��] 8���`� �� ��`ڭZ �] �[ � �����A����5��60-�i�����i��� X����T����  �� ���G 5����)����  ���.4�%� �*���%�" �� r� ~р ��������	 � L� r����
 �`������ � ��������S ���T �� -����`���Y �^�Z ���[ ���S ��T �Z  Fթ �  ��`� �� ������������� X����`����`� �{�#���S��g��������� X����`����`� � � ������^���� X����`��F��`ک�] ������׍ ��؍ ��������] �܀ ���`�m ��n ��n ��m  �π�a��R� jϩ�a�R`��8�a��2�ӍY ��Z ��[ ��S ��T  pԩ��� � ���a��`���M� ��`  ���S ���T ��� �������Z ���[ �V��Y  p�� ������m ��n ��n ��m  �π �Ҁ ���`���S ���T �����Z ���[  5�`Hڪ)�JJJJ�  �ӊ)�  ���h`xH�Z� �a��$��b��%��c��&��d��'����� ���� ��\ �T ��֍ �N׍ �S �- �� i� � i � Ȳ- �� i� � i � ��\ к�S �S z�hX`H�Z
��� ��	 � ��$�&�a��b��Z0��b��0�b�8�7�  ��Ȁ�z�h`�Z�Z �] �S 08�(�S ��i�Z �] �Y 
��A� �A� �Y ������	� i@� �[ �\ �S .8� �S �� m� � i � 8�] ��J�] �S ��@�T ���mS � �N�i � � �- ���] 0��\ �� mZ � � i � �ࠐ�z�`�� �  pԩ�� `� �  Tթ�� `�Z�Y 
��A� �A� �[ �\ �T �A�m[ :��Z �] ��׍ ��؍ ��֍ �N׍	 �S �- ��� i� � i � �] ���)0��\ ��T �A�ʀ�耩z�`� �  ���� �0�`�  ����`���Ս`(Pd������Z�� �� ���z�`H�Z� �@� � � � ����� ���� ��z�h` ��Q ��S �B�T � ,ԩ��X� Y̩�S �\�T �Q  �ө �� � � �� �˩��P� Y�`H ֩P�T �
�S � ,ԩ ��h` 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____Hq���>g���4]���*S|��� Ir���?h���5^���+T}���!Js���@i���6_���,U~���"Kt���Aj���7`���-V���#Lu���Bk���8a���.W����$Mv���Cl���9b���/X����							





H�Z�/���� ���� ��z�h`� �o �p �q  �� �ݜ � � � � � � � �* �� �� � ���� �� `�p ���%�� � �ݭ� � �� �  �� �� ͓ � �ڭq ���%�� � �ݭ� � �� �  l�� �� ͠ � ۭo ���X�p ����| � �ݭu � �v �  =ܭq ����� � �ݭ� � �� �  ���| �| �w � 7�� �� ͅ � �ۭ� ��� `�r �s�u ȱs�v ȱs�w ȱs�x ȱs�y )
���z ��{ �y )0� ȱs����� Ȍr �| �} �w � �L۬~  �� ��s � ��~ ��Ȍ~ �r ���� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��卖 �南 �� )0�� ȱ������ Ȍ� �� �� �� � �� �p � �� )�����q ��  �`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��卣 �卤 �� )0�� ȱ������ Ȍ� �� �� �� � Ы� �q � �� )��@К���p ��  �ڀ��� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��午 �卉 �� )0�� ȱ������ Ȍ� �� �� �� � Ъ��  �� ��� � ��� ��Ȍ� �� ���� 
���䍸 轹䍹 ���s ȱ��t `�� 
���䍸 ��䍹 ���� ȱ��� `H�Z�x )?	@�� �x I��-� �� �} �z��y )@��J��� �� � �8�� ��y )0� Ȍ} �z����} �y �} �� � z�h`H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����΋ �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����Ι �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����Φ �� �� �� � z�h`� `� `Hڍ� �� ���� �h`H�Z�� ���F�� 
��Dލ� �Dލ� �� 

����'�* ȱ�



�� �� ȱ��� �) ȱ�� �( � � =�z�h`�� �* `N�W�e�sށ�    
 (	� # 
 �� ���� ȱ��� ȱ��� ȱ��� )
��卭 �卮 �� )0�� Ȍ� �� �� �� � =ޜ� `H�Z�� ���Ly߭� �� �� I�� )��� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����ί �� �� �� )�� �� )����
�@����� �� �� �( �� ʹ ��* �� � �� ͫ � ��z�h`H�Z�  ܠ  ܜr �� ��~ ��  7� �� =� �� �ݩ��o z�h`H�Z�p � �
�q � ��� �� )?ͻ �N�� �H�� 
���䍏 ��䍜 ��䍐 ��䍝 �� �� � �p �q �� )�����q  ۭ� ���p  ��z�h` 80�!� 8�!� T�!� C�!� 8�!� T�!� C�!� 20�!� T��� ?�3� 2�3� T�3� ?�3� 2�3� 8�3� ?�3� C�3� K�3� T0���     � ��!� ��!� �0�!� �0�!� �!� �!� ��!� ��!� �0�!�     � ��!� ��!� �� � �� � �� � �� � ��� �� ��!� ��!� ��!� ��!� �� ��� ��3� ��3� ��3� ��3� ��3� ��3� ��3� ��3� ��!�     � ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� �!� ��!� ��!�     � ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!�     � K�!� q�!� K�!� q�!� K�!� C�!� K�!� T�!� _�!� T�!� K�!� C�!� T0�!�     � K�!� q�!� K�!� q�!� _�!� q�!� q0�!�     �

		�
	� ��� /2��     � �	� _�	� K�	� ?�	�     � ��	� ��	� �	� _�	�     � ��&� ��	� ��	� ��	�     � ��&� ��&� ��&� ��&�     � ,�&� ;�&� T�&�     � q�&� ��&� ��&�     � ?@�6� G@�6� ?@�6� K@�6� T@�6� _@�6�     � ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� ��&� � �&� ��&� ��&� ��&� ��&� ��#� ��&� ��&� � �&�     �
	�
�	�
	�
	
��

















����������������������� �  ��  ��  d���  $�  x�          ����'�c����	�E�{��g�o�|����S����b��K�X�d�m�q�v�|��������������������  ��)�5�PRESSaSTARTa$PRESSaSTART$CONTINUE$END$BEAM$SCORE$NUM$READY$GAMEaaOVER$PAUSE$STAGEaONE$STAGEaTWO$STAGEaTHREE$STAGEaFOUR$STAGEaFIVE$STAGEaSIX$STAGEaSEVEN$STAGEaEIGHT$STAGEaNINE$STAGEaTEN$CONGRATULATIONaYOU$SEEaYOUaNEXTaTIME$HIGHaSCOREa$YOURaSCOREa$�5�g���˜��/�a�g�k�o�u������	�I�^�s���ў�Q����@�A�B��ȟ
�J���ʠj������
�.���¢.�V�����ڣ
�:�j���ڤ�Z���ڥ�R�r���Ҧ��+�k����+�k����+���+�k����M�t���Ϋ��.�^�����֬��<�\�����ۭ�5�e��������5�G�O�����ǱW��w�W�7���8�@�踘�Ź�׺O�w�����O�߼o����i���S��i���S��  




	 |{~} &'pqrs"#$-./0123456789:;<=>?@ABCDEFGHIJtuvw!%K ����������cc                    !!!!!!!!!!!!!!!          !!!!!!!!!!                    cc#$$$$$$$$$$$()$$$$()$$$$()$$$$$$$()$$$$$($$****$$$************************$$$$$$$$$$%%%%%%cc���,�\�����,�\�������`��.����`��.��	 "$&(*,.02468:<>@BDFHJLNOc
 "$&(*,.02468:<>@BDFHIJKLNPc
 !"$)*+,-./02356789:;?ACEc "$&(*,.023456789:;<=>?@ABCDEFGHIJc	
 "$&(,067<>CHKPRTUVWXYcc�����������������������������������������
������"�&�*�.�2�6�:�>�B�F�$�&�*�.�2�6�:�>�B�F�J�N�R�V�Z�^�b�f�j�n�r�v�z�~��������������������������������������������������������
������"�&�*�.�2�6�:�>�B�F�J�N�R�V�Z�^�b�f��������������������������������������������������� �������� �$�(�,�0�4�8�<�@�D�H�L�P�T�X������������������������������������������ ����������!�%�)�-�1�5�9�=�5�6�7�J�����\�A�J�����\�A�8���8�j������8�j����9�cccccccccccccccccccccccccccccccccccccccPPOGGOGGNGNGGNGNGGG(F
P|2PZ< P
(<Z2(P <Z
(F2ZF(P2Pv(Ft <2ZvP <P(v <Pr2F
<
P2Z(<vP
(F<Zr2F
F
<Zv<Z2
v(<2P<Z2<ccccccccccccccccccccccccccccccccccccccccGG&GG$GG$NG&GGG&$G!!GGN!!G!!!$G!!!!!!!G!!!GG!!!!!G!!&!!!GG!!!!!&GNN$!!!!&Pt<tP2.tcp<t<^ <t(F<^(tP<<(P,2Fc<vbFdF f6Pd2<d <P<Z dd2dV2Z2FZ2c(P< (F( FfPP2<P<P2ZpF(P2P<F22Z<dFcccccccccccccccccccccccccccccccccccccccccccccccydy(yP(q<ZP2K2Z2FZVFy2ZB0XZ<yP2F2Z<Z2ZFqF.D\4JX@F2@zP@2@5q@2P@P(qP@5~@(@P*@FZ@2Z@~(P* R(P&rP7,7=y7(P7y7=,7(Z7qy(y,Z(<P<GGGGGGG&JJGGGGJJLfSfGfGfSJffJLfSQfQf!fS!f!!fQQ!!LG!fQSfJGf!!fGGfLSffJJGGGG!!!!!!&cccccccccccccccccccccccccccccccccccccccccccccccccccccccc*####*%%#%*#%,-*/0-.*&/*0,-##%%*2222-/22,0*##%%&,0-/&#%##%%#%-0,/F(Z<\<ZF\2Z<(P2PZF<((P<^2^F(P<<Z
<Z2Z
<PZFP2Z<P<P<P<
P<P(P22
P2F(PZZ<P(FZ<(Z<P(2F(<Z(FZ(P
<(Z2F
2(<Z2Z<P(2FP<FZ<
2Z
(P<2ZF2ZZZZ
Z
ccccccccccccccccccccccccccccccccccccccccccc!!GG/-*0,GG()()()()(!!!,0//))-/)()()(0)()()(()(,/-0)()30-3)(333-0G-0G!!!()()()()(,-)/0-(<PPF<p
Z<
Z2PZpPZ(2F<P2P2PFZ2PF<ZF(P<"F2 2Z2<F<F2ZF2PF2<(P(F22P<P2Z(Z(F2<BD8F2(Z2<2DDDZ(pZ(2FZFZ2F<P2^^Zccc ���� ��� �������   :�<�>�@�B�D�F�H�J�L�N�P�R�T�V�X�   �  �    
 


 









 
 

		(		

((((((( XYZUVW[\]^_LMNOST`abbPQRcdefcdeghiXXjkggxyggPggPz|{lmmnnmn ���������  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            R� ���