   �P�P�P�P������U�W�_=���_�WUW  ��p�P�ХP�ન�  00��00  P�P�P�P�P�P�P�P�    UUUUUUUU����    PUPUPUPUP�P�   �U�U�U�U�_�S�P�P�U�U�U�U�����P5PPUPUPUPU����                    �     �     �     �     �     �    �    <<    �����    <<    �    �                                               ��0�0�0��𪨪     �� ���  0  <,8<3 �3��3��3��<0<�� �  �?     UUUU     �� ���     <  <30�33�3  �3  �<�<�   �  �?     UUUU     �/ �� � �0  <  3033�033  33�30����  0  �     UUUU     �? �� � �0  <  3033�033  33038����  0  �     UUUU                �����������������������?               �WUUUU�WUUUU�WUUUU�WUUUU=               |UUUUU}UUUUU}UUUUUUUUU�              �WUUUU�WUUUU�WUUUU�WUUUU�               |UUUUU}UUUUU}UUUUUUUUU�              �WUUUU�WUUUU�WUUUU�WUUUU�               UUUUUUUUUUUUUUUUUUU�              �������������������������               _UUUUU�UUUUU�UUUUUUUUU�              �UUUUU�WUUUU�WUUUU�UUUUU�               _UUUUUUUUUUUUUUU_UUUU�              �UUUUU�UUUUU�UUUUU�UUUUU=              �_UUUUU_UUUUU_UUUUU_UUUU�              �UUUUU�UUUUU�UUUUU�UUUUU=              �������������������������              |UUUUU�WUUUU�WUUUU�UUUUU=              �WUUUUU_UUUUU_UUUU�WUUUU�              |UUUUU�UUUUU�UUUUU}UUUUU=              �WUUUUU_UUUUU_UUUU�WUUUU�              UUUUU�UUUUU�UUUUU}UUUUU?              �WUUUU�WUUUU�WUUUU�WUUUU�               ������������������������              �UUUUU�_UUUU�_UUUU�WUUUU�               _UUUUU}UUUUU}UUUUU}UUUUU              �UUUUU�WUUUU�WUUUU�WUUUU�              �_UUUUU}UUUUU}UUUUU}UUUUU              �UUUUU�WUUUU�WUUUU�WUUUU�              �_UUUUU}UUUUU}UUUUU}UUUUU              �������������������������                                                                                              ��P� � �Q��j�������?�����~��������������UUUUUUUUUUUU����UU�}}}_�_�W��        U]UWyg�����{�_UeUeU�U�Uz�~�_�U���w�_=���_�wW��W�\�|����{�^�WUUUUUUUUUUUUUUUUPAQ�$�%AAP_��߭|�|�~���_�u]�_���|�~���_u]�Z�UjZVVUAP�����?TP � � ��Ee�Z�Z)h*���*�)h�Z                                                                                                                                                                                                                        �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                    0 < ����< 0         ����      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ��.�� � �� �@�� ���.��.��}p�� ��}�� �� �@�� ��� ��� ���     � ���� ��� @�� q �� �@�� � �� ��� � �� �p�� �� ��� � �� �0�� ��� ���     � ��� ��� ��� ��� �`�� ��.�� � �� �@����.��T�� �p�� �� ���     � �� �@�� ��� � �� �p�� �� ���  �� � �� � �� ��� �P�� ��� ��� �0��     �.�� � �� ����  ��     �                                                                                                    ��� �� ��������� �� ��������� �� ��@������ �� ��     ����@��@ �� ��������� �� �����@��� �� ��@��f��     �      � �� ��������� �� ��������� �� ��������@ �@ ��@��     ����� �� ��������� �� ��������� �� ��@��@��� �� ��     �������� �� ��@��@��� �� ��������� �� ��������� �     �� ��������� �� ��������� �� ��������� �� ��� ��� �     �������� ��� ��  �     �                                             ��� K�� ��� �� T�� ��     �      ��       �     �� � /��     �                   �          �O"             "E" "u"e"��" "�"u"U"�"     "E" "E" "u" "E" "E" "u"                 "F" ""                                 "" "" "�"                                                         ��� ��� �
��.
�� ��� ��� �
��.
�� �
�� �
��.
�� �
�� �
�� �
��.
��     �T
��}
��}
��T
���
�����}��.�� ��� �
�� 
�� ��� ��� ��� ��     � _
�� 
��.
�� ��� ��� �
�� �
�� �(��.
� ��� ��� �
� �
�� �(�     �      �����������������@����@������������������(�     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ��                 ���                ���;                ����                >���               >�?�               �                 �;               � ?�?                ���               � 0�               ��?��              � ΀�    ��?         �    ? �        �   �         < ��   ?   0      ,  ��:  �   �  ��  �p�:  �    �  ��  � <�+  <      �� �0 ��:        ��  ���+         �   ����;         <   ���+ �           ���? �    �     ����; � �  �0     <  ��? � ��0     �� ��? � ����    0 �� � �  �(    ��  �    � <    ��
�� �0 <   �    �>
�� � �� 
     ���� �� �  �?  �>���� ��    ��  ���< ��   �?<   < �
 0 ��   �    ��  0  �     ��� 0  � �      <0��> 0  <0        ����0  ��     �     ���>0        0     U���?    <         ���
     � � �    ����:     ��     ����*     � ��     @����     0�  �     �����     ��  0     @����      � �     �����     �����     �����     �< ��     ���?     ;��<     0 0     �� �     0     ���� �    0     �����      0     0����     0     0�*
�     (� 0    �����      � 0    �����     ���     �*��     � �     �����          �����           �*��?      0     �����       0     ����        �     ����       ��     � �        ��      �             ��             ��          ��0��?         ���0���        ���0���        ��������?        ��������?      �        0      �� ��������?      >�                ��?                ��?                                                        �*                 ���               ����               ����               ����?               ����;               ����?               � ���               ����                3��              �<0�               � �               8��      ��     � 0��     � <   ���  �       �   ���<  �    �     ���  ��    <      ���p�?          ���<�*   �     0   � � ��;   �     0   < 0���+   0     � �  �?��;   0     ���   ��;    �   ���   ��.    0   ���  �?��?      ���  0���?    �� �  �� �?    ��8 �   <0 �  �  0�2 0   ��  �� 0  �   ����   < �      <���    �   0   ;���   ? �
  �3  � � 8�   ��     �  0��0�   �  ����  0�� �   <  � � �  00�: �   000 <   �  ��� �   �     0    ���   �     0    ����    �         ���?     0         ���     �   �     ��j      � <     ���:      ?00      T��6     ����     ���:             ���       �      ���:      ?�      ���     �����      ���     �< ��     ���     ;��<            �� �     �     ���� �    �0     �����      �0     0����      2 <    0�*
�      � 0    �����      �    �����       �     �*��      ��     �����     �0     �����       2     �*��?       �     �����        �     ����        �  ������        � ��� �           ��? �           �����           ����           ���0��?          �?0���         ���0���          ������?          0�����?      �    �   0      ��    �����?      <�                 �?                ��?                                                        ��                 ���                ����                ����               >���               >�?�               �+               0�?               � ?��                 ��               ��               �?��              � ���                 �                �              < ��
                p�/    ��       0< 0�>   �        0� ��*  �  0 �    �  ��;  �   � 0�    � ���:       0     ����: �           ���* �           ���? 0    ��    ����/   �<��   <  ��>   *�?��  �� ��   �� �   0 ��    �  ��  �    ��#<   ����    �<�   ����   ����  @���� �  �� �� �*���� <<   � ��  ���< �  00 ��  < � 0    � 0�   �� 0 �      ��  ��� 0 33      0�  <0��> 0 3      ��  ����0      ��:    ���>0    �3:    e���? <   ���2   ����
  ��   �/�   @���:  �?? ����   ����*   �� ��? �   @����   < �? �8   �����    �   0�    �����   �?  ��    �����   �>���(?    �����  � � � �     ���?  � �����     0 0  � ����#�      0   0 �����?      0   0�(��(�      0   0 �����       0   0 *���>       (� 0  �����>        � 0   (���:       ���   ����:       � �  ������         0����:         ������:0       0   �����>0       0    ���0        �    ��?00       ��    3��       ��   00<�? �         �������         ������        ��?�����?        ���������?      � �����   0      � ����� ���?      � ����?           �    0           (� ����           ��                ���                 ��                                                        �
                 ���                ���               ��??           ?    ��<<       ��   �??    �   0    �#��   �   ��   �� �   �  0� 0 ����  �   ��  ��0  �       ��?0   <0 �  �  ��     �? � � 0  ��0        � �   ��         0 ��    �  �       0 �0    �           ��    �       �� 0�    �?      �        �ߨ�   �  0       �Ϡ�    �   �    <  ���
          �  ��    �      <   �? ?   �    ��   �? �  0   �0<    � �?    ���     � ��/   *���     <� �   ��<� <   0� �  � � �  �+� �   ���#<    �����:    �,�   ��갪�    <��   ��:��� �  �� �    �:��� <<   �    �: ?��  00 0   �� �    �?0   ��� �    ��0   ��:  33   ���  ���� 3   ����   �� ��>    ����   00���� ��? �   00�����<  �:���   0P���  ��  � �   ���� �?? ��3   ����  �� ��? ;   ����  < �? �  �� ����   �   0  00 ����  �?  �  0 d���  �>���(  3 ���� � � � �  �� ���� � ����:  ��      � ����#>      � �  0 �����      � �  0�(��(�      � �  0 �����        �  0 *���>        � �����>        �  (���:        �  ����:        (  �����:           0����:         0  ������:        �0   �����>        �0    ���         �    ��?          �    3�0          �   00<�0            ����              �� �           ��?����        � ��������       � ��������       � ��������       � ����?              0���       � ����           ��                ���                 ��                                                                                                                                                                                                                                                                                                                     ���\���� �}� �.�� ��� ��� ��� ��� q��     �               ��� �� _� �.� �,��-��+��*��     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          H�Z� ������������ �����r� �Ʈ��������Ʈ������ ��ƬƬ������ �����D�	 � πL+� � 쥮���� π��i��� ����� π��8���� �� I� �� ���< ���z�h`H�W�d���	��
dd -�h`H�V�d���	��
dd -�h`Hd��	��
 ��h`                                  ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�                               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                �� � /2��     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                    0 < ����< 0         ����      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                H c�	�����! ����
�� ����$��& ��<����U ����P��f ����d��w ��<��"��%� ��d� �ɿ�2 �數���"��<��%� ��d��ݩ"��i��%� ��橀��������5 �數� ��"��d��%� �������"��8���%� ��ƩLc���Lc�h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   HکP�d�(����
JJ�	dd�(8�	���8�
� -��� 6���sd�(8�	�d��8�
� -��� 6���Sdd��8�
��(8�	� -��� 6���3d�(8�	�d��8�
� -��� 6������| H��iɠ��L� ,� �� �� �dddd�(�	���
 -� ��h`                                                   ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ����������������������������������?      ��������������������������������?        � ����������������������������?          ? ��������������������������� ���      � T������������������������ �����     �? T�����������������������  ������     ��@���������������������� ��������     ��U_��������������������  ��������?    ��@��W������������������  ������?��    �� �_}�����������������  ������ ��    ��P�������������������  ������ ��   ��@��_}���������������   ����� ��?   �_? �_����������������   �����  ���   �? u_�U__�������������   �����  ��   �� ��W}}}������������   �����  ���   �����_���������������   �����  ����  ��P�W���������������   ����� ����  ��@�W}�WW_�����������   �����������?  ��?@�_��__�����������  ������������?  ��?@�_�W_]}}�����������? �������������   �? ��W}�u���������������?����������  �? ��_}�u�������������������������  �� ��_������������������ ����������  �� �����������������?��? ����������  �� �����������������?�� ����������  �� �����������������������������  ���������������������? �����������  ��������w������������ �����������?  �������׵������������ �����������?  ��������]�����������?  �����������?  �������u�������?����  �����������  �����u}�������� ���   �����������  ����_}}��������� ��   �����������?  ���_�_}����������  �    �����������?  �� �_�W�����������?       �����������  �� �W�����ת�������       �����������  �? �W���湿������     ������������  �@������u�������� �     ���������  �P����_w��������� �     ���������  ��_����]��o�����?  �?    ����������  � �����w�}w��������  �?    ����������  �?@���w����������� ��   ����������?  �����_w����g������  �   ����������?  �����__�]w�������?   �   ����������  <����__��w��������   �  ����������  �����W_�u]�W�����?    �   ��������?  �������_}�w��������     �    �������  �������}]���U}���     �    ������?  �������W}}_��Wu�����          �����  ������_�u}���������        ����  ����_��W_�����_Uu������           �?  �����_��_������_��������            ������_��_����U���������  ������  �������_��_��W���U���������  ������  ������_�W��_����]��������   ������  ������_�_��������������   �  ����?  ������_�_}�_���W���������?      ����?  ������_���������������? �    ����?  ������_��W������W�������? �   �����  ����P�_���_�_��U���������? ��   ����� ����@�������WUU��������? ��  ����� ����?@���W�U����W�����������?  ����� ����?@��U�_�_����������������  �����?  ���� ��U��������U����������� �����?  ���� ��W��U���W��W������������ ������  ������_����_UU�_������������������� ������U����WUU�������������������� ����P��U������_u��������������� �����  ���?@��W������U��������������� �����?  ���� ������_��_���������������������  �������W���T����������������������� ����@����_  U����������������?������  ���? �����  @�_���������������������?  ��������� �? �����������������������   ���?����?���P����������������������  ����C������?@�����������������������?  ������������������������������������   ����@���������������?  �������������  �����������?��������?�   �����������   ������� �����������?  ��������������  �������   �������   ��   ������������   �����?   ����������? ����������������?  ����� 0 ������   ��   �������������  ����  ��������� �����   ���������� �������0  �����   �� � ���������������  ���0 �0  �������� ����?   �?  �������?  ��   0  �����   �� � ���������� ��������   �  �������� ����   �  ������������   �����   �?   ����������� 0 ��  � �   ��������  ����  ��  ����������? ��0 �����   �   �����������   �? �  �� � ��������  ���? �� 0 � ���������� � �� �����   �   ����������?   � � 0  �� �������?  ���     � ���������� �   � �����  ��   ���������� �  � �   � �������? ����   �    ����������<    < �����  ��� ���������� 0  �  ���  ��������� ����   ?    ����������     <�����  �� � ����������      ��  0   ������ ����       ����������  �   �3����  �� � ����������     ��?   �   ������ ���� �  � �����������      ������  �?    ���������� � �  ���     0�������  �����?  � ������������      �����  �   ����������� 0 �  ����?   ��������?  ���? �? < � �����������?�   ������      � � ��  � < �? ����?� ������������������������?  � ����������������������������������������������?����������������������������������?����?������                   �������������?������������������������?���������� �? ������������������������������������ ���������  �������������?�������������?���������?�?   �������������������������?��������?  ������������?�����������?���?������� ��   ����������������������?����������?  ������������          ������������ ��   ��������������������� ��� �������?  ���?  ����������������� �? �3������� ��   ���������������������??�������� ����?  ��� ����������? ���?0������� ��� ���������  �������?�0���?0 ������ ����  0�� �����������?����� ������ �� � ���������   0  �����?������������ ����  0� ? ������������������������ ��   ���������?      ����������?������� ����� 00  ������������  �������� �?   ������������   ��� ������ �����  ����    ����������?  �����  ���� �?   ���������  � � ��?  �����   �����  �����     ������������   ���?   ���� �  ����������   0 � ���  ���    ����?  ��?� �    �������������  �    �����������������?      ���? � �     ����  �?    0 �  ���������������   �������������������� ��   ������ �    � ���� ��     �  ��������������?   ��������������������  �    ���� � ������� ��   � � ����������������<�� ��������������������   0 �? ����������������� ��?   � � ������������������ ��? ���  ��   � �? <   < �� ���?  �����   �����������������    �? �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �� _��     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ���ة��  ��� � �, � � �- � �ٍ& ��" � t ���� �� �� � ����� ��� c� @� � �� ��Lt�H�Z ~��0 �0 ����0 z�(h@@  ����)   � :ɜ ���&  í� ����Ln���L��L� � �  �! �" � �1  �� �� ��ٍ&   � �̩��& � �y  � ?� �� �Ωu� �  �Ω�  _뜨  w� fɭ+ � ���+  _��+ � �����L��� )�7�� � �� %έ )п� )� � ���� �ĭ� �� I� � �L�­ )�  � z�L�© �y  � c� �� �Ҝ  r� �Э �����L��� )������ ,� �L��L�� ,� z�L�©�y  ��� �� �� �� ���  � ?� �� S� �� � �����L��� ����	 �� A�L��� �� ����� L���� Ͳ �i��
�� ͱ �]�[�� �� �� �� ��� �� ��  ��!� ��  �� �����	 ��
 � �� ��  �� ����и Ā z�L�© �y  � �� �� �� c� ���  J� �� ����� ������L��� ���� �L�¢ ���� zĩ �1  �� �� � �ƭ& � �L��L��H� �1  �� �� � c�� ��� �  ��(� �� � ��� �<� � ��� �P� � ��� �d� � ��(� �"� �%�  ����  �ɿ�> �ףּ ���"� �(� �%�  ���� �֩"� � i� �%�  ��� ��������? �ףּ ���"� �d� �%�  ���� ���"� � 8�� �%�  ��΃ Lv���Lv�h`H�Z� �1  �� �� � c쩹�& � �P�
 ��	 � � � �(� �
� ��Q�  -� ������|  H��R�  -� �����թ��& z�h`H�Z� �1  �� �� � c쩹�& � �P�
 ��	 � � � �(� �
� ��S�  -� ������|  H��T�  -� �����թ��& z�h`H�Z c�� �D� �� �  �?�%���  �� �ŭ  �� �! �� �" �� � ��L�ŭ� �! ���ϭ� �" ���í� �  �;�!���  �ŭ  �� �! �� �" �� � ��b�� �! ���ӭ� �" ���ǭ� �  �8���� �  �� �! �� �" �� � ��"�� �! ���֭� �" ���ʩ�� � �� �z�h`Hڢ �� �� ����� �� �� �����h`Hڢ �� �� ����� �� �� �����h`H c�� �� ��  ��� � ��� ��  ��� � ��  ��� � ��  ��� �-� ��  ��� � ��� ��  ��� � ��  ��� � ��  ��� �<� ��  ��� � ��� ��  ��� � ��  ��� � ��  ��� �x� � �� �h`H� c�� �� �	 �� � �F� �$ ��� �n� �
 ��� �� �%�  ��&  �ɿ�< ��& ���� �� �%�  ��& �ة� � i(� �%�  ���& ���������? ��& � ��� �n� �%�  ���& ���� � 8�(� �%�  ���& L.���L.ǭ& ��L� c�� �.� � ��� �V� � ��d ���� c�F� �� � �� ���� �� ���h`H�Z� �1  �� �� �� )�  c�� �� � ��� �<� �	 ��� �P� � ��	� �d� �
 ��<� �� �%�  �� �  �ɿ�B �� ���� �<� �%�  �� �ح i� �� �%�  �� i� �����L�����? �� � ��� �d� �%�  ��� ���� � 8�� �%�  ��� L����L�ȭ 	�  I� �����1  k� c�z�h`H��� �F�� �R�� �A�� �N�� �K�� �$�� �� �� h`H�Z���  6� ���&�$ �$ �L�ʭ$ ���$ �� � 8�� Lh����(��$ �$ �L�ʭ$ ����$ �� � i� Lh����&�$ �$ �L�ʭ$ ���i�$ �� � � Lh����(��$ �$ �L�ʭ$ ���i�$ �� � � Lh����	 c� ��L�����	 �� ��L����L�� ,� ȭ � �� H ?� �� w� ��h�  ��L�ʭ H� �  Y� ��� �	 � !�L����	 � !�L����	 0� �L����	 0� �L���� � � !�L���� 0� � �L���� 0� !� �L���� 0� !� �L�� 0� !� � �h�  ��z�h`H� � �  Y�h`H� � �  Y�h`H� i�  Y�h`H� 8��  Y�h`Hک� �	 ��
 � � � �� � � �  -�� �&�  -�� ���  -�� �  -�
� � � � ɐ�i�  -��� � ��&� � � �ީ� � � � � �$�i�  -��� ɘ���� � � �ީ� � �  -�� �&�  -�� ��  -�� �  -�
� � � � ��i�  -��� � ��&� � � �ީ� � � � �$�i�  -��� ���� � � �ީ� �� �$�	 ��
 ��  ��(� �p�
  ���h`Hڢ �  Y�������h`HZ�� 
��-�� ȹ-�� �� � ��U�� L�����f�� L�̩w�� �0 )
��� ȱ� � �� �����zh`Hک� �	 ��
 � � � �� � � �@�)���  �� -��|  H� �����ک��  w� ��h`H�Z� � )0�0�M� �� )ϝ � ��  �덧  �΀0��� )�	 � � �� � �3� )�	� Χ ��  �덧  �� YΩ��  w� � � � � �z�h`Hڮ � )��9� )��i@� � 	� �i0�  YΩ��  w� � � � � ��h`Hڢ � )0� ���� )�� )�	� �����ۭ )�� �h`Hڜ  �ή � �@��� �(�0�)� �� ��� ����� ��� ���|  H� ���h`Hڢ � ��8�H�i�h���� � ��8���
i� �h`H�� �� ��  ��h`Hک� �	 ��
 � � �� ��  �� ��� ��� �� ��	 ��
 L������ ��	 ��
  ��L������ ��	 ��
  ��L������	 ��
  �� ��L������ ��
  ��L������
  �� ��L������ ��	  �π����	  �� �π �� �� -��h`H� 8�� h`H� 8�� h`ڮ � �� Lu����Lu�����Lu�����LuМ$ �$ ���$ �$ ��LuЩ�$ �$ ����$ �$ ��LuЩ �$ �$ ���i�$ �$ �����$ �$ ���i�$ �$ �����`HZ� �� �� �� � ��� � ���� ���  � �����  �zh`ڜ � � � � ������`H�Z � ���&�$ �$ �L8ҭ$ ���$ �� � 8�� L$����(�<�$ �$ �L8ҭ$ �?��$ �� � i� L$����� �L8ҭ � � L$�����?�L8ҭ � � L$����(� �$ �$ �L8ҭ$ ���$ �� � 8�� L$����(�0�$ �$ �L8ҭ$ �?��$ �� � i� L$�ɿ�@� � � �3� 	�  <� r� ӭ )��  �� <� Ӎ � )�	� L8� ȭ � �� � H �Ң �  <���@��h�  r�L8ҭ H� �  <�h�  r�z�h`Hڜ � � )����"� ��!� ��$� ���|  H� ���h`H�� �#�  ��h`H�(� �	 ��
 � � � � � � �	�  -�1�  -�Y�  -𩁍  -�h`H �� ��h`Hڢ � ��8�H�i�h����8�H�i�h��K�� � )��[�� �h`Hڮ � )�$ � )��% �& �% m& � �"�� )�$ �� i� )0�0���/ L���& �& ��ȭ ��8����% �& �% m& � �"�� )�$ �� i� )����/ L�׭& i�& �1�ŭ ���% �� ���% ��0�� �% ��0�% � )m% �% �& �% m& � �"�� )�$ �� i@� )����� �/ L�׭& i�& ��ũ � ���� �� �0��0�% �� �	i���L�ԭ% i�& �% � �&� )�$ ��i@�� i@� )������/ L�׭% i�% �& �ĩ� ���� ��#�0��3�% �� �	i���L�ԭ% i�& �% � �&� )�$ ��i@�� i� )0�0���/ L�׭% i�% �& �Ĝ% �% � �i�@���% �% ���LNծ% � �&� )�$ ��i@�� i� )���	�/ L�׭% i�% �@�ũ�% � �i�4���% �% ���L�ծ% � �&� )�$ ��i@�� i� )����/ L�׭% i�% �4�Ŝ% �% � �i�@���% i�% ���L֮% � �&� )�$ ��i��� i@� )������/ L�׭% i�% �@�ũ�% � �i�=���% i�% ���L`֮% � �&� )�$ ��i��� i� )0�0���/ L�׭% i�% �=�ũ �% � �
i�@��L�֮% � �&� )�$ ��i��� i@� )������/ L�׭% i�% �@�ũ�% � �
i�=��L�֮% � �&� )�$ ��i��� i� )0�0���/ L�׭% i�% �=�ũ�% � �
i�4��LM׮% � �&� )�$ ��i��� i� )����/ L�׭% i�% �4�ũ�% � �
i�1��L�׮% � �&� )�$ ��i��� i� )����/ L�׭% i�% �1��L�׎. � )�	� �� � )���@��� )�	� �h`H�Z� � )�ɀ��$ �;� )0� ���$ �+� )����$ �� )��	�� ��L���@���$ �. �$ �/ �@�
�8�@��$ �� )�� �$ � �L#���L����L����L����L���	�L:���L����L����LD���L����L����L8���L��L�܊)��% �& �% m& �� )�	� �� ��ڮ. � )ϝ �L%��& �& ���L�܊��8����% �& �% m& �� )�	� �� ��ڮ. � )� �L%ݭ& i�& �1��L�܊���% �� ���% ��0�� �% ��0�% � )m% �% �& �% m& �� )�	� �� ��ڮ. � )?� �L%ݭ& i�& ���L�ܩ ���� �� �0��0�% i�& �% � )�	� �� ��ڮ. � )?� �L%ݭ% i�% �& ��L�ܩ���� ��#�0��3�% i�& �% � )�	� �� ��ڮ. � )ϝ �L%ݭ% i�% �& ��L�܎ �% �% � �i�@���% �% ���L%ݮ% � )�	� �� ��ڮ. � )� �L%ݭ% i�% �@��L�܎ ��% � �i�4���% �% ���L%ݮ% � )�	� �� ��ڮ. � )�� �L%ݭ% i�% �4��L�܎ �% �% � �i�@���% i�% ���L%ݮ% � )�	� �� ��ڮ. � )?� �L%ݭ% i�% �@��L�܎ ��% � �i�=���% i�% ���L%ݮ% � )�	� �� ��ڮ. � )ϝ �L%ݭ% i�% �=��L�܎ � �% � �
i�@��L%ݮ% � )�	� �� ��ڮ. � )?� �L%ݭ% i�% �@��L�܎ ��% � �
i�=��L%ݮ% � )�	� �� ��ڮ. � )ϝ �L%ݭ% i�% �=��L�܎ ��% � �
i�4��L%ݮ% � )�	� �� ��ڮ. � )� �L%ݭ% i�% �4��L�܎ ��% � �
i�1��L%ݮ% � )�	� �� ��ڮ. � )�� �L%ݭ% i�% �1�ͭ/ �$ �. � �L����L����L��Lؠ �0 �0 )?�� )���@�	��	� �� � )���@��	� � z�h`H�Z� H�. �@��8�@����/ � �L����L����L����LC���Ly��	�L����L����L���LP���L����L����L����L��L�ߊ)��% � �& �% m& �� �& ȭ& ���L�ߊ��8����% �& � �% m& �� �& i�& ��1��L�ߊ���% �� ���% ��0�� �% ��0�% � )m% �% �& � �% m& �� �& i�& ����L�ߩ ���� �� �0��0�% i�& � �% ���% i�% ��& ��L�ߩ���� ��#�0��3�% i�& � �% ���% i�% ��& ��L�ߎ �% �% � �i�@���% �% ���L�߭% � �� i��@��L�ߎ ��% � �i�4���% �% ���L�߭% � �� i��4��L�ߎ �% �% � �i�@���% i�% ���L�߭% � �� i��@��L�ߎ ��% � �i�=���% i�% ���L�߭% � �� i��=��L�ߩ �� ��� �*�� �?�� L�ߩ�� ��� �)�� �<�� L�ߩ�� ��� �&�� �3�� L�ߩ�� ��� �%�� �0�� �� �� �  ������ ���h� z�h`Hک%� �  �Ң ���� <��h`Hڜ � � � � ��� ������h`�  �� ��`Hک3� � � ����  7�����6� ʽ �  7�� ��7� � � �  7�� �� ��  ��� ��  ��� ��  ��!� ��  ���h`H�Z�(� �� �$�	 �p�
 ��  ��0� �� ����  7���(��1� �(� ����  7���2��2� �2� ����  7���<��� �<� ����  7������� �� � ��� � ��z�h`H�Z�� 
��k�� �k�� �� ����� �� � �� ����� �Ȁ�(ȱ���� �Ȁ�2ȱ���� �Ȁ�<ȱ���� �Ȁ�z�h`H�Z�� �����ʽ � �$ � � �%��L���L4� � �L�i���� LK� � �L�i��� 8�� LK�� �L�i��� LK��� �Di����� i� � � ���
� �&����� � �J��2��2� � ������LI�$ ���| �5�  H�� �  7� ���� �ʀ� 	� L���|  H�ڊ�ȹ � ����Ȁ���(�+� �� ə��� � ��  �데 LI�� ��  �덯 LI�� � �� ɘ�(���� � ��  �데 LI㜯 � ��  �데 LI�� ��  �덯 � ��  �덯 � � �� �$ �$ � � �)�� � � �4�  �� �� ���� ��� � �� ����(� ����� z�h`H�Z�� ��
 ��	 �� � ��� � � ��� �� i �� ��� �� �����ѩ� � � ��� �� i ��2 ��� ��z�h`H�Z 6����� ��� L������ � ��� L������ ���� L������ ���� L���� ,� ȭ � �	�  ?� ��z�h`Hڜ � �(�	 ���
 ��  �� �� �� ��	 ��
  ��� �4� �	�	  ���  ��� �h�  ���  ��� ��� ��	  ���	 � �0�
 �� �8�  ��� �"�  �� �� �� � �
  ��h�  ��� ��  ���  �� �A� �� ��  ��"� �4�  ��� �h�  ��� ���  ��B� �� �4�  ��� �h�  �� ������  Z���/���h`H c�� ��� �! ��� �� � ��� �-� � ��� �<� � ��� �K� � ��� �Z� � ��� �i� � ��� �x� �  ��� �"� �%�  �윩  �ɿ�= �ﭩ ���"� �� �%�  �윩 �ة"� � i� �%�  ��� LW����L^����L�� �ﭩ � ��"� �x� �%�  ���� ���"� � 8�� �%�  ��Ω LW���LW�h`HZ�� 
����� ȹ��� ��� ��/��zh` � ��`HZ� � ��8�Ȁ����� � ��8�������JJ� zh`H�� �#�  �h`Hڜ � � )��@� ��C� ��|  H� � � �� H� � �D�  �h� �h`H�Z� � � ������ )������/��� L��� � � �/��� L�� ������ )�� ��4��0��,��(� � ������ )�� �� �����
� )�L�� ��4��0��,��(� � ������ )�� �� �����
� )�L�� 8�� ������ )�� 8�� �����
� )�L�� i� ������ )�� i� ������ )�L��z�h`���(�	��� �����#��$��,��(��/����� �`H�Z � ���2��$ ��$ �L
���$ ���8�� �����L
� � � L�����2�,�$ ��$ �L
���$ ���i� �����L
� � � L�����4��$ ��$ �L
���$ i�$ ��� �����L
� � � L�����4��$ ��$ �L
���$ i�$ ��� �����L
� � � L�����L�� � � � )�� � �D� ��|  H� �L��� ��  Z� J�L��8� ����L�� 8� �� )�L�� m J��{��w��s�"�o��� ��d��`���� ��S��O�� � �G� 	� � H�  Z�hHm J�� �  Z� � � �@� �  � h�  J� �� � L
����L����2 ȭ � �� � H ��h�  J�L
� H� �  Z�h�  J�z�h`Hک� ��� �% ��2 ������ ��� ��
 ��	 ��  �� H� � �C� �  �h� �h`xH�Z� )�g���) �" �"  ��" �`�"�" �! �!  ��! �`��! �  �   ��  �� �� �   ��� �� �!  ��!� �� �"  ��(z�hX`�# )�
��m# )��# ����# )�i	�# �# `�Z�0���� ���� ��z�`�  ���� ,� � � � ,�`H�  ����h`�Z�� �  ���� O� ����z�`H�* �  ����* �/��h`H�Z� �@� � � � ����� ���z�h`H�Z
����' ���( � �'�$��a��b��c�8�7�  ��Ȁ�(z�h`H�Z�)�JJJJ�  ��)�  ��(z�h`xH�Z� �a��$��b��%��c��&��d��'����� ���� ��$ � �a�� ��� � �-) �� Ȳ-) �� ��$ ��� � z�hX`H�Z c�� �� �	� ��� � �  ���� i � �� ��ީ� �g� �%�  ��� � ��  ���  ���  �쩇� �� � ��&� ��� ��  �� �� �� �� ��&� �� ��  �쮦 � ��i���& ���/ ��. �
�� �  ����L� �$�B�. ��L��. �. � ڬ Z�. � �/ � �$�  ��� � � �. z� �� ���%�L��. �"���� � �& i7�� �& � ڬ Z�. � �/ �  �� �. z� �� L����8 �� �
�i� �&�  �쭄 i�� L�8�� �&�  ��΄ L����8 �� ��8�� �&�  �쭄 8��� L�� � �&�  ��� L����J �� �� i`� � � �&�  �쭄 i�� L�8� � � � �&�  �쭄 8��� L����I �� �n��� � � �&�  �쭄 8��� L�i � � � �&�  �쭄 i�� L����L�$�& �� z�h`� � �$�  ��`H�� �	 ��
 � �  -�h`H�� �	 ��
 � �  -�h`H�� �	 ��
 � �  -�h`H�Z� 
��_�� �_�� � � �� m � � i � ��� m � � i �  &� � ڱ� � ���1�
���Q���	 �����
 �%� i0� � i � � m � � i � ��z�h`H�Z &� � �� � ����U� ������ ���� � � � ���	 ����
 �� i0� � i � ��z�h`Hڮ �a�m � ��i � �h`� �1 �2 �3  �� ��� � � � � � � � �* �v �~ � ���w �� `�2 ���%�Z � ���S � �T �  ��Z �Z �U � ��3 ���%�g � ���` � �a �  x��g �g �b � (�1 ���X�2 ����> � ���7 � �8 �  I��3 ����L � ���E � �F �  ���> �> �9 � C��L �L �G � �� ��� �� k�`�4 �5�7 ȱ5�8 ȱ5�9 ȱ5�: ȱ5�; )
��@��< �@��= �; )0�A ȱ5����w Ȍ4 �> �? �9 � �L'�@  �� ��5 � ��@ ��Ȍ@ �4 ���P �Q�S ȱQ�T ȱQ�U ȱQ�V ȱQ�W )
��@��X �@��Y �W )0�\ ȱQ����w ȌP �Z �[ �U � �� �2 � �| )�����3 �]  (�`�] �^�` ȱ^�a ȱ^�b ȱ^�c ȱ^�d )
��@��e �@��f �d )0�i ȱ^����w Ȍ] �g �h �b � Ы� �3 � �| )��@К���2 �P  �򀍬B �C�E ȱC�F ȱC�G ȱC�H ȱC�I )
��@��J �@��K �I )0�O ȱC����w ȌB �L �M �G � Ъ�N  +�� ��C � ��N ��ȌN �B ���y 
����z ���{ �z�5 ȱz�6 `�y 
����z ���{ �z�C ȱz�D `H�Z�: )?	@�j �: I��-j �j �? �<��; )@��J��j �j �A �8��A ��; )0�A Ȍ? �<����? �; �? �j � z�h`H�Z�H )?	@�j �H I��-j �j �M �J��I )@��J��j �j �O �8��O ��I )0�O ȌM �J����M �I �M �j � z�h`H�Z�V )?	@�j �V I��-j �j �[ �X��W )@��J��j �j �\ �8��\ ��W )0�\ Ȍ[ �X����[ �W �[ �j � z�h`H�Z�c )?	@�j �c I��-j �j �h �e��d )@��J��j �j �i �8��i ��d )0�i Ȍh �e����h �d �h �j � z�h`� `� `H�Z�w ���%�x ���w �~ �x )?
����� ���� �  "�z�h`�~ �* �v `� ���r ȱ��l ȱ��m ȱ��s )
��@��o �@��p �s )0�t Ȍ �n �q �r � ��� `H�Z�~ ���L��l �u �r I�u )��u �q �o��s )@��J��u �u �t �8��t ��s )0�t Ȍq �o����q �s �q �r )�j �x )����
�@����j �j �u �( �j �v ��* �v �n �n �m � "�z�h`H�Z�  ��  +��4 �B ��@ �N  C� �� I� �� �����1 z�h`H�Z�2 � �
�3 � ��} �| )?�} �Q�� �K�} 
��$��Q �2��^ �$��R �2��_ �P �] � �2 �3 �| )�����3  (�| ���2  �� ��z�h`H�Z���|  H�z�h`CHOOSEaAaGAME$MINEaDETECTOR$FORTUNEaFOUR$CATERPILLAR$HOPPER$CHOOSEaMELODY$MELODY$PAUSE$RESTART$CONTINUE$END$a$WONDERFUL$aaGOOD$aCORRECT$YOURaNAME$CONGRATULATIONS$BYE$PROGRAMMEDaBY$FRANKaGU$SC$HISC$LEVEL$CROSS$PLUS$FIREPLACE$UPaARROW$PYRAMID$DIAMOND$SOLITAIRE$CHOOSEaLEVEL$YOUaWIN$YOUaLOSE$ANOTHERaGAME$INVALIDaLEAP$MINEaNUMBER$�������������!�)�2�6�8�B�I�R�\�l�p�~���������� � � ����������������������� �� �0�@�P� �� �0�@�P�`�p�������0�@����� �                    @��(�8�H�X�                    p�����������Ї��                �� ����                       � �@�����   � �                (08@HPX`hpx���3�;�C��ޑڒ֓ҔΕʖƗ������	18?FY`gn����"	}��������)�\�����$H|��c���d�
K�� 9ڲh�!��~�P�X��^_`abcdefg�����������L{���&_����9h����qrstuvwxy?Qcu���������dh�b�~���X��(:L^p�����1CUgy����ӄ����� ��^M�p{,�~�YmX��9_����"Df�������������^����IJKLMNOQRSTUVWX���������������t���!ڇ�:C�������v��%&'()901234 D����˷���������:D������Ȼ����cd��7<JKLM BFh�������۝��� �R����K�k��L�8\����)Mq���>b���/Sw��� Dh�����
	,<L\l|
�;�l�������0�                                                                                                                                                                                                                                     0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^_____  0@P`p��������  0@P`p��������  0@P`p���������������������������������������� ��@�����J�f�r�v�z�V�n�t�x�~� � ��� �p�� � ���Д �p������������� �`��� ���   �`��� �����@�   �`���   �          �  �   �

		�
 �
�  �                                                   Z� �s�