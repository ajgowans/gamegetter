�P�А ��� �@���                ��������������������������������d���j���"���*�����������i�f�Q� �������U�������������������������j���U�U�U�e���j�������������������������������(� � �� �� � ���U PE  T  PD�f�*&����������� ` � b�� ���ha��@� P � @ � @    ������UU��������Z��������������� � � � � � � � ��f������ff�Uie��"��**������j�������! � � 	��@@@ T @     A        @@@P@U U TEDDD�U���Y�f���jj����jj����  ���ii�fUYUU@UUT                   @@PQT ��f�j����������� )�fd� ��Y�ff     DA   @ @ @@P P@UAFUJT*�E*��d������j���� @���ffYUU PUUU                  ��U���VU��U� T  �U���Zjif�fei�Z�       TP@UTU        A       @@D Q@   D            @DAQUVEYQfUZ�Y�V�f��  jUUEUUA U       �eh�VeU�Y�ffYYfV!�@� � ��� ���     U"A(A� @@AUUETQAD        @@           A @ @ PP    QQDUUAUPUUU@UUUUU  UUU              T  T @  �$AQ���Y"�����           @ UPDUDUDDUTUQT               @                  A @  AP  @ @ @UU  Q     UU T                 ��XUXUXUXUXUXU����`f���f � f � � P  @PUT�QUPUUU@UTEUPTTU U  U Q  TP      ��FDFDHDHD`� �a� �`d !`d !eH%`H `F `F �D��D��D(h�"!fH��� ( ��� ��� � � � �f�	f
�)f&����UU  �����ViY�VUUTA@UT U T   P  P  �B����J�"�f�"���������F��F��F��F��F��F��F��F��F��F��J�"����F�������
�*���Z��           � h�h�h�ZhUVUUUUUUU                           @     @ ��DDDDDDDDFDFDHDHDdD!dD!�D��D�DFDFDHDHHd���  �*����"�
*      � h�hATAUTUZUUUUUUUUUUUUU        �     @ �`$@  �"U� ���              	A a d a$!$!T$EaU$ a$ ! $ ! $ !  	  	        
 "         X XV       U U U U  U                        EPUP   P                         @QQTDEUUUU  UQ��QT����QU      UUU�U�ej��ef����A �!
��jVZV�UUU@PQ @T     @E        P       @@@                   A   @             U P        �  �������	 ��@e P      U@UPAU UUUQT@TU  TT  UT           APT@@@  QPEUUPEUPT@   P     @ @T   A                    Q  P             ��
  �`          @PATP@UUPET@      A@AP@PAAAA@E��B����D� A    *j��jf�UUUUUU���                AP          @P@@ UU �  � � � ���*Z�U������Df        PUE AUU PA                f��jUUUUUEPDTi@� T P T   @  �h���R�Jh�J�Jj��
�(j��!����f���  �* � * � ��T�T      " �  Q  @  T      UQU       U UE         U E T P D     U*����PU@      UUUUUP EPUUUUUUUUTUT��������U��T� ���������PU @    ��������������*� � � � � � � � �P ETAU@TTP@PU A   P P PPQUTQQUU       @UDTUQETUUEUU�Y���fQUTUUUUEETUVU���j������������UUVUfU�Uj�Z��������fY�*(*�����UZ & 
 � *F��"*�����f$�	j��)��j�"���B���V�����*����*�������j�������������jUU          AEU AUTEUTQUUEUU   DTDAETQ  UDDDD@ @ UEEUUEUUQTUUUDQDUQUUQQUUUUTUUU    �Z��U%�&����*�������      D������� � ( *�
�� ���������j������*         ����*�������UUUUF ���f��V�UP UTQUUQUUUU�U�ZU�  * � �
�U�              ��&�j�����@    �j������"������@DQADTQUUEQUUU   D DUDTUU  * �  � *�(���������&��                � � � � � ���            �Ad       j��� �ai���j����UUTU  ` Af�jUU @PATP@UUP � @   `@ �@���   @ U       UU     @  @        @ @DUU            QE   @                  A A              @ @@@ P           @    P  P@        @          P                 d���U�@U@  T QEA A  PU              P  @                                    ATEUTEAQQQ  QADAAEQEATQP@@ TP AQT Q@PP @@     @@       TA    E       @  @     P           � � � ��T�E�U�D@ATQEE��             �E�U��T�U�D���@ @     D QU     @ DDTQQUU    E  f���&�������E  EA               P   E    P   UP    @   P@  @          @              @  ��X���i���������               @     P D E  D    @  E    DQDPEUQUUUU TDDQEEUUUe�(��� � � � � @ � � � ��� * �     � � �   � ���*�
�*��"�
*Z�������j�������                                           A            T @@UQ@@@T     @                D��D��D��D�U�DDDDDDDDUUDDDDTDUUUUUUDDDDEUUUUUUU@DD@P@ DDDDDD TDDDDUDQ   D��D�Q�� � � � � � � � � ��Q�           TUEDTU      PDDDDDQDQ P�
�B@UU    ����@UUUQ    JD �D"�j   ` `��* ��""��DD     � � � � � � � ���f������iY��jff��ff��if�YY�e��efZ�e��YeeVU��UUYQ�eUQQYUQQUQETTDEAUQPTD     � � """(��f&f�i  Fe������j&���F�������j���f�������Y���f���f���i���Y�e���f�����Y�e�U���U�Q�e�Q�Q���Q���E�T�E�U���P����� �� � �DDDDDDDDQQ  E      D��D��D��D���Q� �� � �� � T   @               @    P  P  P                  @    @@   DU@      TDD             @  @ QDDE   T D P EAQ@@DQTDDDDD @ D U EAEDEDDDDD           @  ����UUU               P @      @TDU   @ P P@E        TT                 T  P   @P D T  @ AQDDDDDDDT             @ @AE@EUD   P  @EUjVjV���ij�����j�      @P     DDTDDD           @   @   U DA � �@�� �@�P��D��D��Q�@� � �       A P P      A D DDDQEQDDDD @@  PDDEDQEEQDDDDE Q@DUDD EETEDDDADDQDDDDQETDDDDDDDQEQDEDDEQPQDEDDDDDTDDDDDDPE PQ@DEPDEQDDDDDEDDDDD    @ @ADEUTDDDDEDTADAPUDEQD@QDUQDDDDDDPD@QTUADTDDDDDTDTEEPDTE  QED  DAQ@EQDDDDDDDDQP DQDDDDQ@    QQDDDD ������D��DDDD��a �U�Q� UQUTU    D�� ��� ��@D      DD TD@ A      EU            �D��@� � � � � � � � � � � � �                 FD  DD  DD  FD  DU@           DDPP         DD  DU@     DT D D T               � b�X	��j�Z�Z  DDPT @        DD  DD D    DD  DDU  E  P PE  @          DD  DD DE @ bD	 FD  FD	 IDDDDDUUTQEUQDDDDUUQUUTUU      PETDDD        DQDD              QDTDDUUTEEUU PDDDUUUDDQUU     TAUUPQUUU        UUPQEEUUPP   UUTUUUU@  @    UUQUEQ� � � �U�U�E��UEQUQUQTDQQEDDD@@U�E��Q��Q��D��Q�E��D���@�        @  �� � � �� �@��
Xe���������TPD PT���������������i��iUU  DD  DD  DD  D�  D� �D�  D�  D� ��bUUDD  UU��  DD  DD  �DVIA	IAIA	AA	AA	IA I@ QF� HD      
�%H�$a$��$�$X$��@ �P��@$�$�Ud�d�dQZ�ZDj �D�  DD  DD( � � R � $ % 
   hD� R�����RJB�Q"�  � �U�U�UiU �DV�UdE`dXX
 eD� TFUPFT	PIXXEXUXU��XU����U	TIU	UI�
UI�
�J��@DQATU����  @DEDQ��� 
*(���
����� " � 
�*������U�UUVUhU��    ��j�U%U	�*         ��	"%����  �" ��&`���F  DD  DD  DD  DD% eD& JD  DD  DD @               P                DD �Dd HDF�E�E  DD HD  �F ( � FDH `D�  DD �D
   TTZ� *J���� �$ ��Dh �Dh� `&��&&��b�`� �Dd �D�  D� `D`�A�        ��  �D���d�X�X��  ��
`�Z�DDV)VJ� DD  DD  DD  UD@ P @ @     �D� �D� �D� �D�jVjV���ij�����j�  DD �D$ DR�
  DD HD  �D� UFDU�U����� eD	 �F* h�"���&��Xb�$�@@�� b

�D& �D& ID @@@�@� % e � �                 � � � �
�*������� �� �� � ��D��D��D��D�U�U�Q�U�U�E�U�D�        DEQDDD@DDUUUUQUUUUUEUUDD�
�
U*P)               
 *��*�
��VjUUU        P� � ��j�VP      
 � ���������������� � � � �@� � � � � � � � � � �*�����Q�D�� ��U�U�Q�T�@� �  @    @ TDP@ @ T@ DPPD@U E  D  P   @@      T UUU   @PU PUUDEUQU@TT @ UUUU@UU        UUU            P   Q  P @  D��� � � ���  @            @ @    @ @ @      @    @@@@@   P @@DEQDAUU @U@UDUUPUE   @ U      T              @  U @@UPDUU     @           @� ��� � � � �      TPPPD  @ @@       T ETP     T@@@@E@Q@  @A   U UU UU@@ TU@ E@U   @ A @UU          TU  UUTUP@         U                      TEU@  @  D D UP      UU    @    UU   @@     D@ P    @U   UAUQ  @T UUT  U  UT@U               PDP@@ @@ @           U  @PZ�������j�������@D    @      A@ E  @             UU        PTAAT@QPU           @QU T        E   DU  A                          U@E@AD  DUU  PQ               � j�UV@                    � h   F�VF@ @ @       UEP        T DTPUDUTTPUU          QUE P U@                   @      @ T DTUTTUUTAT U   @Q  �Ua�E�e     ��VVAU @P  Q       @          A                   P @ @   @U T@P EU �d@e `  P�
e�P @D PV�d PYD P D Q D PTA V@     @ ` jU@                  T @U         � X �     ��UVD V D @  @         @TEDA   P UQUT     �T� dQT   � V�UD P             ��UU              �U) � P     @          �	T$�@     ��UV F A @            UT�@a�`@� V�U A@PV UD Q A  @   @   @                �*Z�EAT@A                 ���������������� � ��Q�T�Q�� �   @DPEDTA     @  P        @ Q @@ @        @@      @                         T  @       @      @ UP@AUUV��YiAAP  @A @TEAPQAP   EEUUUTUQ@ PP PTU@P  A @@QTEADD@ � � � � � � � �     P @ PAD  PUP@     Q DTAPE@ @ @@TQA@@@@@@@AQ Q  @@@@TUU@T U   TTT@PPUQAEQAA@EQDP     DE P   A DDPD  @T D U DQD @@A  TE   P  PE@        UE  DT  Q@@DQTPP@QUETD P T  PAPQQTPTDQ@@  @D@@PPQUUEEAPPTDUUTEPDPD@PD@UAQUTPDUPETEEDDEQQDUEQPTQADDD@D  PPPPAETDPT D D D T UUDDT @ P @ DEEPDUP   PAPP       A           AT@ EQUUUUUUETTA@TDUUEU@TAUEQUE   P QUTUEDDTUTPTATTUTPUQQQUUEUUUUUDTDUUDUQUAEEDUDQTTQDPEQEEEQTQDUEEUTUUDDQDUAQPDQAUEQ Q@AU@PAPUUAUQPE A@@T@@UUUAQPUEP @@U@UQUAA DUU@P T PA   ATTDTP          TEPQTUUTUUTUUTAU@TADPTAAA P     @ � � � � � �P�E�P�E�Q�A�U�U�U� �U� �D�Q����� �@� � ��D� � �     ATA      PDDTQ@        @UU@ D @ @ @ @DDPUTUQE@EEPA@ P@P@A       TPDU  E@@@E@Q@TPE P@    AP  QPT    T      fY���Z�f������fZUU�jj��Z��������T UTUE  *(��Z��j�Z������j���@ E@   	 � U�jU�Y�f�i��      �
�)U��������f��f���Z�����  
 �f	f%�&�&�%V��eV��j����i��� ) % � � � � �f���V�i�������i�jf	�	�
Z*Z)i%�&���j������������i���i���f��������Zf���j��j��jf�U�e�fZ�Y�j�j�f�Y�PUEEQDE   U TUTTPU   @   PD          D @      PPPPTTT     @ P D DU@TTTTTTTQUPDDD@   A @ @ ED@D QQDD T PD        AD  P@U @@  QP  UUUUTUUUUUDDEUUUUUUUDDTUDD@D    QDDDD @  TUUTQUQPU T Z�������j�������     D T     @ D@   UUUEDDATDAT UUUUUUUDDQDTUU@UTUD                �*"�*���*�*��������������������UUUUUUDDTU�	�b�*���
 @TQ   �
�*���"�*��""��������������"��B�
�B�
(� T��T�� �T��T� �U����������� �������i�����U�@�P�A�T�Q�$�h���h�T@UT@   TDTA@@PPDUP   DU PU TPAAT@@PAPDDP EQ PTU@@ � � � � � � � �U U
 ��"���*�� @ Q    *������������jf��ff��f���fj���f��ff��ff��ff��ff��f��)����f&�J�PDUPf
�IfJ�&DIEJERUUUU@UUUAUUU @  @   " �   UD          ����ff���f��f�������ff���
jP@TU&@Jj����U TUUU@UQTVUZUPQUUUUUUUUTU�E	V�TEQUUUPUUPUUUUEQED      @ T           T@     ��Z
RUEUUUPUU  UUPUUPUUUUUUUUUUUPUUU@TUU@TUUUUTUUUUTUUUUU�U�Tj���f�  EVUYTJ
UJD        @@���         P *@��UUUUPUUUU@UU��UUAUZ�jPUUUUEPUUUU PUUUUUUUU@�U�U UUUU UUUU@U�Q�E�TAUAUUZU�T*T@TPDD         P �P �� "�
"��*���
����UUT� h���aY��������Y�Z���j��� UUZUQUU@UUPUU  UUAUUUTUU UUUU QUUUTTQD@PUUeT��D�D   P P  ! � �
P@            ��ZU�TZRf)��U��
  U��UP@U*T@U PUUUUUUTUUUU�UUU @UUUUAUU@UU�Zi
�JZ)�
�P  PQUTU UUUTUP    @ P        @U        �� 
* ���*@UUTUUPU��UU UUUUUU PUUPUUUUUUUUUU� UUAUUUUUUj�V*UUPU�Z�ja���� @AUUEUUABUTED E  P     �   T@  ��������jP�UTUEUUP��ff���f��f��hfUUUUUUUUTUU���f���UUUUUUUPUUUU�U��Q��UUTUUVU�����
D@@� �����P�� � � � � ����j�����f���f��ff����������f���f���ff��ff���U@U��f���f���f�����UUAU�UUUJ�@h�j�������j���f���DTQQDDAEQTQEEAQDATADQDEEADDDDTEEQADEEDQQPQQEADAQEDEADDDQTTDDUEQQETDQAQAQDQDDD@DDEDEDEEEDUDQQDDDQQDQEEQDQEQEAAEEE@ EAAD       DQA   DA DE�Q������Q���A���A�Q�E����������A��D�Q���T����Q�Q�Q�D�@��������Q�E����A�A�E�E��E�A�A���D���A����D�U�D�@PD P@TQPDPPEDAPPATQQUPP@                 TQP U           A@UPT   QP@    � ��U�Z�f�e�e�   @�T�VV�VUVT  � � � � � � � �UUUU�U�VV�VURUT @UUZUbU P   T P�P�VR�VV                           @ P T      T
UfT!       � ��BVPB  PTTTP@@ UUUUUUUUUUUU     Z &Ue    � � � � � � � �   ��YU*����     @��iU(�UV��Df���f��@��% ��DDU��� j �U*��Z�Z�Z�Z�Z�Z�Z�Z%%U%%%%%%�Z�����
(      �*
*   � h�h �Z�Z���*� 
  � h�hQ P  %* 
  � h�Vh P  @   @   P    U Z�U�j��@PEPT@ P  Uj P��VP          �U��U� U         �����V�P      j��Z����@�@U P             TU     PP @U   UAUUUUUZUfe % %%U%%%%%%��Z�Z�����   �%
* 
  � h�hUU h�h UUPUUPQ U @PUEUUUUUUTTUUAUP@@@UUUUUUU U      PP   TU     P @  @U �j���jUU   P  PU����AU     UUUUUUUUUUUUUU%U%%%%%%%�Z�Z�Z�����

   %U%%*�         ��UV  PUUU��UUPUEP@@PQEUUQUU UU@ UUUUUPUEQPUUUUQQUU E T          UUUU UUPU            @  U P  @ T    UU�����UU        �Zj�UU P @  U  �Z�Z�Z�Z�Z�Z�Z�ZUU�U�VV�VUVV  �Z�Z�Z���      %U%%%*(* �  ��UUU TP   � U* �T@     TPUUUUU UUAUUU T UUEPUUUUUUUUUUPUU UPU TU U ��V�RP TUPPU  QT @            U UUPUU @       U�UjP� U @ UU   ����jUU      �Z�Z�Z�Z�Z�Z�Z�ZUUUUUUZUfUdU T   � �   ) �@) �%*U*  ( �    @  UTUUUTUUU) �@)U�DAU   UU UUP  U@UUU@PUUQUUTUU@UUUUUUUUUU U    UUU@UPU      ����UU @        Pj���UU@ T�Z�Z�Z�Z�Z�Z�Z�jUUUU�U��VUVUVURUUUUUUZUfUeU!   &U** 
 �     @UUPUUUUEUUU@) �Q)�UA      @ @        U    U P        �V����UU        UZ���VU                  %%U%%%%%�%*�Z�Z�Z�Z�Z�Z�� �%%U%%%%%& �     ) �@) �*U*  ( �      @     TPDU) �@) � UT�����Aj����U� U @    e����ZjEUT  @�Z�Z�Z�Z�� � �   PUE AUU PA       * ���UZ � � � ���V�U�P�VUETUUQ    U��E�U� � � � � � � ���i�(�U���D��U����j���*�%�%�%�%�%�%�%�%�%�%�%�%�%�*�*�*�    � ��V E        J&!@                  UUUUUU         @ @     @UTUUUUUUUUUTU     PTUTUPPPUPUPUPUPUPUPUTUUUUUUUUUUUUUUUUU           U U      U U                                                                                                                                               8<HIR       chi:=JKST	)*7dejk?ALMUV+,9ofglmCENOWX -.;npqrsFGPQYZ_>!"/0  
  [\   @#$12  tu ` ]^   B%&34tu       ab D'(56                                                                                                C#               %&      1 4  ')       2358:<*+   ,-0"!  >=.>=>=>=>=>=>=>A?@67?@?@?@?@?@?@?B;;;;;;;;;;;;;;;;;IDDDDDDDDDDDDDDDD9/EEEEEEEEEEEE
	$FFFFFFFFFFFFF(KHHHHHHHHHHHHHHHHHJ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������t�4�d�Ę����ԫ�$�                EE       @@TA UDP       @  @@UUT QQA   P  @@@A   AP        @ @    @   @               @       A @       � �@��E� �@� �           @         @     @P @A      �@���E�U�Q��   @Q@Q@DTE     P PF� � � � � � � � �      �                           "     ( �                 � (        P P                � � ��� ��� � �� � �@�@� � �� � �� � � ���   � "�     ��(       ���*����	 (	  ��(( �     � � � ��� �)X� �   ��U�
(" ��VUVUVUVUVUVUVUVU% ��eY��" ��eYUYVUVUVUUUUUVUVUVUeY��" ��eYUYUYeYVUUUUUUUUUjU�j ���" ��eYUYeY��*        � `*`��Q��        ��UV  * � ( � � �    @P  (�� (� 
(�  ��     � � � � � ���� `(X�V  
 ��U	U� � `UZeVeX�b�XUVUUU% %P		 	  R VUXUbUXUVUUUUUVUT    Yi	�XUbUXUVUU�V��
 	 ) � 
  � �       � � ��%U$�   
                    
 X (PT       �  ��P U   DH" T   V B���U  HT            ��V( @UU@   UU   UU �` XXff���� @ @`U H H XU���U`U`�`���(@@ @ @UU   UU @���V�� � XU XUUEU�( " � �        @ @ UUPUXTTQUETTAD PP  ED@QU   D     Z�@ UU UE   � �UU  UU   UU   UU   UU  @ @UU�� � UVAB��U� TUA@��������h�� �UU@P@������hf����TPU@ A  @    P  @            
 �  U	 � UU   UU  BP      % � 
%�U� j)V&B��@� � UV B)f)V&)�ZU`  DUPQUQ    @ P   D     @   @  E   P       @    T        P   U PUXUT���  E    UUU���*       @@E          D Q T    @      � V@U � �     UUj	�      @@@ UPU     @ @ PPD TDUUE  UUUU TTTUUQUUEPUU  UUUUUDUP @  UUUU@���� � � ��@@UUUU@ @ UU�U�T��U��D�U�UU@ @ UUEP@��U����P� �TD@       QTDU  @@U @   Q @  P ADPU    @P@T @  QD @ �U��E��U�� �     @ U@U �        U UjU�                            @    A               D             P@     ��"�������������EAU@ �d�����������������U�U�������������DUU���*������� UUT�"��Qf��  QUT   DTTU T   "��*�
(*�� *��"����������  UUUUEETTU T  UUUUUUUUTUT aUUUUUUUTUUUT � � � � � � � ��DUUVUQUTUUUTTUU������f��fU�YU UD���U��YUVU���� @  @ @ @ @ @ D   P  PPPT E@PDDDDD             @            T@EDDEDDDDD   @ TPEDDD           @ P PDDDDDDDDDDDDDDDD��D��D��D��   @ UUDDDD        UUDD  EA D ����U�U�UUjV��E D  E  @             P   PP     E E��� ��D�P�U�      @  QU  T DTDD            Q DDDDDDD      DDDDD�UV�ZUeU��j�V� ����
�*��� � � � � � ��Q�   @   TDDDDDDD @EQDDQDD  @ @ @   @D@@QPDPDDD� ��	 ��YU��
��� V�j `��Ue�����   @Q@D@ADQ" �""����������  @QDQDD��U�jjUUeeEUUT P@Q@DEDDDEQUDUQEUUEUUEU�DDDDUUU�U�U�V�Y�f���������j��UUV��Y�Z�i������D��D�Q�U�E�U�U�U�V�������������ET @@A   EAU@ DAT@TPTTQET   ETQT  DPQUTUA@��������h�D ATUT   PU��U�j�U�e��U�T�D��T�U�T� � ��T� � ��T�� � �                �� ��@��@� �E��U�D�Q��Q�D�Q�D�U�D�Q��E�T�Q�U��U�Q�U��T�U�U�f�U�U�V�T��j�������������������������������V�Y�Z�Y���������U�U��f��j���f�������i���j�����U����f��f����VZUUU��������U�����������h���UY�������Y���&���������didi�������j� � � � � � � �@� � � � � � � � �                            @dF��������*����� D�eh�a�����������*����Y����������*���Ye�����������j�������j��VZe��eiY��UYeeYVjj���������j���fUUU�fUUUUUVETUU��ff������fj��ifQQUUUQQUUEUTT���e���fe��ef���QEDUUDQQUETU           U	Y	U	@"j�V  F�F���b������ @���j��j�����(�����UU������*j�Z�"��UV������EQUDQQQDD              A @@ @  VUVUZUZU�����j��U�U�U�V�U�U�U������j��jj���jV�VUUUUUUUUUUUUUUUUU @ � � � ��� * �ZUUUZi�� P P @ @ @       @  PP         f ���������eVYff���U�U�U�U�U�Z�U�UUj ��*f��UU������    j UU������������i���UYeeYV����������������U�U�UeU�U�U�U�U�����������������ed����U�U�U�U�U�    @@������*���� � � � % % %@%         � h�VhE    E    �     ��`DFD `   H  H  F VDDDDDDDDUU   V V  UV������  UUUU  UU���������������������������������j����������U�����U�UU����������������EUUUU�U�QUUUUTT���������jUUQETU        
 & & �               �  ��DDDDDD    * �D!D��������ZZU�U!V�V�*  �
 �       D    @
��j�V`U        �j������j��f��������eUVY��������j�V���U�VU�UZeZUjUjQ�U�V� � � � � UUU��V�V�F�U�U�QUUXU`U�ZU���UUUU��& * ��VZ�VUfV��`UXUXUXUVUVUVUXU               XUXUVUVUVUQ� i�V 	 $ ! $ � � � U��Uiej��*�
�&V%  � �   �U������        UU������     
 
 
 �ZjV�f���������� @ P @ @
P � Z�Uj��i�Z�*���j���f                 �U� �U�� � � � TU@T            UU PU  T @    UUP            UU TU     @U@      TU       @U U U @ U @ UP        P  P  @ @ @ PU@  U  T  T  P @ @ @ @ @   @U  T  P  P  UUU  U  @ @ @  UU             UU @U@    � � � � � � � �����UU  ZDeU�U�����U�T�T�T�P� ����UUUU ��Z  UUP  U  T  T  P  P  P @ @����UU  D�UYU�����U� �D�U�U�������U�U�U�U� ���j)Y�DVUDQF�&��UUff������j���fi��ff�UVi��ffZ�efU�f�������i���e�����������j�Z�f����������������"  �����*�����*���i&�	QVV  @DEDQUUEUU@ T       � � `         @  ` `   ` � �@��TEUUUQETUUTU@�Q�DaUaUdQTYU��&U��JZbf��bf�Z��E��UUUUIY�j���j��Rj�����UEUUEYUEY��    UU��UVUEUUTTQ PU � U
�% �
UQET�E�(�              � � ! ! YTHQRU       EDTUT�� D��UU @ QDU�VUh��e���U���U�@TPQDTQ T @��TU��U���U��aUb�ZV D    @
��j�V`U           � V��             � Z`
�P X UX�Ze��� `      ` ` `�
��P�@@
@*@� � ` � ����@�@�@�@ ���P@  	 �   )�@ @e��*	       T d � � @      U����j�Z�fTj@� �i�Z��jYe� � � $�V���U�U��VU@VP  UUUUUUUUZU      UUUDUUUUU�        ��UU�j �          
 % � UU @ @UU�� P P�i�TE	U	j	e�jV***�%�$B�I	�U���jfe ii!i%Z%*�"�*�*j%Z%Z Z ZZ%V%			@	�VX�Zh��
���*�@*��%  @�Vi���
 ��	��j	Zh ���j V  U@UUU�����Z�V����ZU�jjUV�U����j��P�      UUTUUUUU�� P   UUUUUUUUU�U@T@                       
 % $ � � � � � � � � $ $ $ $ $ $ %��h�i        @ T@UT�U������V�j��j�UUUUUE e UAUU��U�U�U�������������*�������U�P�@�@�P�P�T�      ��`E   ` a e �U�Tfe�UUf�������jf�f�f��U�ZffZ�ef  UU  UU  UU  UU �U� �U� �U� �U�                E��D�Q��� �D�E�U�T��D��D�� ���U�U�T�U�E�U��
�%�����U�U�D� � � � � � � � � � � � � �A�� �UDAUD@ DDEEUUUTQUDDUDT�*U�UUQUUUUUTTUUVY��e���V��jZUED 
 % � Y�
e%��           TP DDQPTPDDUEUTDUDUQEDU�UUUUQQTEUDUUUV��ee��UV��e��ZU�UUUUUUUUUUUUUU@DDPDD�@��D��P��D�UV��e���UV��UY��            � U*EQEDDUUAEDEEUUEUQTDUEE             �*�*�*��*""""��UUUUUUUUUUUUUUUUUUUEEUTTUDDTQDUUUUUUQUUUUUUUUUTQQUDUUUUDQQUUET@D  AUUUUUUUTQEUUUTT@ UUUU@ jU�*U�B UUUU@ UUUU               * �������*�*""�"U*U�UUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUEUUUUUUEUUUUEUUTTUUQUUQQDADADDD   �   X �U XUQDPEQTEQE DDUUEEQUEUUEPUUUUUUUUUUQEUUUTU 
     �������������U*U�UUUUUUUU  VU) �VU)U�UUUUUUUUUUUUUUUUUUUUUUUQUUQUUEUUQEUQEEQEED@UU@ jU�
U�UUUUU  �   X �U  XUTDPEDDAUTUUUEUEQP          � *  ��� � ( * �PU
U�UUUUUUUUUUUUUUhUVUUUUUUUUUUUUUUUUTUUUUUUEUTTUUQUTQQDQDQT V�UXUVUUUUUUQEU   �   ��U
V X X   T @     QTUEDUQ@UUQQUDUUETQUTD              @ 
U% �U)U�UUUU             ��ZEUUUUUQUUUUUEQAEEDPQD(       � ZjUUU            ��
             UT TDUQDEQUDTDD@jUUEUUUTEUUQQU ��U)�)    ��    �`@X@X
V�UUVU)U�UUUUUUUUUUUUUUUUUUUUUUUEEUUQDTQDEAAA@E             �U� �U� �U� �U�QTEETUQTEATQTT��UUUUEUUUUQEEj��U V V�U���*�    @  @P  �
UEEQDUAQDD��UUUUTUEQUETUU	 �U)�)    *  	 % � UUU	U	UEUTQEQDTEUUUUUUUUUUUUUTUUUU  UU  UU �
(��ADE@@@ HFE@@@ ZUfQJjD!UTEPEV�X�b�`DUXJPEVEQUUTUQQZUjTJ�YYUe�UVVU�UUYUU�J�j�j����V�V�F��YYUf�YV�U�V�Z�Z	"�%� ��@� @ �"��e�V��Vee�YU���(%���!���%���UUTQEPDUTEPE��E��	�@*@ (h���h(����"")X�Z&�H V�%V�F%X�R%��
T�EPE 
�����(�
���*�
((��
���Z�TJff�������j��jj���������j��jf�������ief�VY��fe��V�ee��U��Vee�YU����
( ���"(�VEQUUTUQQTUUTE�����ijf�V���f�� � ����V�eY�f�����������j�������������j���������e���Y���e�����e�����V�e�Y���Y�e�U�V���U�U�V�Q�U�U��T�U�E�U�T�E�P��T�E��A�D����@��@�EDP E  @                      �j�j�� �
�����
��YeeeUfVe�U�UDDQD                       �   ���*����"����"�� ��         DDU T          DDDD@D  P @          ����         � *"��"���(���**�� �� �*������"��� (���"�*�� � � � ��(��   
 
 * EDDDPD@@D  
�� �*��*��� P @�@( ��"��DDDDTD@ �"           ���*"���� ��(   DDTE @      DDDDDDED             @    @�Z *@b DDDQ                 � "��      � ��� "  ����"�      DDDDQDQ   DDUT              �� "��**�������" 
 �
 * �D�� � � � � � � � � � ����"���*����� � � � � �DDDDDDDDD��D��D��D��DDQDQ       UD  @          ���"�
����  (�����ief���ff"e DDEDP E  b��DDDDDTf� ����"�� � �    �"*��* �" 
 
 
 DDDD@E  P  DDDDDDDEQP���e��U��Vee�YU               DDDD��&
�
"DD�D���������� �  ($�d���Dj�����������JDDDDDDFD��������D��DDFD�jD��j�����VQUdUa�Tj�b��D�)D$!D�DDJD�jD��J������D��D��D��������������������������������j�JD����DDDDDJD��F���*���j)D��DDDDDD������������D��d���U�@U@  T D�DDDDDDff
�����j��Rj�V�ee��U��Zej�Z����*�F�*�F�D�V�ee��U��Vee��V������"� ��(�(�(���������j���f������������
@BX� $�� I�&U�b��e������ihf�VZ��fh�                   @@ Q  b%ZI�R%ZEUUEA% 
             U�U�Y*�*�&�&�%�%UUUU� � � � UYeieieU�UUVUVUY     �*���� U
U�)�"h��U�UjUUU	X	V��Y�YV�UUU`aT�UUTUUDD VU�U�UUVVV�V�ZZ`U���� � ��%�� Zf��b X�VUUUUVUVU�XV�V	V�XUXUXU`U��jf���i*������ ��%`�X�Xb���h�� � � � � � � � �            V VBUP@VEU    ��X��
 @ `
`&j� ��` UU��""UU  ���UfDeU��""��  ����fZ�� %�%�����V��@b*��H��j"�"Q"�e�%�E��E��E��H"Y"D"Q"D"Q"D"�"����&������dU�� "�""
" "�Z ��  UU  UU  UU  UU �U� �U� �U� �U�  UU@U        D��D�� � �� �  UU  UUDP @   @U P            UU  UUD U  @ @U  P  @ @ @ PU  P  @      UU  UUP      @U U          UU UU       UU U          UU@ T @        UU  UU P @ @ TU@  U         UUPP         @U UT        TU        TU      �P� � � � � � �   XXXPYE	T XXUU@X XT	@	R
F��

��P X*�h*����YU��""�jE��fZ��U��""�j  ��U�f��BeX	J�(�*�%�!b�@b*��H���"U"E"%b!b%b!b%b!b%b*�""f""E""E""�" b*�(b"�(b��`X��@"�"�"("
"�Z����f���U�V�U�����         V B UUQDEQTTTED B " b b�� "�� D@D  A    `U��$"TiPE��hV�         ��� "��`� �`� �hf"�h�*f������ ��  �����bf(fbf(fbf*fjf(����je���U�e��i��f&*�j�&&j�Y�	Y��    X H  X X       T @ E T     ��U ��@@   ` `��f ���PUU��""U�  ���U�DVU��""Z�  ��eXh��eU����A���Ubj��&���)b*�%b!bbIbbEbbEbbE��&b"b$b!b$b!b$b*�b ��b�"b���X�� b*�"�*" �������        V BU�Q�D�Q��T�E��VBU
X%*H�
�! � � ���� � �U%�*""U  �*U&@�d���U�@U@  T ��@&*��(��jfe"a&��b�����������"�e�a�e�a&e�a�e�j�����*���������j�`�j�h�bfhb�����                       ��**    � �          �
UDU     � *    
  PT  ��
�  �@@U Q@ U                    ( � �  UUUUa���j������ T@P   U   P    P U P PD  P         @            ��f���f���f���f�a�����Z���������DEUV��ej�������� � �A�T�E�T�U��� � � � � � � � � @ P @ QTUFTU     D  EEEYEZ�jfj���j����jVVE�j���j���f��������f������������j�����������           @            @ A @EQQVUVZUf��eDUDUUUUZ%f�j���j���fe��UV��jj��f����fi�VeZ�         EP    P @T  @TVETUEbU�Yej��QATEUEFUUUU @ P DPDU DP        E  T PDPDTUUUV�Q    EDUUY����Zf���j����������j������f���j��f���ff��f������������������ff�������f��ff��ff��ff��f����f�����Qfj��f*�BPU���f��f�����j@U��fj��ff��f������jf���f���f�������fi��f��jf��f��������j��ff���f��U�
T� � �TBUUUZ� �
�*EU��ff��ff��ff��ff��jf��P�PQ T                  U             UUUUU             ADQQEUT              UUUUUUU       @UUUUUUUUUU   T UUUUUUUUUUUU  UUQDEQTTTED    DDEEUU��EDETPef����ff��ff���U U��ff��ff��ff�����TU@� h ��j � �Tj��hf��jT�Pj��ff��ff��ff��ff��`f��ff��ff���f   � ��e ��f��`f��jf��ff��ff��ff   � ��f���f��jf��ff���fE��f��ff � h �  P   ��j��ff��ff��ff��ff     � j��hf���f��hf��jf��ff��ff         ��j��ff               ���ff���f��ff��ff     @�J��ff��ff        * ����ff      �*��ff��ff           ���jf  QPTUUTQ    @ @PUUTQUUUUUTYU�ff��UTTeUiU�ef������    @ P@QUQT       @ P AATUUUTQYf�������UUUUUFQ�e��f���   EUEUT  TQETUUUUUUUEEUf��Y�����                 ��D�U���f�����      @eY�����    "  f ZDf�i��%���%���%���������������%�%�%�%  " "�� *������``U`@`U`dUijUFF		X*��` `U  � � V� VJJ         & & �  
�%`�`��*`�`�`��j%��*�%�*�%�*�%a�e�`�e�a�e�d���* � � � &"��UU`�`�`�`�b�h�`�e�������e��������� � � � � � � � �ff���f���f���f��ff��ff��ff��ff���f�Z�j�����������Z�j���j���j����ffY�ff���fi��Z��ff��ff��ff���e�����j�������fi����e���Y���j������ff�YffeYi��f����if��i���i�j���j���������������������f�����j�����ff��ef�Yf���j���f���f���e���f�Zjf���j������jj�����������ij������ef�Ye��Yi��Ui���ff��ff��Zf�Yj���i�Z���j���������������������j��������������������Z�ieZ�iff�ii���UUUUUUUUUUUUUiV�ff��ff��ff��ff��Z�V�����ff��ff��UUUUUUUUUUUV�Z�YUUUU�U�VeV�YeZ�eef��ef��j���ff��iZ��ff��ff��ff��UUUUUUUUeU�U�U�VUUUUUUUUUUUUUYUjfV��f���ff��ff��Uf��ff��ff��ff��UUUUUUUUUUUUUUY�UUUYUfUjUf������fi��ff��ff��ff���V�V�V�V�j����feUUUUUUUUUUUUUUUVUUeU�U�U�U�UiV�V�Z�Yff�if���ff��iV�Vf���ff��ff����e����������f�YUUUUUUUUUUUUUUUUQEUUEUUUUUUDDDUUEUUUUDDD@QUTUUUUUUDQEUUUUUUUU@QDDDDDDTADDDD       D A               �E�U��T�U�D���              QQDDDDD EADDDD�����j�Y�Z�Z�j�j�����ei�YeZ�V�V���h�������������Z�V��iYf��fj��fj�i�Z�ZfZ���V�V�Z�jjZ������U�UiU�D��D���U�U�U�U�U�U�UjU�UiU�U���Zj�ii�ZV���e���je����fZYY�V�V�������e���e���U�V�V�Y�i���je�YjZej�ii�����f���jj�j�Z�V�Z�j���j��j����jj��ij�j����������f���j������������������j�UUUUUUUUV�Z�V�Z��V�Vf�Z�Z�����j�i�ZUYUV�fef��eiVjV�UU�UUU��U���Y�����j�Zff�Zjf�j�Y�Vj�YeZ�YeV�VeV�Vf�i�fejUj�f�Ye���U���ef��if��UjeZej���Z�Z����jV�V�U�U�U�UfUjUjVjV���ij�����j�Z�V�V�VUYUVUYU�U����������e���e���j�UUV�fU��j��������Z�VjUYUZUVUjeV�U�U��feZ�Z�ZVUVUUUUUUUU�UeUY�Y�VZiV�V�V�V�VUeZ�Y�V�V�V�U�U�UUUU�UeU�U�U�U�U����V�UiUjUYUZUZUU������f���V�U�UVUZUeUfUY�Z�Z�YeU���eZ���f��e���Y�Y�V�Z�f�Z��Z�Y������U�U�UiU�U�UfU�U���e���e��j�iUj�������V�UiUZUUUU�Uj��U�Uf���f�j�j�ZUZUV�V�UVUjU�UVUYUVUYU�Ue�������j���f��f����i�����j�������i�����V�U���U�U�U�U���i�����������j�����f�����U�U�U�U�U�U�U�U�U�U�U�U�������V�U�U�������f�����Z��fV�UeU�V�UUUU�Z�U��V��iVZ�YfZjU�UZVYYf���e���                ��*�*��(�*�������*�*��(�*�����U�V�V�Y�Z�i������&��Xb�$�@@j�������
��(����f���fd
�b$������ff�&f�$F�ff�Yff�&f�$F�ff���U�VeV�Vi��Yf���f���f�i���������ff��ef��f���f���ff��f���Z�����j�ff��ff��fff��eiVff��ff��ff�Y���Yff��ff��ff��jf��f���f���f���f��� � � � � � � � �ff���f���f���f��ff��ff��ff��ff���f�Z�j�����������Z�j���j���j����ffY�ff���fi��Z��ff��ff��ff���e�����j�������fi����e���Y���j������ff�YffeYi��f����if��i���i�j���j���������������������f�����j�����ff��ef�Yf���j���ff��ff��ff��ff��f���j������jj�����������ij������ef�Ye��Yi��Ui���ff��ff��Zf�Yj���i�Z���j���������������������j��������������������Z�ieZ�iff�ii���UUUUUUUUUUUUUiV�U�V�Zei��ii��f��Z�V��f��ff��ff��UUUUUUUUUUUV�Z�YUUUU�U�VeV�YeZ�eef��ef��j���ff��iZ��ff��ff��ff��UUUUUUUUeU�U�U�VUUUUUUUUUUUUUYUjfV��f���ff��ff��Uf��ff��ff��ff��UUUUUUUUUUUUUUY�UUUYUfUjUf������fi��ff��ff��ff��UUYUiUj�����ff��UUUUUUUUUUUUUUUUf���ff��ff��ff���Z�Yff�if���ff��iV�Vf���ff��ff��jf��ff��ff��ff��UYUiV�Yif�Y��f��QEUUEUUUUUUDDDUUEUUUUDDD@QUTUUUUUUDQEUUUUUUUU@QDDDDDDTADDDD       D A               UUUUUUU�UeU�Vie�              QQDDDDD EADDDD � � � �D�Q�D��E��D��D��D���Q�U�U�U�U�U�U�U�U�U�U�U�U�U�U�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������0
�����6����7�ŀ�8�ƀ�9��:�@�;���1��2��3� �6�4 w��:�>�;�? ���6��7�:i�:��;�3���3�:iX�:��;�;�1�1��о�2�2��ж`�4JJJJe9�=�4)



e8�<��=`� �������<�>�>��?�����>i.�>��?����`ˀ�[�{�;�k� (  (((     ( )*((  (((  (  ( }+h[ZIH/ (  ( (   �|{fdYP?>. ((      (�zyb`ON=<-( ((  ( ( �wu_^ML;:, ((        sq]\KJ98  (  !01@AQRaQRar��� ( ("#23BCSTcSTct���( (($%45DEUVeUVev��� (  &'67FGWXgWXgx�� (  ( (QRa1@AijQR���� ( (( STc3BCklST����((((( UVe5DEmnU~����(   ((WXg7FGopW����� ( ( ((  (           (((( (((  (  (    (   ( ((( ((((( (( (((((	(((
(((((  ((  ((((  ( (((                                                                  	          
                                                                                                                                            5 9   >?G@MH #6784;<=####N####23  AB###O ####01  CD#SW  ###/.   EIT    *+,-   FJUV  ##(:     K#Y   #'    LRZ     #&     QX    !$%       P           )      																		
""""""""""""""""""

""""""""""""""""""

""""""""""""""""""

""""""""""""""""""
																		 @T�T�T�� �T��* ��0�����������������0�� �   � ���3�3�3�3�3���    ���������������  �<<<<<<�? < < <<<<�  �<<<<< ��� � < < �?  �?|�\_�p�p��W?|��_ p��W�W}|U��    �p5p5\\ \\\5\5\5\5\\�  �U�5�5�������U������   ��W��ppppppppp���W �  �����\�\��� � � ���\�\������  ?�5p5p5p5p5p�UU�5p5p5p5p5p?�  �W�����W�����W�  �?U5�?      �U�      �?U5�?  < � � \\\5\�\W\_\s\�\\\�  � ׀� � � � ׀� � � � � � � �   * � ?33� * ���k�[�[���� @T�W�[��+�kի������TP +�k�k�k�����UU  P�������UU�������k�+�k����[�[�j�����+�k�k�k�+�j��*                             P �                     = � ��9             ������� �   9 9 � � � �                 ��:Z�V�F���� �T�Tk�V��E�A�Q������� �nQnPnPnT[T�����������������������F�Z髺������[�k����                 ; : � � ����V�� �          ����� 8 � � � � � � �j � � ����PP�@[@[U�����Ð@�~��tG� 0����U�TTAU��Z �����嚥����+�k�n�n�l�l+�+�+���P�P�Q�Q�A�A�A�+�����Z�����A�A�A�F�F�K�K�F�Z鯾������+�jբ*B�A�A�A�E�V����+         �44�        9������[������VjU���� � �       � � �Q��k�V��Ao@n���������/��@�
  @}������Q�@��  @ �@}�      @���}������kU[  TT��?��U� P  U�V�k������������k�k�+�+lk[����������[@TV�[����������k������j��k�k�+�+�Z��* �         � �T� � P @    ���W� � �0                                  ��������30���   _ �             W � � � � ,,>, @_�����T�@� ��6 6 = = ��>��������A�@�P�        �+効���+�
�R��*�9�6���i� �  @T�T�T�� �T��*       � � � p  �T��Z�����/ �A������*���������J�������*���������J�������*������ZT����J����k�[�k����                �?��k������                ��������V:�6f��~� � [P[@l��V૕���e�[�~�������� � �T�T�T�� �T��*��iiY���iifje�ڦ��Yi�if��if��Vf�i�f��i��fi���Zf�fp����e�Yך��� ��=e楙�Y��e��[  VU[e�j�k � p p � � g g���o��k�k�k�kU���� @R�[�k�+�+�kի����Z�F������k�k�k�k�k�kծ������������jU   P���A�@�P����������*�����Z髺��
@Z�Z�Z�
�
�R��* @_�����T�@� �� �ԫ�VllPT�������A�@�P���[�kQ�E��Z�k���*�䊐���A.A� �T�T�T�� �T��*����Z�k����� �����ZU[ [U���� @T�V�V��
�Z��* � � � �        
@V�V�V���Z��* � p � � l � � �               �
@V�T�T�� �T��*E����@�U��+�
 ����jUU  UU����@[�n���钥���Q�����UU  UUUU������.U�@�U�U���������.���钥���Q��*��T�T�� �P��*E��Z�kQ�E��Z�k                UUUUUUUUUUUUUUUU                 � � � ��������� � � � �������������������������   ��������������  ? � ���?��                ����������������  ? � ���?��������� � � � �   � 0  � 0     0 �    0 �  ? � ���?������� � ����� � � � � � � � ����� � ������� �  ��������������������                ���� ? ������<?���������                 <    ������ ���?�?�����������   ����    D      D �0_��W�W=\� ? �\�WpUpU\U\U��  CUCUCUC�CY�� � �U�U�U�j�E�CYCYC	CUCUSU����E�E�@�U�U�U����� \W5W\W� ����������?�?������T� m mT~�������k����z]y��?�?�����������|UWUWU|UpUpU\U\U���������������UpU��<< 7� ��_����o����������   7=��UUUUUUU�0W�WUUUUUUUUUUUUUUUUUWU\U_UUUUUU5U�50<           � _UUU�U�U W \ �      UUUUUUWU\U\U\UpU           ��upU�U?W \ W�U�7W�U�] s �    �\�WUWU|U�U|UWU\UpU\U\UWUWUWU|��� 3   � p p p p �    UUUUUUUUUUUUWU|U�� �            UU]UWU\UWU\U_UpUpU�W \ \ \ p p p �                              UUUUUUUUUUUUUUUUUUWU\�\��5                   � � � 5  5 5 5 � � � 5 5 5 5 5  �  5 � 5 � �                 U�UUUU��3�s5]�_U�U�_U�W�  0  U� ��3_ \ �� p               3 � � � 0     UUUUUUUUU�U5U7�U5U�UUUUUUUUUUUU0��3<50  UUUUUUUUUUU�U5U5U?� �UU�0����0 ��WUUUUUUUUU�    ? � 5 �U�UuU]U�UUUUUUUUUUUU3 ��U�U}UUUUUUUUWU5U�UUUUUUUUUU            � |� �    �       �s��U5�?     3��UU�W �    WUUUUUUUUUuU�W \       � \�W\U\U     � s�]uUUUUU  ��U�U]UUUUUU W�UpUpUpU�U W �UUUUUUUUUUUUWU\U 0   � � � �    \UWUUUUUUUUUWU|U�U�U W W \ p p � �         � p �    ? ��U_UUUUUU      0�5W�U�U3UUUUUW��0 5 5 � � W�W]WUUUUUUUWU_U\U\U\UpUpU�U�W \ \ \ \ p p �  ? � UU�UuUUUUU�U5UUUU5U5U�UUU� UU� ppp�         WUWUWU\�\�\�\5\UUUUUUUUUUUUUUUUUUUUUUUUU�U=UU�5                 <3��UUUUUUU  0 � UUU5UU5U�U�U�5�5�                U5U5U5U�U�U5U5U5UUUU� 5   ������'���3���?�ŤK�ѧW�ݪc��o���   #                 #      #   #                                                                        #	     #	#     	#      	                                                                                            !"!"            #    !"#     "!                                              
	         	
          !"     #     $  $  
  #  
  "      !              	      $
  #                                
   #  $!	  ""!                                                                      "    "                                                 $  ##  	  	  $    ##                                                              "        !  #"  "# !         #      #          "                                         #!!#              	       !      !       	    
               
   	           $                 
$            "        
"       	            !   	    #      	     	!                           	#                                                   !             "   ! 
 " 
    
      "   ! 
    !             "              !               ! !        !       #               #        #           #  
     " 
 "     	        "    ! $ $    $"! $     	                       !      
                         
                     !                        #$
      !      !      #   !
#  !    #$   
            $      
$        
            $                    "   "   	     $ #         #       	   
              !	    $$   !      	           $    $     ! !    	            	     !      
!  
        "  	##  $  	  $		  "      	     #  	   	          #           $               	 "            #"    $  #    
  	  !     ! #  	             ""                  #       
   !!  
                         	    $     	         $       
  !!   
	
	 		
 
               !  	                                              $	  $!                                                                         !            !      " 	

! "

 	            !                              "         "                      " "	                         	  	  	     $    $     "                                 "   
		$		 
$ "
#"##            	        	    
    $        $            #		$$	   
"  !	  
  !                            #   "  #  #	#    	
$##
$"$""#

"#$   !! !!!
 
  
 
	!			!#"!#!""!	"	 $  	

	 $
$
$##      #  "          
  	  
   	        "   #    
                     
     !       
       "              $$       $        $!   "
                                                
  
   
 
                                                                                	"    	"    
      "" 
                                                       
       #                !   #$#  !  $#
                        

"!"  !#	
! 	" 
"$	!	$###                                		  $  	$	        ""                                     
	  "#	  #"$  #$
  #  !!  		""                          $    $"  "
"  "!  
  !    

               
#    
$! $	 	  
$"""$"!
#       !      
                         
                     !                                     !"                 "     $   !       $    "     "           !$ 	"$ # #	 !	"	 
 
##  

$$	!
!
$           $   	  $""  $#  	"#  	"           
      
# !"	!#"	"# !		"!  #  

                  "  	!  ""  "	  	  
!    $  	$  
$$           !
 $ 
$
 !		
! "!"#$	"$"	#"		"!$! $"
"
 #$!
	# $	 #!#
           
!    
$    !#  !         !   #$             

$!  !  "
                 #                 # "     $  

#  #	
	!$!$          !   !      $ #$		#  �����                                                                                     )3== [       9
 *4>HR\fpz  �w1	!+5?IS]gq{���v0",6@JT^hr|��eu/#-7AKU_i }���t'$.8BLV`j ~���s&   CMWak           DNXbl           ;EOYcm         (2<FPZ          ���o%           ���n            Gy�             Qx            d              :                                                                                                                                  huvLY"#   @MN[ ijw Z\$%34ABOP]^kl!.gq&'5 CDQR_  n/0m`()7 EFSTabop1:86*+9 GHUVcd r >2,-;<IJWXefst?K            
	                                                                                                                                                                                                JI     /=>KLY <MT '"#0 ?@@@[ NO;:$%34ABBB]^PZ98`\.7b!a2_X,+
1WV*)	56CDQREFSGHU&&&&&&&&&&&&&&&&&(((((((((((((((((dddddddddddddddddeddddddddddddddddedddddddddde V   dddddd        ddddd 7FG       ddd 89HIW      
ddd	 :;JKX       #,-  <=LMY     $%./ `>?NOZ_!""""&'01"a@APQ[^()23bBCRS\*+45cDETU]                                                                                                                       "               #-7          )$.8B D   I?4!9CM:ZVQH>3 
&0N/]YULG=,	'1;EO%\XTKA6+(2<FP[WSJ@5*GGGGde^YGG_`jGGGGHGGGGGgZ[UVabGGGGGHGGGGGGG]WXcGGGGGGHGGGGGGGGGGGGGGGGGHGGGGGGGGGGGGGGGGGHGGGGGGGGGGGGGGGGGHGGGGGGGGGGGGGGGGGHGGGGGGGGGGGGGGGGGH"&*+GGGGGGGGGGGGGH#',-2GGGGGGGGGG@AD#(./4589IJMNQR<=BE#)0167:;##OP#T>?CFhhnmnmopLop	S$ik	%Kl\3
               ! "  #$12    %)*+,0      &'(    -./   @34KLW B56MNYZ D78OP[EF9:QR]^GH;<ST_`IJ=>UVa?AAAAAAAAAAAAAAAAAXCCCCCCCCCCCCCCCCC!   
	
	
	
	                                                                                                               
	                                                    "#  VWZ[^_9 !$%?@XY\]`01*)'&25AB4444444444+(36  CF444444/.-,87    D444444=<;:     GE444444     IH4444444    KJ44444444     ML444444444    PON4444444444UTSRQ44444444444444444444444444444                                                                               	
                          CD FCD FCDIJQRghszABGHABGHABKLSTijt{=>?@=>?@=>OMa_klu|<<<<<<<<<<<NU`mnv}'(+,/03478'PVbopw~)*-.125)9:)*Wcqrx))))))))))))Xd��y�))))))))))))Ye6;�f"#^]\[Z !$% !&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ 
��)@�� � ������ � t�`�Z�K��[�_��\�����[�s��� n� C� C��[�\��` 
%*5AFLSZ`fiou�
	
	                      ��)�7��)���H���Z��� ���H���Z������ �l��� ������`CIILPKLRJJHIFHJKMS�u����[Io>`��<��<    �Y��,���Z  ��Y��,���Z  �`���& ��0  ����� ��Z���V��  � t��� ���� ��B�ɍ& `�B��]� � c� 5� �� �© �B`�� �t�v�r�r��
8��r�tL��`� �����r������`� ��������`�v�vɥ�*�v� 	��q� 	�q��w� �� ���p`�৐��v�vɦ�֩�G ��`��� �� � �ʥ��/ T˥��( �̥��!������x�  ͥ��榥���� ©�p`���� ©�p`�w�wৰ�v� 	� 	���p`� �p`�]�����p� #�`�� ]�`��� ��`�^ �ѥ^���G�G�'Å�*Å�@�����-�0�� n��������� ��������C`nkn 	�� ��m0C�)?�=�l�9��l�m�I0 � �`� �G ��`� ��nȩ��n�ni0�n��o�	���`���; Lå��x�)��r� ������� ������� 	�\���P���Q�Q� �� 
�� t�`��A��ɴ��)��4� �� ���`��� 	�� �� 
��%�j ���`汦�ഐݩ� ��`������ 	�� �� 
�� 	�j ���`汦�ഐܩ ����� 7�`� �A��@�P�
�@i�@����Q�
�Ai
�A��� ��`�S�W�P�R}�ąV��W�Q�V}�ąV��W�W}�ąW� �b�b��ąc��ıV�d 2��b�b��� �� �` 	
 $6Zl~����� 2D              " �Q)


��P)�� ��e� �����e������`� � ��������� ����`�dJJJJeU�Y�d)



eT�X��Y� �c��f�X� ���f�������`�a�P�P��� �P�Q`�B� Lĥa�� t� hũ �B`�a8���� 
�� � 	���j �� hũ �B`�j
����ཎ�� �������� �`�D�\ƍ& �
��oƅ�nƅ���g���S�W� �R�V� ��V C��V�V��W����������D�8ƅ$�& �Jƹ ��T���U�$		�$�& `������������������  

������������������ �h����P��� ����X���LӼ�T��ش�քש �P�Q�a�B�� 	�ഐ��
��E��y�ƅ��y�ƅ���� �k��g�
�f��� 	��k���f�����g��`   ���������� �� 
��)�@��� � ��DǑ������ �����B��� � ��=bǑ������ ����Ɖ�` ��? � � � � � � � ���? ���?��?��?��?��?��?��?��? ������ �� 
�� 	�	�P �� t�`�j ��`����ǹ� ����}�Ǚ� ���������� �ǥ��� ;˩ ��`    �������� 	�2戥�����������`��	��ť�ƈ`����� 	�� 	�� ��膦` &�`�_�B�p��<�v� 	�)��w� 	� ����_ �� �ǥ��ƈ �� © ������ �p��v��w`��� �ƥ) � ��`�)� �`����������� �����=��� ��搥���쥄���`� �����=��� ��搥����`�������� �� 
�⥞����i&�j ��Ɵ��`���P���Q�Q� � 	 t�Ɵť���Ɓ�`���<��)�6����� ����� �恥�ŀ��`�� ��`����� ��Ɓ v�`�p�� �vŤ�ť�
�wŤ�ť���v��w� �p` Oɥ������������ ����������k�k�k� ��`�_i�_�
��	�_ ���D�D��� �D��)��^�^�
��	�^���� ���]��`��� �P� �� 
�� �� t�`��Q�P��
8��P�QL��`��� � 
�� ��@�4ʠ �:ʙ������ �` <Zx�       TU ��@��@��@��@�U@�@�      U �_ �����U�@�@�@�@�@�U@��@��@�� �� TU      @�@�U�������_ U       @�@�@�@�@�@�@�@�@�@�      UUU������������UUU      � ����8塅���8壅������������`���
��������� � 	� �ഐ������ ����� `�𵠅��
��i������`� ������������˅���˹� ����˅�ō�'����}�˅��� �(��� 抩����}�˅�Ŏ��拥�����������`���륊)�������`����    ����������8��˅�� ��˝@�䀐�`����� ����8��˅�� ��˝@�䒐�`� ����)�
接�) �接�)�
接�) �掦����@��� �` ��)���
���D̅� �˦�� �� ̥�)e���Œ���)�JJJJ)������ �˩ ���������������������� 	�j� �� 
�� �����`� ����������� �|��˅���˹� ����˅�ō�+����}�˅��� �,��� 抦��|�����}�˅�Ŏ��拥�����������`ɀ����`����� �������e�����ͅ���ͅ���ͅ��������͹� ��� ��������e����� ���-敦���}�ͅ�ŝ�ᦦ��ͅ���ͅ�� ��Ƙ�攦��xЖ`ɀ�ߩ��`��������  ���������� �˦���� ������ ̥�e���Œ���JJJJ)������ �˥���������I������ �急�����)�e���������JJJJ)�� �� ��`� ���������`���d�� �ʥ�����!� �� ��`�`�� T˥������ �� ��` &�`�� �̥������� H�`��妦�x��  ͥ��н����΅� ��` ��i0�����`��



���� ��Α������ ������`  �??????????�  �������  �????��< �?  �????�????�  �?????????�? ?  �?? � ?????�  �??? �????�  �? ? ?����  �????�????�  �????�? ???���H



����h��� ��ϑ������ ������`� ��Б������ ������`  �<<<�?<<  �<<�<<�  �<   <�  �<<<�  �?  �  �?  �?  �     �< �?<<�?  <<<�?<<<  �������  �?   �  <��?<0        �?  <??�<�<�<�<<  <<?<�<?<0  �<<<<<�  �<<<�    �<<�<?<�3  �<<<�?<  �< � <<�  �?������  <<<<<<�  <<<<<<�  <�<�<�<�<�<<  <<��<<0  <<<����  �? < �� < �?                      �?�?         � ��?��   Rҩ����v�������� �C�p������`�V�ᩩ��^�� ��`�#)���хE`      ���B��  ��)��� �B�� �ѩ ���D� �& ���^�_`�[����_�� ��`�D�ᩩ��I�� ��`�<�m��l�F��o���⩹�n��� ��ȑ� ޢ<� ���ȩϑ� ������ ��ȑ�`��I � ҩ�����҅⹕҅㾒Ҡ ��ґ������ �������� �� ��` 8pASX������\]u5\s�5��?7\�5�� 7�� 7��?7�  7�  7\�5\��5\W�5������\UU5\_}5���5���7���7���7ܢ�5\�z5\�^5\�W5\�U5\UU5������\UU5\�5\��5\_�5\_�5\_�5\_�5\��5\��5\_�5\_�5\UU5���������`                                                   %&             ?A  '(     367 ;=@BCEF )*+ 154T89<!\]DHGJKL,-.RSUV:YZ[^_I!!!MN/0!!!WX!!!!#!!!!!OPQ!!!!!!!!!!!!!!!!!!!!!
	`b""""""""""""a2"$                  CCCCCCCCCCCCCCCCCSCCCCCCCCCC78CCCCCSCCCCCCCCGH9:UVCCCSCCCCCCCCIJ;<WXCCCSCCCCCCCCKL=>YZCCCSCCCCCCCCMN?@[CCCSCCCCCCCCOPABCCCSCCCCCCCCQCCC3DCCCSCCCCCC$*-CCCCCCCCSCCCC%+.CCCCCFRCC&,/CCCC	0E 'CC5
14(62) !"""""""""""""""""#                                                                                                                       CD FCD FCD FCD FCIABGHABGHABGHABGHAJ=>?@=>?@=>?@=>?@=K77777777777777777L'(+,/03477'7	6<E)*-.1259:*8;"#
!$% !&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&                                                                                     )4>              5=@AHK        bfg*+67BCNOZ[opu !,-89DEPQ\]qr"#./:;FGRS^_st($%01<  ITU`    &'23   JVW             LMXY     nmjk  cda 	       lhie   
 	           	
           
                                                                                                $%6            &'89           ():;           *+<= mnuv}~PQ,->?  opwx�RS./@AHLklqryz�7TU01BCIMst{VW !23DEJN\^
	XY"#45FGKOZ[_`             ]ab            cd           ef           gh           ij                                                              "#*+23:;BCJKRS$%,-45<=DELMTU&'./67>?FGNOVW !()0189@AHIPQXYZ[Z[Z[Z[Z[Z[Z[Z[Zl\]\]\]\]\]\]\]\]\m^_^_^_^_^_^_^_^_^n`a`a`a`a`a`a`a`a`obcbcbcbcbcbcbcbcbpdededededededededqfgfgfgfgfgfgfgfgfrhihihihihihihihihsjkjkjkjkjkjkjkjkjtvwvwvwvwvwvwvwvwvuuuuuuu
	                                                                                               }~�              �e            ���2|�{       
 AP\]&Iyzyz	uvw3@w'45BCOwf()67DEQR[w'*+89FGSTQ^ghw,-:;HJUV_`ijox"#./<=KLWXabklqr$% !01>?MNYZcdmnst����������������������������������������������������������������������������������������������� ��@��/� ��� ����`��� ������ ��� �� �䨑��������` �ݥ@JJe����`�AH)���݅�hJJJJ)����yޅ�` 0`��� P���@p��@@@@@@AAAAABBBBB 	��i0����`�I�  ��  �`���& ����������  � � � � �* �	�
� ���[�� ������& ����� �� Hߥ��������i<���`���`���>�]�:��8� 5�i0��i ������������i0���i �������  �ߥ�a�.�]�*�D 5����ȑ���� ��i0��i ������ ��_��a�Ș p��a����`�`���`��K�]�G��8� 5�i��i ��i0��i ������������i0���i ������� �ߥ�a�0�]�,�D 5��ȱ����'��� ��i0��i ���ߩ���a����`�`



}������i ��J��� 5๑�e��i ������`� � ��@����������`H)��P��hJJJJ�
ei@}`��` 0`��� P���@p��      

�� ���� � �����`� �/ ����� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                  �����ȱ�� � ����0��� �J���� � ��� �* ���`����Q� �  �ܥ
�������`� � � �� � �����
����`
��������
���ȱ���� ��	�� ��L�� H�L�� *�0Y���JJJ����	�Bȱ�4�

��4� �)�7� �� �"JJJJ�%�)pJJJJ	�1 �� � ��`� �.�>�����k�L\��+��%8�(�%���)�+ �� h�`� �.�% �� h�`�+���(}%�%����)�+ �� h�`�.�� �� �� h�`�+�Ž%8�(�%��")�%L�")�%���ǽ)�+ �� h�`�+� �� h�`� ���)����1��)pJJJJ	�1�

��)�%�48��4��7� �4�7�4� �7� `�4e�4���7�7��ީ�7���4�ҭ �

��)�JJ%	J� `���� �.`
em ������ )�+�JJJJ�(��.`�����e`���ȱ������.�@���*����Q� �  `��ý
��
��L*���ȱ��
�L*���ȱ�L*�
qm �����ȱ�� �L*�05

������� � ����)� � ���� � ��� � �	�	�c��S)x�OJJ�����C��?�0&�8���
�� ���� � �� � LN�e�������ܩ ��	�� � � �0

�������( ���) �
���* �
�	�
�� �* `� o�_Cb4 � ����%�u�}���I���K����+�S����c��y�c�o�%��������@!T! <a@!T"<!TA}  !@ � <a!@"<!@AT  !T! <a@!T!�!TA}   �0�@� �!!@!}A�   +�+��.. �.}.� � �ThT.T��A}@  i�i���!@!}!�R  ���.	@h	.@	h�	�A�   ����	@	@h	@ !@1��!}!��<!�A�!�1h}!�!@!}� } !�  Ha� Q� 	@	@h	@ !@1h!}!�!}!h@h!@ �1h!}!�!}!h1@�  � � �0��!@ � } 0��	@ !@!�!}0� � � � �0��!A@    i�i��@1. �!!.!T} !}!.A�  1. �!!.!T} !}!.A}    �����1}T!}a�1}T!}a�8�  �a.9 !a}9T !T1.!T1}T!}a�9T !T1.!T1}T!}a�8�  �0��!.a`�!!}!�1}�!��<    ����� �  "� � "  @ @ h h A�@ � �  "� � "  @ @ h h A�0 � � 1�� � !�  � 	� 	� !�!�a�    ����@"<� � ���}T T ThT@  .�A  !T@ @T!}!@T T}!�!T!}!�!�!�A}  "<� � ���}T T ThT@  .�A  !� �!!@!T!}!�!�!�!}T@T } A�    u�u���T}� � !���< < "<�}T T T}�}!T} !}T}� � !���< < "<�}!T T�}  z!T!}!� !T!}A�T!T !T!T!  @ �@�  �@ �@� ���  � !T !T!}�}!T T�}!T!}!�  Y�Y���!�} 1}�!}. !.!T� � 0�!.!T!.  !�} 1}�!}. !.!T �T 1T}!�!�!�  � �  �!}!. !.!T� �  �!}!. !.!T� �  � �!!.!  !T.0�	} !}!T!.   � �  � �!!.!  !T.0�	} !}!T!}    1�1���A�!T 	T ATA.! 	 1 1 !.!@�AhA.1T A�!T 	T ATA.! 	 1 1 !.!@�AhA.1T    � �!`� � �� @�  �  �!.`��  � 1 A�!T 	T ATA.! 	 1 1 !.!@�AhA.1T   �����@1@!T!}!�!}!T!�}T@}1T}!�!�1� 1@!T!}!�!}!T!�}T@}1T}!�!�1� 1}T!@!}1T@!!}T.!�� � � �1 1@!T!}!�!}!T!�� � � �1@!T!}!�    �������<��@aT�<�<�Ta}<���<������  PT}�}T}a@ T	} }�}Ta}@ @ !@aT  !A@  @ @ !@AT!}a�} } !}AT  T T !Ta�} } !}A�!�R�   Q�Q���!@	@} } }	�}	h!}  !h�	@!}  !�<	�"�  q�@h}�}h!}  !�} !}�	T�� .�}!h }�!@   ��h} � ��<���}h  �����@�}h@!@!h!}A�}h@!@h@h}�}Ah�}h@!@! �!@@!�}h!@!}!�    O�O�����}T.T�T. .	A.T.T� �		.	T	}T T	.1T T.T� �		.	T}�}T}�� ��}.T}�}� �
\1�   ������!@T	}1��!�"<"� �!} }!T TA@0 	@ @T}	� �	��	@ @T}	� �	�	� 	� 	� 	� 	� 	�	�!� 	�	�
< 
< 
< 
<	�!� 	�
<�!@}�	���� < "�    ������� �}T T}� !�! 	T T T}!�}T� � !�  @ @ !@ ��@!T!	@ @ 	@ !@ ��T! 	T T T}!�}T� !�! 	T T T}!�}T� � !�  T T� �T}�}T!@}�  �!�"<!�"<���}AT �!� �!!�A�@   {�{���� � ��}	@ A@Ah} } }���b<  < < <��	� A�2� � "�<����}@ !@@h	} A}B<h !h}�}@��� � ��<�@ !@Ah� � �h}�a�    +�+��!h!@h� �h��2 @�h!@!�ah  @�@1h @�@1h !h!@h� �h��2  �1� @@ �!@ah   �1� @@ �!@1h@��h@ah    ������h 1h !�!h1@ 1� !!@!!A@ h 1h !}!�!}!h!@!1} 1�	� A�@ 0� !!1 1 !@!!h!@1}�� h !h!}!h!@1h �  !!@!!1 @ !!!!@!h1} !h!1 1@	h Ah    ���	�T T	}	�	}	T	@		T		T�	�	� } }	T	}	�	�	�
<
�
<	�	}	�	}	� � !�	}	�	�	�}T@� } }	T	}	�	}	TQ� 	} 	}	T1@}	T 	T	@1T  �	@ 	@	0����T� |	. 	.	0�.���.@	T 1T	@	T	}	T	@		@	(�		@	T	} )}	T	}	�	}	TA�    �����9�W�u����������)�G�e������������7�U�s���������	�'�E�c������������5�S�q��� ����������?�� ��������?���+�+ �+ ���������������?��?���������+ ��
������������?��? �?����������?� ������?��?������+�+�+������������?��? �������?����?� ������?��?���+ �+��+���
�+����������?��? ����3��3���� ������?��? �3����3����3� ������?��?������+ ����+ ������������?��?0�<��������<�������?��? �<�?�<�<�<� ������?��?��������������������������?��? �?����?����?� ������?��?������+��+��+(������������?��?���+*����������+*���������?��?��������������������?��?���������+ ���������������?��? �?����<����� ������?��?������+
�������+ ���������?��? ������<�<�<� ������?��?���+ ��
������������������?��? ���0���� � ������?��?��� ���+ ��"� ���������?��? � � ���� � � ������?��? �?����<����?� ������?��?������+
����+
������������?��? �?����?����?� ������?��?������+����+������������?��?����*����������+����������?��? �������� ������?��?���������+ ���������������?��? �?��<��<����<� ������?��?������+��+��+ ������������?��? �?��������?� ������?��?������+�� ��
������������?��� � � � � � � � ���������� � � ����WU�WU�������������������WU�WU�������������������WU�WU������ꫪꫪ��������������� � � �* �	�
`��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xة �& ��  5� O��F�
�� �� �� �� �� �� �� yťa���� y� 7� ���]��C�L�� ��Fп�� ���^�L���� �� ���H� �B�B����)?��H�H���)����_��_`�� �� ���H� �B�B����)?��H�H���)���`�D�B�� ��`	
�������
��O��ׅ� ��`8�
��O��؅� �ΩO��օ��� ��`���& ��0  � T�� ���H�]�� ��ɍ& � �B�B����)?��H�H���)�����&  ��`�)��)��������F�����V�� n�`����)���+��b�-��c�V����b�/��� n��b�����c��`��  ���&  �ݩ�������� � ��� � �F�B�0  �� �� ���ɍ& �B�� ���)���)@�� � ���FI�F� �B�ک ��F�
���� �& `��� ��� ��D�E�B ��B���)��إ)@� ��� �B��`�E�E��� �E����� ���D��^�_�V�᩟��E���� �ΩV�ᩝ���� nϥ�b�b�b�
�8�
�b�V�ᩙ���� �ΩV�ᩛ��b�� ��`H�H�H� � ��  �� ��B�	 &�惩�B��#e�#h�h�h(@������������������������������������������������������������������������������������������������������b�����