L�L��1��� ���������2��3`�1
��4��-�5��.l- H�d���������WWXXDF�Ʃ �<������/ ނ � +� E��1`慥<
��w��-�x��.l- �����QJ[JQ�����XUJJI������)�6��)��)���)����
΅ E�� �`������ E�� �`�<��� �/�L�$ 怩�/�R�$��#��(�/�#��$��}��+ 2��/�#�#�(��`��)�
�� +�L ��+ /��)�+)�3��/)� �<��/�L�$ 怩
�/�R�$ � +���`� �/ ނ�<��)�����)�����ߩ �+ /�� +�� �`���ȩ �+ /�Ά +�� �`��)�
�� �L���+ ��)�(��$)�3��� ��<��/ ނ��/�R�$ 怩�`� �+ �· ���`����� �+ �� ���`VXY�8����+ �����
����� 2�`��̩��+ ���S����(�� 2�`��� ��� �!�/��������"�
��
�"�!���N��/�
iH��!i<�+ 2��/�/��� �/�*�(��J�'�(i �(�
8�'�(�)�*�'��*���'�B��+�M��/
i�� 2��+�O��/
i� 2��/�/�
��` ��� �(�/�8��+�@���D�� 2��/�(�(���`UZXM XYFWY          � 0�� ���� ��`��2�3`慥�)������/�
�(��# ���/���+�R��#� 2��/�#�#�(��`������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������1��&�
�"� i��9�� ���i� ��`�9�� ��1
��=��-�>��.l- ���� �Q�����/���⌃�7�#�YTUXHTWJXYFLJXUJJIGFQQAAAEEEEEJJJJJNNNNNSSSSlnp�����lnprt�����lnprQT\RJI MN�1 ��� ���'�B�U��+�k������ 2��'�'��� �� А��'��#� �"���!�
��
�!�"���'� i<�+�K��#� 2��#�#�'�䭆
m��'��(�p�#�'����+�P��#� 2��'�#�#�(�� ��� �� e���)


�>�����T�

i�=��=� �� 
��h��=��� ������?�8�?�@ c���
�A`888888000000000((  慥�)�`��%@�'m�ee5���'� 
��?�>���+i� � �)���JJJ���'�@� 
�(� 
� 
�(� 
�@�?�>�(� � 2��� �����=��1��i� ��`� �� %��1`�����������:��� �:�;`BBAA@@??d_ZUPKFF慦A���<�#�A���I��9�1��� �:�;���� e�������� e�� �!�" ����i�����!���" ��`����=����N� �!�" �����d���H��H %���������h��h���d8���������б����� �!�" �������К����� �!�" ���Ї����������������������� �����������
�1� ������������ ��`�1` (#	 
#� �/�,�)0�p����


e������������T����	�����E���@���, <��/��/� �+�" ߏ��I����)���� ����� ��L���e,���)��慤A�����[��� ���(��)�	�)�L����W���L�����)�k���g�������'���(�( y�� �L����


e��� ����1��� ���!��������������� ������ ����
� �x�����/����+���" ߏ`�)���)����ޥ��'���(� ���)��)�5��iŃ����' y�� �� <��/��/� �+�" ߏ�'���(��L�������'L닥����'���(�(L닩 �/���-���.���# ����-���.���#����-�!�.�-�4��+ ���8逅�� 2�Lz� ��/�
�1�1�1 *�`�1 ��� ��`慥���	�#��2�`�2�+ ��`�3�+ ����`� �+���� �� �� +�����1���� ����1�� ��`慥�)����� ����


e��� �2��.��)���)��	������	���憩 �+ � 2�惥����Ƅ�����1`� ��/)��� ��� �+�� � �H)���JJJ��� � 2�Ɔh���x�ǩ��`� �/��������� ����#���-���. ��惥�)����愥���ԥ/��18��1 *�`� �� ���1�1`LFRJT[JWXYFWY �������������������IIIILLLLXXXXXOOOOOPPPPPRRRRRSSSSS

�����	�����	��������2�&�' k� ��� �/�ԍ�+������� 2��/�/�!���` ���5)�
��� �+��҅+�O��� �� 2����2�3`XYFLJHQJFWYW^SJ]YXYFWY����̺���ͼ���ξ���������GGGGGIIIIISSSUUUUXXXXXKKKKKLLLLLNNNNNOOOOOQQQQQ�����
��������IKMOQ�����IKMOQ�����IKMOQ���2�&�' k� ��� �/����+�Ŏ��� 2��/�/�/���` ��� m�i� �� ����� k�� �������	��3��2`���̏�H��3��2`� �H���"����H� ���ȏ�����eH�H����� �1`
	DFGIJLMOPRSUVXY[ � 2��"�+����#�#L��$�#8逅#��$�#��$� 2�` ����
i�#���)��#i��#�Ϗ�$��#�`�%��&��+)



e��i ��+JJJJe���-��.  �`� ������ ��� �����`� � �(


e'�� �������� `���� `��%���&` ����'��#�'�i<�+�B��#� 2��#�#�'��` ����'�l�#�'��i<�+�G��#� 2��#�#�'��` ����'��#� �"���!�
��
�!�"���'� i<�+�T��#� 2��#�#�'��`

4  5

�������/��/� �+���4��" ߏ`688  67   6  ���Y�$���#��

�'��(�'�Y��+�$��#� 2��$��#i� 2��(��'�#i��#�$i�$��` 0`��� P ���@�$���#��JJJ�e$�$�Je$�$�)���e#�#��)����$���e#�#�$i �$� �'�'�!�+�$��#� 2��#e��#�$i �$�'�'���`��)������!�����"�������������� ���B�B��� �B�A�A����A`UFZXJ�9I�9� �'�(�/ ����#�(�)��#i��#�Ϗ�$�/� �+�9��+�� �+�#��$� 2��/�'�#�#�')�'���(�(����1��B�9�2� �+�" ߏ� �'�ǅ#�'�d��+�O��#� 2��#�#�#�'�'���`���+���" ߏ`�9��`�.


e-�!��$�-�%��!���������#�	�%�$����-��!���������#��$����$���/�!8�-e%���	�����$���$�.�%��!���������#��%�$�8�����.��!���������#��$�i����$���/�%


e-���	����i��$��`� �����H���+�  � 2�h�����惥����愩 ����`� ��)�)�� ���� �� �������`  (08@HPPPP  @P`p������ 0`x��������:�;��`�;��



e;��Q��'� ��!�����'�
��
�'�#��"� �!u���
��
�������� А���������� ������ ���� ��L��� ��� ��� � �:�����` 戥���I���E�/ ����H��H� ��� ����+� �)���JJJ�� � 2��/�扦����֩ ����h��h��` ��� �/�����+� � � 2��/� � �/�/���惥�)�������`�5)�)��/��I����/��0� �+������� 2��/�/���`�ԍ�+��@�:� � � J�-�@-��� � 
������ ��)�� ��-��I�L핹���	���`��� }T	}!!T!}!T} 	}T �	��  �!T T	}T} }T	}!!T!}!T} 	}T� �� � �!!T  x}	��< }	��<0 <�
<� � �
<�2�   �	� � �	  �} �}1    ����..Th���!h!�AT �@� � \ � � \ B )����!T!�!}!��
<�
<!}  !@!}!T!}�
<�
<!�  !T!�!}!T@	�@	�� 	�}	@	hT	hT}1�  f��2�� a�  �@  	@T	@! �!!@T	�T	�!}  !@!!@!T}	�}	�� 	��	�!}!�!}!T@	�@	�� 	�}	T!.! �!.�	@T	@T	}  �@X � < � < < �0 � � < � < < �0 X � � < � � � � < < < � � X �  � "�  � "�!�!�!�"�"�"�"�#X#X"<#�"�"�"�#X"<"<"�"�"�"�"�"<� � � � "�  "�  #�"�"<"�  ���@@}�} � @@}�} � @@} @@} ����  P\ �  \ � ����!�  ����!�  ��� ��� ����  �A} X!}!@@}�!}!�@@}�!}!�@@}�@@}�!�!�\�  ���"�  ���"�  ��"�� "!�<�    �E��` ����������������������	  @	 	2��!� �!�!}T	h}��� ���  @  [�ћ�T T}T@!@ @T}T!�} }�}T!@T T}�}T T T}T@!@ @T@�	�	}T T�@T}�A�@   ��CX  X�B<  �<B�  ��CX  X�CX  X�C�  ��B<"<"�B�#X  X < X � � � � � < � < � X < � < X < X � � X � � < < < � �  � < #X   ����2��	} !}�!}!�A�@ 	} !}�!}!�A�@ 	T !Th!T!�!}  !�  P  !� �!�!ā�   !� �!.!Ta}  1}T1}T1.T1}�!� �1��a�  1}T1}T1.T1}�!� �1��aT  1T.1T.1.1T1.1.Ta}  !� �1��1�}!.  1T.1`�    < � < � X < � < X < X � � X � � < < < � �  � < #X   ۝y��@T.T}�}T ��}��}T T.T}�}T 	T  L}��T�  � }��T!�  ..T}T. 	.T.T}�}T ..T}T. 	.	�	�	h	T.T0   �@� ( � ( �  �  � ( � ( �  (  J "�  � � � \ � � ( � ( � � \ � � �  �   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������1
����-���.l- ,�{���C�ġYMNS HMJS HTRUFS^� �/�c�# ���[��#��/����+ 2��/�#�#�/����1� �/ N�� �����E���C��D� �G` 8p8��6慥�)�.���/ ����JJJJ)��w��/ ���C�C)��D
�1� �D���C` t�慥�)���Cɏ�
���/ ��Lؠ�i�/ ���C�C�~��C)��E�E��� �/ %�� ���1`Ɏ��!�I�G��F� �/ %���JJJJ)��5��/ ��`��JJJJ)��w��/ ��` #F# 0H`x���إ5)�b慥���[�H�9��/���%��&� �(�*�S�$���#�/�ȥ�+�*
e#��$i � 2��/�(�*�(���*��֩ �*�#i��#�$i�$��`����1�H�	��P��(�/ N�`��H���	���2�3`��3��2� �J`��� !"#$%&'()*+,-./ 123  6789:;<=> @ABC 123  67DE:;JFG @KHI 123  6789:;<�� @A�� 123  67DE:;J�� @K�ߩ �(�* ���S�$���#�/�ꡅ+�*
e#��$i � 2��/�(�*�(���*��֩ �*�#i��#�$i�$��`���%�ۅ&`     	
        !     "    #         ()./4$%*+015&',-236   :987   ;  @   <  A   =>?B  JKTU CDLMVW^EFNOXY_GHPQZ[` IRS\]a   b  f   cdeg                                                               � �(�*�C�#�A�$���%���&�/����+�*
e#��$i � 2��*�/�(�*eD���(�8�'�ѥ(eD�8��(� �*�/eD�/�#i��#�$i�$Ь`   OPQR  UVWXYZ[\]^_`abcdefg    lm          xyz{|}~����������          ���� ������������� ������  ����                                     ��ŷ�  ��  ����ô��������  ����ô�ȷ��ɻ��������                �E�(�*e/�/�C�#�A�$ ���/��+�*
e#��$i � 2��*�/�(�*���(�#�'�ԥ(eE�#��(�E�*�/eE�/�#i��#�$i�$Я`� �(�* ���G�$�F�#�/�}��+�*
e#��$i � 2��/�(�*�(���*��֩ �*�#i��#�$i�$��`�G���S��Fɀ�`��)��0�/ %��Fi0�F�Gi �G�S��Fɀ���/ %��H�	��<���/ N�`� �/ %�`    	
'!%("&# $)*/078+,129:-34;<.56$ =@AH  >BCI ?DEJKFGL MQRYZ NST[\OUV]PWX^ _cdk  `efl aghmbij^ nrsz{ otu|}pvw~qxyL        ��   ������ ����  ���� �����������������������������                        �� �_\�  � � �� �U��pQp��  \ �  UU @  DUUUU��? � �����k�[U[Ul�         �=|�AlelUlU�����������W?��X�� _�}�U���~�_UUPU�W\U�U5UU� =     p p � �          �\;���{0 ��_U @@�@]��?~pp\UEGAU�E�4@� 4 TU�Q��_uUUU     �?|�PEQUEUUUUUUWU|U�� �E�U�U5U��k�  �����kUQA    5 ��>Z�� @    � U�  = � ?    5                                               9 � �         � � l l  [��F��������E��E��F� [  l � �       E kU����        @U����?�@@ 9 9 9 � � � � � � � � � 9 9@@�� >      �� �_\�pQp� �� �U��UU   D�  \ �         @TUUU��?         �=|�A�W?��      ��=���_���� _�}�UU�U5T��U�PU�W\ p p �U� =           �                � \�WU@WU����     �U= �@__��fvj��ZUUEUUUU���QEQD�U�U5UUWU|U�� � � ���U��k� 5 7 �           5 � ?                               9 � ��@�>U� � @        �ZkUE            � � l l [ ��F��F������E��E��F� [  l � �         E kU����        @U����?    @ 9 9 9 � � � � � � � � � 9 9@@�� >                    ��    �  � � �� ��_\�pQp��  \@U��UU   D @TUU �              U��?                       � 0 �             �=                |�A�W?��X�� _�    �����UuT]}�UU�U5TU� = ���p@p    � � p p   G  @@ A@T��pU\t}Gs��=  ut�t��m�[��F�                                    �_�T       �=|�WPQD uAt�@� � ���D�5U�> � = P�Q�D}Q�Gku[��  ��>U�� @  [                                                               9 � ��@@ 9 9 9 �����E��E��F  [ l � �       D VDkU����         @U����? � � � � � � � 9 9@@�� >    �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`L�L��1��� ���������2��3`�1
��4��-�5��.l- H�d���������WWXXDF�Ʃ �<������/ ނ � +� E��1`慥<
��w��-�x��.l- �����QJ[JQ�����XUJJI������)�6��)��)���)����
΅ E�� �`������ E�� �`�<��� �/�L�$ 怩�/�R�$��#��(�/�#��$��}��+ 2��/�#�#�(��`��)�
�� +�L ��+ /��)�+)�3��/)� �<��/�L�$ 怩
�/�R�$ � +���`� �/ ނ�<��)�����)�����ߩ �+ /�� +�� �`���ȩ �+ /�Ά +�� �`��)�
�� �L���+ ��)�(��$)�3��� ��<��/ ނ��/�R�$ 怩�`� �+ �· ���`����� �+ �� ���`VXY�8����+ �����
����� 2�`��̩��+ ���S����(�� 2�`��� ��� �!�/��������"�
��
�"�!���N��/�
iH��!i<�+ 2��/�/��� �/�*�(��J�'�(i �(�
8�'�(�)�*�'��*���'�B��+�M��/
i�� 2��+�O��/
i� 2��/�/�
��` ��� �(�/�8��+�@���D�� 2��/�(�(���`UZXM XYFWY          � 0�� ���� ��`��2�3`慥�)������/�
�(��# ���/���+�R��#� 2��/�#�#�(��`������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������1��&�
�"� i��9�� ���i� ��`�9�� ��1
��=��-�>��.l- ���� �Q�����/���⌃�7�#�YTUXHTWJXYFLJXUJJIGFQQAAAEEEEEJJJJJNNNNNSSSSlnp�����lnprt�����lnprQT\RJI MN�1 ��� ���'�B�U��+�k������ 2��'�'��� �� А��'��#� �"���!�
��
�!�"���'� i<�+�K��#� 2��#�#�'�䭆
m��'��(�p�#�'����+�P��#� 2��'�#�#�(�� ��� �� e���)


�>�����T�

i�=��=� �� 
��h��=��� ������?�8�?�@ c���
�A`888888000000000((  慥�)�`��%@�'m�ee5���'� 
��?�>���+i� � �)���JJJ���'�@� 
�(� 
� 
�(� 
�@�?�>�(� � 2��� �����=��1��i� ��`� �� %��1`�����������:��� �:�;`BBAA@@??d_ZUPKFF慦A���<�#�A���I��9�1��� �:�;���� e�������� e�� �!�" ����i�����!���" ��`����=����N� �!�" �����d���H��H %���������h��h���d8���������б����� �!�" �������К����� �!�" ���Ї����������������������� �����������
�1� ������������ ��`�1` (#	 
#� �/�,�)0�p����


e������������T����	�����E���@���, <��/��/� �+�" ߏ��I����)���� ����� ��L���e,���)��慤A�����[��� ���(��)�	�)�L����W���L�����)�k���g�������'���(�( y�� �L����


e��� ����1��� ���!��������������� ������ ����
� �x�����/����+���" ߏ`�)���)����ޥ��'���(� ���)��)�5��iŃ����' y�� �� <��/��/� �+�" ߏ�'���(��L�������'L닥����'���(�(L닩 �/���-���.���# ����-���.���#����-�!�.�-�4��+ ���8逅�� 2�Lz� ��/�
�1�1�1 *�`�1 ��� ��`慥���	�#��2�`�2�+ ��`�3�+ ����`� �+���� �� �� +�����1���� ����1�� ��`慥�)����� ����


e��� �2��.��)���)��	������	���憩 �+ � 2�惥����Ƅ�����1`� ��/)��� ��� �+�� � �H)���JJJ��� � 2�Ɔh���x�ǩ��`� �/��������� ����#���-���. ��惥�)����愥���ԥ/��18��1 *�`� �� ���1�1`LFRJT[JWXYFWY �������������������IIIILLLLXXXXXOOOOOPPPPPRRRRRSSSSS

�����	�����	��������2�&�' k� ��� �/�ԍ�+������� 2��/�/�!���` ���5)�
��� �+��҅+�O��� �� 2����2�3`XYFLJHQJFWYW^SJ]YXYFWY����̺���ͼ���ξ���������GGGGGIIIIISSSUUUUXXXXXKKKKKLLLLLNNNNNOOOOOQQQQQ�����
��������IKMOQ�����IKMOQ�����IKMOQ���2�&�' k� ��� �/����+�Ŏ��� 2��/�/�/���` ��� m�i� �� ����� k�� �������	��3��2`���̏�H��3��2`� �H���"����H� ���ȏ�����eH�H����� �1`
	DFGIJLMOPRSUVXY[ � 2��"�+����#�#L��$�#8逅#��$�#��$� 2�` ����
i�#���)��#i��#�Ϗ�$��#�`�%��&��+)



e��i ��+JJJJe���-��.  �`� ������ ��� �����`� � �(


e'�� �������� `���� `��%���&` ����'��#�'�i<�+�B��#� 2��#�#�'��` ����'�l�#�'��i<�+�G��#� 2��#�#�'��` ����'��#� �"���!�
��
�!�"���'� i<�+�T��#� 2��#�#�'��`

4  5

�������/��/� �+���4��" ߏ`688  67   6  ���Y�$���#��

�'��(�'�Y��+�$��#� 2��$��#i� 2��(��'�#i��#�$i�$��` 0`��� P ���@�$���#��JJJ�e$�$�Je$�$�)���e#�#��)����$���e#�#�$i �$� �'�'�!�+�$��#� 2��#e��#�$i �$�'�'���`��)������!�����"�������������� ���B�B��� �B�A�A����A`UFZXJ�9I�9� �'�(�/ ����#�(�)��#i��#�Ϗ�$�/� �+�9��+�� �+�#��$� 2��/�'�#�#�')�'���(�(����1��B�9�2� �+�" ߏ� �'�ǅ#�'�d��+�O��#� 2��#�#�#�'�'���`���+���" ߏ`�9��`�.


e-�!��$�-�%��!���������#�	�%�$����-��!���������#��$����$���/�!8�-e%���	�����$���$�.�%��!���������#��%�$�8�����.��!���������#��$�i����$���/�%


e-���	����i��$��`� �����H���+�  � 2�h�����惥����愩 ����`� ��)�)�� ���� �� �������`  (08@HPPPP  @P`p������ 0`x��������:�;��`�;��



e;��Q��'� ��!�����'�
��
�'�#��"� �!u���
��
�������� А���������� ������ ���� ��L��� ��� ��� � �:�����` 戥���I���E�/ ����H��H� ��� ����+� �)���JJJ�� � 2��/�扦����֩ ����h��h��` ��� �/�����+� � � 2��/� � �/�/���惥�)�������`�5)�)��/��I����/��0� �+������� 2��/�/���`�ԍ�+��@�:� � � J�-�@-��� � 
������ ��)�� ��-��I�L핹���	���`��� }T	}!!T!}!T} 	}T �	��  �!T T	}T} }T	}!!T!}!T} 	}T� �� � �!!T  x}	��< }	��<0 <�
<� � �
<�2�   �	� � �	  �} �}1    ����..Th���!h!�AT �@� � \ � � \ B )����!T!�!}!��
<�
<!}  !@!}!T!}�
<�
<!�  !T!�!}!T@	�@	�� 	�}	@	hT	hT}1�  f��2�� a�  �@  	@T	@! �!!@T	�T	�!}  !@!!@!T}	�}	�� 	��	�!}!�!}!T@	�@	�� 	�}	T!.! �!.�	@T	@T	}  �@X � < � < < �0 � � < � < < �0 X � � < � � � � < < < � � X �  � "�  � "�!�!�!�"�"�"�"�#X#X"<#�"�"�"�#X"<"<"�"�"�"�"�"<� � � � "�  "�  #�"�"<"�  ���@@}�} � @@}�} � @@} @@} ����  P\ �  \ � ����!�  ����!�  ��� ��� ����  �A} X!}!@@}�!}!�@@}�!}!�@@}�@@}�!�!�\�  ���"�  ���"�  ��"�� "!�<�    �E��` ����������������������	  @	 	2��!� �!�!}T	h}��� ���  @  [�ћ�T T}T@!@ @T}T!�} }�}T!@T T}�}T T T}T@!@ @T@�	�	}T T�@T}�A�@   ��CX  X�B<  �<B�  ��CX  X�CX  X�C�  ��B<"<"�B�#X  X < X � � � � � < � < � X < � < X < X � � X � � < < < � �  � < #X   ����2��	} !}�!}!�A�@ 	} !}�!}!�A�@ 	T !Th!T!�!}  !�  P  !� �!�!ā�   !� �!.!Ta}  1}T1}T1.T1}�!� �1��a�  1}T1}T1.T1}�!� �1��aT  1T.1T.1.1T1.1.Ta}  !� �1��1�}!.  1T.1`�    < � < � X < � < X < X � � X � � < < < � �  � < #X   ۝y��@T.T}�}T ��}��}T T.T}�}T 	T  L}��T�  � }��T!�  ..T}T. 	.T.T}�}T ..T}T. 	.	�	�	h	T.T0   �@� ( � ( �  �  � ( � ( �  (  J "�  � � � \ � � ( � ( � � \ � � �  �   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������1
����-���.l- ,�{���C�ġYMNS HMJS HTRUFS^� �/�c�# ���[��#��/����+ 2��/�#�#�/����1� �/ N�� �����E���C��D� �G` 8p8��6慥�)�.���/ ����JJJJ)��w��/ ���C�C)��D
�1� �D���C` t�慥�)���Cɏ�
���/ ��Lؠ�i�/ ���C�C�~��C)��E�E��� �/ %�� ���1`Ɏ��!�I�G��F� �/ %���JJJJ)��5��/ ��`��JJJJ)��w��/ ��` #F# 0H`x���إ5)�b慥���[�H�9��/���%��&� �(�*�S�$���#�/�ȥ�+�*
e#��$i � 2��/�(�*�(���*��֩ �*�#i��#�$i�$��`����1�H�	��P��(�/ N�`��H���	���2�3`��3��2� �J`��� !"#$%&'()*+,-./ 123  6789:;<=> @ABC 123  67DE:;JFG @KHI 123  6789:;<�� @A�� 123  67DE:;J�� @K�ߩ �(�* ���S�$���#�/�ꡅ+�*
e#��$i � 2��/�(�*�(���*��֩ �*�#i��#�$i�$��`���%�ۅ&`     	
        !     "    #         ()./4$%*+015&',-236   :987   ;  @   <  A   =>?B  JKTU CDLMVW^EFNOXY_GHPQZ[` IRS\]a   b  f   cdeg                                                               � �(�*�C�#�A�$���%���&�/����+�*
e#��$i � 2��*�/�(�*eD���(�8�'�ѥ(eD�8��(� �*�/eD�/�#i��#�$i�$Ь`   OPQR  UVWXYZ[\]^_`abcdefg    lm          xyz{|}~����������          ���� ������������� ������  ����                                     ��ŷ�  ��  ����ô��������  ����ô�ȷ��ɻ��������                �E�(�*e/�/�C�#�A�$ ���/��+�*
e#��$i � 2��*�/�(�*���(�#�'�ԥ(eE�#��(�E�*�/eE�/�#i��#�$i�$Я`� �(�* ���G�$�F�#�/�}��+�*
e#��$i � 2��/�(�*�(���*��֩ �*�#i��#�$i�$��`�G���S��Fɀ�`��)��0�/ %��Fi0�F�Gi �G�S��Fɀ���/ %��H�	��<���/ N�`� �/ %�`    	
'!%("&# $)*/078+,129:-34;<.56$ =@AH  >BCI ?DEJKFGL MQRYZ NST[\OUV]PWX^ _cdk  `efl aghmbij^ nrsz{ otu|}pvw~qxyL        ��   ������ ����  ���� �����������������������������                        �� �_\�  � � �� �U��pQp��  \ �  UU @  DUUUU��? � �����k�[U[Ul�         �=|�AlelUlU�����������W?��X�� _�}�U���~�_UUPU�W\U�U5UU� =     p p � �          �\;���{0 ��_U @@�@]��?~pp\UEGAU�E�4@� 4 TU�Q��_uUUU     �?|�PEQUEUUUUUUWU|U�� �E�U�U5U��k�  �����kUQA    5 ��>Z�� @    � U�  = � ?    5                                               9 � �         � � l l  [��F��������E��E��F� [  l � �       E kU����        @U����?�@@ 9 9 9 � � � � � � � � � 9 9@@�� >      �� �_\�pQp� �� �U��UU   D�  \ �         @TUUU��?         �=|�A�W?��      ��=���_���� _�}�UU�U5T��U�PU�W\ p p �U� =           �                � \�WU@WU����     �U= �@__��fvj��ZUUEUUUU���QEQD�U�U5UUWU|U�� � � ���U��k� 5 7 �           5 � ?                               9 � ��@�>U� � @        �ZkUE            � � l l [ ��F��F������E��E��F� [  l � �         E kU����        @U����?    @ 9 9 9 � � � � � � � � � 9 9@@�� >                    ��    �  � � �� ��_\�pQp��  \@U��UU   D @TUU �              U��?                       � 0 �             �=                |�A�W?��X�� _�    �����UuT]}�UU�U5TU� = ���p@p    � � p p   G  @@ A@T��pU\t}Gs��=  ut�t��m�[��F�                                    �_�T       �=|�WPQD uAt�@� � ���D�5U�> � = P�Q�D}Q�Gku[��  ��>U�� @  [                                                               9 � ��@@ 9 9 9 �����E��E��F  [ l � �       D VDkU����         @U����? � � � � � � � 9 9@@�� >    �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`�3�r�����!����"�y����%���&� �!�$� ���!�#� ���!�) ���� �/� �!�����)�+LU� ���!�+ ���!��+��, ��� ��/�8�� �$�#i��#��$�#��$���$��8� 
e#����,�� ��L=�`�!��"`������������@  ��()�-�* 

4  5

 -�* � .�,+ � -�* � -�* � .�,+ � -�* � -�* � .�,+ � -�* � -�* � .�,+ � -�* � -�* � /�01 �  !'% � $ � & 	�
 �9@  ������������fgjkno  �������hilmpq �������FI[JSYZWJ�������{������|��}��} XYFLJ��}����
��}����
��}��} XUJJI��}�QT\  RJI  MN  �}��}�R^ KWNJSI��}�MFUU^ RTWSNSL �}�SFZLMY^ LZ^��}��~���@                       !"+,56@A   	#$-.79BCKL 
%&/0:;DEMN  '(12<=FGOP   )*34>?HIQR                     �J  uv���wx���yz����{|�����k}~������l�������V WXXY  mn�������  Z\]`adehiop���������[^_bcfgj qr�����������st�����������@  ������8�
�						@  �	�
�q%34GH[\�&'56IJ]^�()78KL_a��	*9:MNbcs  �	+;<OPdet  �	,=>QRfmu  �	-?@SThiu  �	.ABUVjkw�/0CDWXl� 12EFYZno�*@    ��z } }z z}  zz�����{|~|~{|{~||{{��  � q	 #q	 x �  � r
 $r
 y �  ���������������  �� � � � �����������������������������������������������������������������������������������Q@  �	E\]qr�������	F^_st�������+,G e`uv�������-.I�wx�������/0K�y�������12MNabz{������34OPcd|}������56QRHf~���� 78STJg������	!"9:UVLh������
#$;<WXij�����%&=>YZkl�����'(?@[ mn��)AB  op�*CD�p 
  
�%��&��+)



e��i ��+JJJJe���-��. ��`��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������1
����-���.l- ?�(�`�XYFLJ >AXUJJIQT\RJIMN YW^FQQ XYFLJ HQJFW�J
��P��-�Q��.l- ^�����Ő���� �I��K�����J�G���F�1`�F�G��F�1`��I��K�����M�٩I������
�M�G���F��I�G��F��K������I�1`������K��I�R�G�d�F�1`��I��K�Y�G���F�1`������I��K�T�G���F�1`�1�1`������I��K�T�G���F�1`慥�)�,����%���&�I���+�F��G� ���F�F�I�K��1�J`����2���]��3� �J�K��`�1
�����-����.l- ���H���INWJHYTWFSI^ HMJSUQFSSJWQNS HMNS SFSFWY^FSL \FS LZFSLUWTLWFRRJWRZXNHFR^ HMTZXTZSI JKKJHYYJ]YHFWTQNSJ XMNMUWTIZHJ G^YMNS HMJS HTRUFS^=EE>�K��)������K�1�K��� �K�J�J��`�1�1`����i�/�
�(�W�$�J�# ���s�/��(�Y�$���# �����/��(�[�$�Ѕ# ��� ��1`�0��
��` $5?LX
'D\			��9� ��8��J����/����(�X�$��# ���J����/����(�[�$����# ���1`23 ��%���&�/�����+�K�����+�#��$� ���(��/�#�#��`                    �<<<    <<<�        �<<<<<<<<<<�        <<?<?<�<�<�???<<<        �<<<  �><<<<�3        �<<<<<��<<        ��<<<<<<�?<<<        �?�����������        <<<<<<<<<<<�                   �?      �������������        �<<< � < <<<<�         ������ � 0   < <      ��u|��G[�����s���s����G[��|t�] ���pp\\��UU            UU��pp\\��    �<<<<<�            � ��k�V�U����    �<<<<��?<<<<�        <<<<</>������                     ?���Gp|t�\p  �W5G���4T44p�  \ �      �� 4 5U5p��A�ApG\���U� � � � � � � � � � � � �                     � � �          U���p�\��o           � ��k l [<[�V�V�[�Y�V�VkUVUUUUUUU�����VUVUYUUU�U�����         � p \ W   ��o|UWUUU�U�W W����supu\u\U\�W]U]UuUuUuU����v\�l��[��pl _ Z!��8�     �pp������Q@p�    �pQ��U  @ �� mp�  l l ��P�_�U�@� � � @��n۾��V^V9[�l�    k�V������U�Z[�VUVUUUUUUU�n�[�[�[�n������UUUUUUU�U�U�U�U�:�:����� l lU:U:�:���:�:� l [ [ [�Z�j����  �U>U�UUUUU�UW ����Vo��U�W��U�UuUuU]U�U�o��]�]�uUuUuUuUUUVUA��Q�0�oU�U�V�[@n � � ������P } � � � @ @      @��v�}m|��               �|u_u_}WmWW�   d � � � � 9�T  @ �U骿�j�V@�� > � ����Un�Y�U�U���U�V�������������V�V�V�U�U�U�U�U��������?    U�U�UiUVUUUU����� �?��U�UUUU���� � �P: �A�Q_D            9 �E��_�����9 � � ��UUU��U�U�U�U�U�V�V�  ��  ��  ��  ���� ;       [�[�n�nչ����U�V��pp\\��W�����V�V������:�:���� ?�?���P@ �/�,���  ��  ��  ��  ����p@ \���� 9 � � � � � 4 �?W���p�\��    UU��pp\\��?             �� � ? ?         � ��:���?                                    �?    �     �?    � ��?4�3�4�8�P3�4�8�P3�4�8�P3�4�8�P3�4�80000000000000000��3�4�=�7p3\�      <<<<<<<<<<<<<<<<  <<<<               @���,tt8p=��    @���,ut�      @ ��t48,p� �        �6p�,��@    �|,84��@                ��8�4p4p4p�,��@@        @ @ @ � � �  s � ��A  � ��o��w =      , t � �        U�[� 4 � @  4 � � ���   �� 9 � 4 @� ��@U            ? 9 4 4@4�4t      4���W�} 4t�P                                     � �48l�            @��  @�? ��p  �� � p ��,  p �  p�V        l l  ����               � ��y���@� � � P�    l l l � � � � � �     �             �9 ��������� � 0p�pа��A�B � � � 0 �������� o  G  l p � �U� ��� �T���=A �              �?        � � �                                     � � � ��뼖       � � � � � � ��k�VjUVU����kUVUUTQQ@UU����     ����ZkVTQ    ����UUUEQ@T QDT Q D  D@PUEUTEUEUUTEU @  @  �@�Ы��TUQD�����������^�G������oo����������[��P�WP����ZZU��  �����ZZ U�o ��C�^�����������������������9 ��VU    �� \��P^ � � P l l �Q����n�o  @��E�_}��_[n[mnm�m�nU�V�[�U�����չu����:�:n�i��fU�UiU������������:�?      ? � �@ 9                 9� �� �@A           9 U U�o����������9 9 � � � ��������o[W�����Z���VE@[����j�t��F  @U����       UU��  �� :�6��|���|�����������������>��m���U�kZ  �? ��U��  � ~�~@�U��m  P��Z^U�U��[Q�T�U�U��o�� �]�W�V�W�]�U��k�[ � � � l � k�����Z�V�UfUYUVU������U� �U���   : � � ��E_� 3�?s9p9������� � � � �@n� > �Q99 @�G����u����Ζ�A�� dt?p<��6�:��������l�           ��W�UETPUU���� � �����������       > � � �                    � � ��������������������/�������������� � � ���                            ? ? � � ����;�98�0�p��� � � � � � � � �       � 0 p �                           � � � � � � � � � � � �                             ����������       / ? � � ����?��ӑ�G�]9�yC���<��� � � �                   � ����           ����������������������[�E�����o� �l�U��V�V�Z �𯿮DG�����몪꪿���l  ���V[@�� � � � ���������F � @ @          �l   WU��kl  �@        l�/�?�� � ��     Po�������/�?���� � ��Z�UlU\m[[�[�V�V � � � �        �V�V�V�V�V�W[[l[�[�[ � � � � | | p �                    �����        � ��>�;���������������������[oA �[       > � � � p , \@��o�����[on�����[o�ef���o�UV     �����                �����P   �      ������є�� ������P/Pj@            @� � � @U ��j��   �U        U�U�UU�ZU�U�U�U�VU����9 9 : ?��WU�U~��]uU�E�m}WD     @   D�WEF%�P @   P �@4D� 9   �V�                                          � � ���������� <                  � � x � @                              9 9       n �? 9 ���������? ���������   �[=U�� D   @o     ���9�䰐o��п�������������oAnFny������п��@o      ��� � � � � �                 � � � � � y@n@         @ �@�>��_���V������S�?            ������         4 5 4 5           � �મj�Z   ���������Y�U��Z�j���������갺U�U����������������ejUoU�W �        � � k��   ����_=��PU�_l@��48� �p �������/����������       ���            4 �M�,Ь�z<=��P        ��kz�9��PGS�C�   V �U����OU�U�s 0 � �@�����U�D�T��C�S���������� � � �G}?���� � � � @        �������  ����j�Z�V�����������Z���o������j�������U�U�V�Z�j�j�������������������������j�j�Z�j�j�j����U�U��� � � � � � �    ꪺ��������                      ���U� T          � �P: �   @ @ � � t��[NxUu�� ��<| } � � � � � � <|?�?�VG�E�l  � P                                                @ @ � �     TU����WUU @y�^�   � [�lW�U0��? �~��<0�                      ���������U�U��Y������������j����U��������ꪺ������꯾������j�j���UuU]UW�V�Z�j����j�����������������j�Z�Z�j�j�����j�Z�Z�j������� � �            ���������������              �                �9n5[�WՖ�U�U�u6          ����[}��U�_n�[U�A~@�@�V}[_�_�5������;@@@�@�@n��ϐso�����1�?:�9 �p�\9\9���^�009           �5��l�\1W0�                 � 0                              ����U�����     ����������������U�U�����Z�V������ꪺ��j�Z�ڪz�������]�[�U�U�U�Z������������Z�V�U�V�����������Z�V�U�U������������V���U�U�V�Z�j�������� � � � �����p9��������ê � � �p9\\��� � 9  �              9                                              � � l [�����    : >     ����~�뵪�������   � �����[ZVVUZUj����������n��������ڪ֪֪���������eUUUUU�ڪꪺ����������UUUUUUU�U�U�V���������j�Z�Z�j��������ꪺ����e�����jUjU��������U�W�W�� <       ���������� � �  ���@T T@ T @ } � < } }T@ } T � T  T T@ T @ � @ �  T@ }@T � }0 �� ��� � � � �  � ��� � � � � � � ��� � � � �  � ���� ����p   �@#X"<"�"<< � � � < � } � X � < � X < � < � � X � � < � � X � 
< 
< 	� 	� �  T   @ } �  � � � � T  T �  T  � @ � @ T  } @ !T!A�  ����@2<�!T!�!}!T!@  2<�!}!�!�!}!T  1�}!T!�!@!@�  \!T�!@T�}T}������ !T�!@}�a�    �@X � < � � X �0 � � < � � � X0 � < X � � � CX  |� < � X < � < "� � X < � � < X0   ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L����ϓۓ�/��                ��?���������?��l6��g��g�9��0����0���?�?���?�?��l6��p��l�9�  <<������<<   ?���l�k��[����}k�k�k�k�k�k�y��[��k�lѬ��� ��?��W�@W�������_���G9�:�� � ��:G9��[��?�����������������������U��������������UU����������������j *U*�+	������������������������ککک�Uکک��?�������U���U��������_����_��U���?|��s����V���:�:����?�絛����������ꪪ�������U��U���������V�����W�g�g��Z�3 ��0 �0� <� �  0 ���3�: � ����������  � ����������������������몪����     ���_?|��s���_V������������ ���?�<�̿������������������̰���������������� ���W | � ���������  UU��  �������� �U�j�`�`�`�`�`�`�`�`�`�j��@���@��j�`���UU  ��  UU��  ?	?	?	?	?	?	?	?	?�?U� ��� ?U?�?	?�?U? ��������UU  ����������j��@�����������P�R  �RP@@@ TP @@< �W>�W�~�} <���[�kս���@}          �����l4�l4�l4�l4� � 0� � 0�������UU��UU������?��?����?�  �?����<<�?��  �?????�  �������  �????��< �?  �????�????�  �?????????�? ?  �?? � ?????�  �??? �????�  �? ? ?����  �????�????�  �????�? ???�  �<<<�?<<  �<<�<<�  �<   <�  �<<<�  �?  �  �?  �?  �     �< �?<<�?  <<<�?<<<  �������  �?   �  <��?<0        �?  <??�<�<�<�<<  <<?<�<?<0  �<<<<<�  �<<<�    �<<�<?<�3  �<<<�?<  �< � <<�  �?������  <<<<<<�  <<<<<<�  <�<�<�<�<�<<  <<��<<0  <<<����  �? < �� < �?��
�*�*�*�*�
��
*(�*�"�*�*�*�
�*�*�** * �*�*�*�*�*�*������
*(�*�"�*�*�*�
�
�*�*�*�
*****( � l      ? ���W���A�A�A �\  pU���A�A�A�A��W� ��lU@ 9 4 4 4 ��P� �@Us���t�t�t�t�t�����        � U�AU@              AAAAAUW��         ���������,< 3�0000�03<�?�����0� 00� 0 0     <  � ���0�033?3�0�����33�0000�0?0� �00����0 0 ��00�?�         � \ \ �   ��۰�t�lŬ���l�l�l�l�l�l�l�l����l�t���� �    ����UU  UU��������UU  UU����     �SC9W:�?99999999�?49K[�            � C� ��   � 0             ��WpU\U\U\U\�p�z�z    �pL�1p| ��@�@  � � W�W_^UUUUU��� � ���U�UUUUU������@  ������ �  � T         �]P������ � ���W��   ��UlD[D  ? ��:D��DDQ�j������U�UUUUV�DD*���������U�V��U��@U      [U[UU�U���� �    @ � � � �� �@@~@�|  @ �U���@��?�?��?�����k � � l W WUW���7���}�}U_U_U��   � ��
����         : � � �������ο��?� : :          �� = 4 4 4                         � ���              � �������� f � f � ������ � � � � �������          ������ � � � � � � � � � � �                          � ���������ff��ff�������� � � � ] ���]    UU��������������UU��?/|||�p����=�= ������UU�������UU���������������������������������������?��������?����������������������������������                       � � , ���     � p p p �  |UWUUUUUU��Wz ����<��     � �0�@ �                 p ��p~������     � | �PU    ����[�U���UU@U      ��[�ED�F��       9 5 � � U�UUUUUU��U��Q�� � UU�U�[������C �?�?_:��� ���@�@�@���WW\�P�����n���4�=|=>?/����n�ne�U��UU  ����?            ������4 4 ? /   < � � � ?                                                  � �  �0�3 < �                   � �� 0p�} � W     � | � � � �   ��޷z � � � � �      �z������_�T� �     ��VlU[U[��W_ � |��kU�[�}U�W  <��p��5? ��@]t�@��@ @@}���� � � ��M_5  �A�A�Au 4 �W�]�U�U�׵T    5U�V��Z�UP     �QD45F��mԹѵ����6�6�W[]]]]_m�� �=�|��?A                                                                                                                                    UU��      UU� p�p�s�s�s, �?��� ��UUpppp p p�UU  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ���?�?��    ��h)h)��    ��((((��  ������0000�0�0                UUUUUUUUUUUUUUUUUUUUUUUUU ���V�F�� [ � � �                n����jP ZU���� ������������S�����������T��[999999yyyyyyyy99A-P�� /   K�Ŀ���������������������������UAU���[���ll@n@����n@l@l ����[��U��������������� ��������������_�o��U�P    P��[l����l�[�P    PU�����T�S�O�/�?�������������? /     PUCU.U�T�P�S�KPN@@.999A9@.@P�K�C�R�P.TUPU����/�/�?�?�����������?�?���[999999��iQ��999999[9���?�?�?�?�?������ � � � � �UUUUUUUUUUUUUU�W             � ��:U� PU ��  lPmCmm9myl�l�l�l l l l l l l � ��l�l�l�l�l�l:���?�������? ��?�����?�?�����?� �?�������?������������UUUUUUUUUUUU_Uz�               媐UP  T@�P��� �U�^@y��[�l���� � � � � � :  �������������� ?������������������������?�?�?�������� �?�?�?�?�?�?�?�UUUUUUUUUUUUUUUU      �\�WUWU��          � ���l  ��  ��  ��  ���W��u�u��<, ��?�C3TOUSUPUPU p�p��� _��p�?��������������0?������������������������ � � ������������?�?�U��]W��U�_� < �  4555�WP� [����� �y�{_}uu��@W@^@~  ? � � <@ �U���@~@~�ה��>�;��?���������?�?�?������������������������?�?�?�?�?�����������������  UU����             � ������_������_�W}UU�p�^�W\�\\�WW                ���������������?U�T�T�T?U UU?U���������������?    ? � � � ?                                   ��  ��  ��  ���?�����������?���������??????�? ???��??????��� �?  ����� ���? � � � �����       �� � ? ?��  ���������������������      ����������        ����� � � � �  ��������� � ������      �����        ����� � � ����  ���?�?������� � � ����      �����       ��3�3�3�3�3�3��� ���3�������               � � \ G �E�pDp\DGD ����Vl    ~D�Q��@�@n � �  [ [oE�V���� � �@���䫹Vn ��k�������k�VT       n��[k�V��nn �V꫕>U�P�@� � �          �� < ��������<��������� �0���������������������A< � � � � �   � 0�C��|�|�  ��0� � 3 3 <�M�M\��u�� ���Am��4 � ��Ъt�]�Wt5@]�uu�Q^DQ]DGMD}�D�QODQGQGTWUן�����k�@���Z�UUV�[�n��n  V k��V�[@n�n�����o�n�@� � � � �@�@������꫻�n�[������U[      ����[�o@�@�@�0�0?������������???�?�?�?�?���_����1�1}��?�?�����0� ��������0 0 � � p������??��������3�3�1T �W�S������p���������������W�~����_\A_��_��o�����������������z�z�z�z����������������Z�P  ������������              P���k�����nZ����讀TUPA @  oU����뺮o���     @�U�֫�Vn������n麔� � ��� �U��4 444p44�u~]         5 � @���]Wu�t��������UmU[DEDWDQ��ֵ�m���E_]E\^Dz�EUUDD�E\E\O�����ѫ�Vm[�_��Z�P�o�n@� � � � �T�          �����V�� @ @  [PZ����﫺n��n�n       @ @�V�������Unn[ VV    � UQ�D��D�9D99DQT��� � �@@A9W9^:�����V�V�V�V�U�j   : ������@�A��k�@    F��o�o�[�[�[�k�� _ z��W��@�@��됛�V�����Z�P         ���Z�T      VT 9 9 � � � � 9 [�n����Z�n_^U:  � �P 9 9 �                ����V���V��F�F�R�F�����F�F����������U�E��Q�D����D�U��D��P�A�����A�Q�Q�����VU&VPFFDFDQQFPFFFAAFF��k][[]��[U@@[U��[][����U���U��WU@@WU��Uu t tUu�� ����V����V �����UU      UU��           ��V`A`U�Z �               � j�e      ��VY       QVE�U �      DUe�U�U Z �      
�%Z�@       
 % �@� d@T TUU�X
�   A  TU��*)              * �P	 %U	�
                                  � p  G      ��_UUD         ? � @                          � � p p�\_GwGבW�_���D A_U��UUUU_U@�P_�UU��     4 4 � �  p p p p � �    ���ꐪ@��P |���������ZU    ��Z       @ �� � � � 4 4          ?��pp]���W��{��U�4|��  UU����UU@_���P��믶V-Q�s���   �@0�5?                       � | �Ep    ��_UEDDDQ         4 5                                 pE\\EpUp������_D�Q������_UW�U�� ���UWUU��u�P   � UU� � 7          � � �   W�U|�W�UmU[UW_�Z�U[      P \4�Q@    4 4 4 5                 �G  \ p �         t�W��� �  ������_��           � ���UWUU��[�@   � UU� � } @@@�t}�P� 0� � =  4 4    A@� =  P��               �Z�U[       D @G��}|��<                                                  � �����k�[U[Ul�  �\;���{0 ��_U @@�@]��?� U�  = � ?                                  �         �=|�AlelUlU����������~pp\UEGAU�E�4@� 4  5                    �� �_\�  � � �� �U���W?��X�� _�}�U���~�_UUPU�W\TU�Q��_uUUU     �?|�PEQ           pQp��  \ �  UU @  DUUUU��?U�U5UU� =     p p � �        UEUUUUUUWU|U�� �E�U�U5U��k�                                                                                  � �            5 7                                                                                                                                                                     �  � �   �=|�A�W?��      ��=���_��  � \�WU@WU����     �U= �@__           5 �   �� �_\�pQp� �� �U��UU   D�� _�}�UU�U5T��U�PU�W\ p p ���fvj��ZUUEUUUU���QEQD�U�U5?           �  \ �         @TUUU��?      U� =           �              UUWU|U�� � � �  U��k� 5 7                                                                                                                                                                               �=                                                                            ��    �  � � �� �|�A�W?��X�� _�    �����UuT]    �_�T       �=|�WPQD           �_\�pQp��  \@U��UU   D @TUU}�UU�U5TU� = ���p@p   uAt�@� � ���D�5U�> � =                  �              U��?              � � p p   G  @@ A@T�P�Q�D}Q�Gu�                                                          � 0 ��pU\t}Gs��=  ut�t�                                            � � l l ����k��� } t ��>U��@           9 � �  [��F���� � � � d   � @               �@@ 9 9 9 � ����E��E��F@ � }   d d                � � � � � � � 9� [  l � �       E kU����        @U����? 9@@�� >     ����ZkEE    ��>P� � @     �����k��E�� � � � � � t } @ ��>_��@                ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��P4�QO�����_��    4 4 4 5            @@@�t}�<�����V��  0P5�  � � =  4 4                                   ��pUp@p@p@���� ��k ��UUU��?T�� �@��WUUU�UG^�  p \      U�1t t��@�@3@3�UL ���� 5 4 � � � 4 5  p � |  ����< ��W������ZW[\�sE_�V��_�����1�   � O|�? � � [=�l�l�l@��� k � �  ��]�� ��ZU����T 0}���U������ t@���_}jU��w�P  TT���� � � �����W�99A9@P�� >    ? ��?�������������� � � � � � ��~p�0�0�0p�_ \�s]�4 4�ZU���� ���<0 ����� �0<����< �_���C10001 �T�C0L@@@ L?p�@U��������]���pU���o�_�_����m��mU�����~��z���^}jU�� ������������������� ? � �0��7��7�53�07�t�P  TT����? �������?�?��?               ��������������� � �                 � _�p p \     = � @� ���Mw��<          ]n�n     ������^�   �]t t�ZU���� � ��Z�[     � �P: � � @ @   � \� ��_�_   u�_ ���@��_P� T} ��}@� � �UU| �<G�G   � mm}�VU����� t tA��^}jU��     � | �~ n     � P   4�u��� � � � � �q7��<3          ������ � � � � �����W�99               < � � � p �             � ��w��    � ��S0 � < �@�?�ꫪ��������������������W�\�p������^�~�^�z�ꪪ���Up p   9 9 ��������@z@z@z@z� � � ��UU�����@z@�P���]}jU��   > � ������U?�5�ک������?�?�?w�� ����]t t�ZU����s�P  TT����   �   �           � p p p � �   � W  \ � �   ?��]�t 4�ZU����?��_�0s s�|�|�U��Wpp���_Uu!P0      ��p�T@@P_|�W��?�0:�����=���ʬ��°���j�A�VU������w�T��]}jU��       4 5�5\          ? � � 5�A�A�����ս5�7=             _==P7�5mF��P  TT����  � �<�<�0�  � p   p p �                      �]4 4�ZU���� ��[lE�ku���y��U��@} �pW|�t�� t ?w�W��|]mU � �PW��Ѱ��A�A�A�@�P����^��m������ќ��|��U����A_AG����_}jU��     9 5 5 � � � � 7 9 ? =��20�4�KO�          ������ � ��[|�0�@ , p��7 ? 3 � � � ��3]� 4�ZU���� ��Vo�������� �P���������P���׿E� �  ��Po?�?���   �?������0�0000<0��< ��<��0�� �<�<U�������0���\}jU��      �����o3        �< 0 � � ����0����<      ��0� 3������]4 4�ZU�������<??L�ZK�    4 4 = ; � s ǿ �C��[��[�� � � = � �l?���j|U�AUW�����ꯗ����^}jU��     �:��^�y��?s�P  TT����       � � � � � � 0 � � � �   p �    0 � \�]}� 4�ZU����  0 ��G[l � 0     = � @�P��s�<<0?��@����LO ��p]s�|<|<�7W�@   �|p|plp\     |�UU���� ` `PA��]}jU��                        �[�u 4 4 8     �  < � ����:�1             � �����������@� � � p �����4:W?�K۫[���l�l������3>|�<>�?]�� 4�ZU����     ��_|� �    ? �@����V�@������P���37??T  �}������@�  P��    @��o����U������������\}jU��       5��\]��}            �]���@@@>O�sw           ��1���5�9 �s�P  TT����xآ��� � ���& �� �� �� �������� �7� ������������������ �2���  � � � �  �� _���2� �3���  � � � �  ����L]�����e-e.ee�� ���2����(���&  ��  ��3�Y��& ���`�� ��� �1�2L���3� �LL���  �LL���  �LL���  �LL���  �LL� {��2��� �2L�􉉉����		
� �g����� ��`� ��m���)��������� ��)�� ����I�L��������`� � �������-���.� ��� ��`�i0���`� � � �* ����� ����`�  I����I�%��`���`�� ��`H�H�H�2�
 � *���2�5�� �� 	�h�h�h(@���& ��� ��� � � �* ���  :�����[��� �����5����& �5Ť���� �� d������쥣����5i<�5��`���Ơ`栥��>�]�:��8� Q��i0���i ����������������i0�����i ����㥢���  	����a�.�]�*�D Q�����ȑ���� ��i0��i ������� ���_��a�Ș �����a�����`�`���ơ`���K�]�G��8� Q��i��i ��i0���i ����������������i0�����i ����㥣��� 	����a�0�]�,�D Q���ȱ����'��� ��i0��i ���ߩ�����a�����`�`



}�������i ���J��� Q����e��i �������`� � ��@�� ��������`H)��l��hJJJJ�
ei@}|��` 0`��� P���@p��      

�� ���� � �����`� �/ ����� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                  ����	��ȱ	�� �����0����J��� ����� �* ���`��� �c�� �  �ޥ
�����	����
`� ��� �������
����`
�����	����
�
��	�ȱ	���� ���� ��L� \�L� <�� 0]���JJJ���� ���Bȱ�3�

��3� �)�6� �� �!JJJJ�$�)pJJJJ	�0 ��� � 	�`��-�>�����k�Ls��*��$8�'�$���)�* �� �`� �-�$ �� �`�*���'}$�$����)�* �� �`�-�� 	� �� �`�*�Ž$8�'�$��!)�$L+��!)�$���ǽ)�* �� �`�*� �� �`����)���0��)pJJJJ	�0�

��)�%�38��3��6� �3�6�3� �6� `�3e�3���6�6��ީ�6���3�ҥ�

��)�JJ$	J� `�����-`
ee������)�*�JJJJ�'��-`�����e`���ȱ������.�@���*��� �c�� �  `��ý	��	��L<���ȱ��	�L<���ȱ�L<�
qe�����ȱ���L<��05

�������� � �����)� � ����� � ���� � ���c��S)x�OJJ�����C��?�0&�8���
�� ���� � �� � L^��e�������ܩ ���� � � �0

��������( ����) �����* ��	��� �* `�oU \ :y|I)O1 o�y� �, ��ߗ�ߙ��ߚ#�՝U������������ ����.}.�.�@�   �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������9�S�S�