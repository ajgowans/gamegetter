                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �� ���             ������           �_U��_UU�      ��    |UUUUU5          �UUUUUUUU  ���WU�����WUUUUU�          pUUUUUUUUU���UUUUUUUUUUUUUUUU         \UUUUUUUUUUUUUUUUUUUUUUUUUUUUU         WUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        \UU�_UU�U���W�UU�_U�UU�U��UU        \U���_��W���W��U��U�UU��U��WU        \U���_��_���W��W����U��W�����_U        \����W��_�WUU��W���W��_���_�_U        \�������_�UUU��_�W��W������_�_�
        \UU�W���_�UUU�_�U��W�����W�_�        \UU�U��_�UU��_�U��W�U�_��W�W�        �U��U�_�_����_�_�W�W�U�W��_�U�          W�U�W�_������_�_U�W�U�W��UU-         �U�U�W�W������_�U�W�U�U�U�UU-         �U�_U���W������_��U�W�U��U�UU�         pU�_U���U�UU�_�_U�W�WU���UU�         pU�WU��U�UU�_�_U�W�W��_�UU�         pU�WU��U�UU�_�_U�W�U���_UU�         pU�U�U�_�UU�W�_U�W����_���WUU�         p��U�_U������W����W����_U����U�         p�U�WU������W����U����WU����ի         �UUU�UUU�����WU��U��_�UU�����*         �UUUUUUUUUUUUUUUUUUUUUUUUUUUU�          WUUUUUUUUUUUUUUUUUUUUUU�����+           \UUUUUUUUUUUUUUUUUUUU�������*           \UU��_UUUUUUUUUUUU����������
           \UU5 l����_UUUUU�������
                \UU5 �5 � �U��������                  pUU5 �6 � ��� ��*                     pUU5 �: � ��� ������                pU�? �: � ��� + ;   ����            ��� �: � ��� � ;   �   ��?          ��� �: � ��� � ;   �   ; �          �
 �: � ��� � ;   �   ;               �: � ��� � ;   �   ;               �: � ��� � ;   � ��;�             �: � ��� � ;   � ��:�             �: � ��� � �� �� ��;�             �: � ��� � �� ��   ;�           � ��: � ���   �� ��   ;�           � ��: � ���   �� ��   ;�           � ��: � ���   �� ��   ;             � ��: � ���    �� �� ��;             0 ��? � ���    �� �� ��:             0     � ���    �� �� ��;�           0     � ���    �� ��   ;�           0     � ���    �� ��   ;�                � ���   �� ��   ;�                � ���   �� ��   ;�                � ���   �� �����;�                � ��� ;  �����������                � ��� ;  �꿪�������             � � ��� �  �����������             � � �� � � �����������             �� � �? � � �����������             �� �    � �������������?           �  �� �    � �����������             �  �� �    ���������?                 �  �� �    ������U��                  �  �� �   �����_U]                   0  �� �  𫪪�WU�                   0  �� ��  �����UU0                   0  �� ������� pUU��                   0 ��� ������  pU�X�                    ��� ����:    \U�X�                    ��� ����    \Uը�  ��?               �������     \��0  ��>               �������      �? �?  ��{               �������       � 3  ��{              ������       ���  �{	              �����?        ��� ��O	             �����            ���SA	            ������:        
  �?0< �PI	            ������        * �?�?��<PI	                          �. <� � 03PI	                          �� ��?   TI	                          ��� � �?TB	                          ����    � TB                          ��00  �� TR                          �2�  <� ��                        �* ��2� �   ��                        �� ���> <   @%�                        ��
������   @%$                         ������?��   P	%                         �> ����/   T		                         ��  ��*   UB	                         �   ���  @�P                             ��   P%�                           : 00  �   U	%                          �:�   �+  T�B	                         ��?   �
  T)T                        ��� �? �* @�B�                        ��   � ��
  U
                        ��� ��
�< �+TU�                          ��?����; �� �                           �:�j�:�*                               8 ���:�
                                : �V��                                 > ����                                ���� �                               ��? �?��*                               ��:   ��*                               ��:   �                                �
8��+                                   8��/                                   8��>,                                   8+ �,                                   � �/                                   �
 �/                                   � �.                                   �   *                                                                                                                                                                                         �                                      0 �?��� ��?�?������                   �� ���� ��������                    3� ���� ��������                    3� �?�� ��?��������?                   3� ���� ���� ����                    �� ���� ��0�� ���                    0 �?��� �������?��                   �                                                                                                                                                                                                             ?  ?  ?                               �� �� ��                               �� ��  �                                �  �  0                                �  �                                  0  0                                ?     ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �  �5 ��� p�U\�U\�UW�e5���5W�e5W�U5W�U5W�U5W�U5W�U5���?  0       ��    ��  � ���+���o����_��[�>��� �� ��     ���* 8�BU9�BU�RUN�R�N�R������~9D�B9T�R9U�R>U�RU�CU�N�����? �� �����?�>�Z���U��o���k���k��������������?���?��������?     � �      (     �  �         
    �       �    �     �
 �                                                                   �?  �� ��V��V��V ��  �� ���pW�p]u=|�_2�V���j��W�ë�?0�� �?  �� ��V��V��V ��  �� ���pW�|]u��_=�V�2�j�W�?������ �?  �� ��W�5\�?� ��  w� �7�p�|�v��_=�V�2�jç�?������ �?  �� ��W�5\�?� ��  w� �7�p�p�v=|�_2�V���j����ë�?0�� �?  W� �U%�U%�U� ��  ��  ��  �� ��� pY? �V� ?�*�U���� � �?  W� �U%�U%�U� ��  ��  ��  ��  �� �Y? �}5 ��:  _5  ��  ��  �?  W� �XU�XU��U W�  s�  s�  S?  [�  �e \} �� \�  �?  �?  �?  W� �XU�XU��U W�  s�  s�  S?  [� �e _�����WU����� �     �   ����<0?� �     � ��0�?�ڿ]�՟]�՟����y�?�z5�?�UUUUUUUUUUUUUUUU ���uU\�U\U�W_7 W�5 W]5 W]5 W]5 W� |U ��                   �� ������w��w�?|w�=|UU=\}}5\�5WUU�wUU����\UU����?�5���   �� ������w��w�?|w�=|UU=\}}5\�5WUU�W�����Wp5����?\  ��00��00�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���*      �?�?                                                                                                                                      @0   PpPP  � ��0000 p ��    	    	 	%% 	  00 %05@EP                                                                                                                                  H�Z�z � �Lܠ�� �Lܠ�w �Lܠ���� Lb����� Lb����� Lb����� Lb���� Lb��� �� �� �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� ί �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� ί �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� ί �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� ί �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� ί �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� ί �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� ί �Lܠ�� �� �� �� �� ��  ࠭� �� �� �� �� �� z�h`H�Z�� � �L��� c�L��� ��L� �z�h`H�Z�� �� �� �� �  㫭� ��0L<� ū�� ��0��r L_��� �� �� �� Ι  㫭� ��0Lr� ū�� ��0��r L_��� �� �� �� Κ  㫭� ��0L�� ū�� ��0��r L_��� �� �� �� �  㫭� ��0Lޡ ū�� ��0��r L_��� �� �� �� �  ū�� �� k�L_��� �� �� �� Κ  ū�� �� ��L_��� �� �� �� �  ū�� �� ��L_��� �� �� �� Ι  ū�� �� ��z�h`H�Z�� �� �� �� �  㫭� ��0L�� ū�� ��0��r L���� �� �� �� Ι  㫭� ��0Lʢ ū�� ��0��r L���� �� �� �� Κ  㫭� ��0L � ū�� ��0��r L���� �� �� �� �  㫭� ��0L6� ū�� ��0��r L���� �� �� �� Ι  ū�� �� ��L���� �� �� �� Κ  ū�� �� ��L���� �� �� �� �  ū�� �� ��L���� �� �� �� �  ū�� �� k�z�h`H�Z�� �� �� �� �  㫭� ��0L� ū�� ��0��r L��� �� �� �� Ι  㫭� ��0L"� ū�� ��0��r L��� �� �� �� Κ  㫭� ��0LX� ū�� ��0��r L��� �� �� �� �  㫭� ��0L�� ū�� ��0��r L��� �� �� �� Κ  ū�� �� ��L��� �� �� �� �  ū�� �� k�L��� �� �� �� Ι  ū�� �� ��L��� �� �� �� �  ū�� �� ��z�h`H�Z�� �� �� �� �  㫭� ��0LD� ū�� ��0��r Lg��� �� �� �� Ι  㫭� ��0Lz� ū�� ��0��r Lg��� �� �� �� Κ  㫭� ��0L�� ū�� ��0��r Lg��� �� �� �� �  㫭� ��0L� ū�� ��0��r Lg��� �� �� �� �  ū�� �� ��Lg��� �� �� �� �  ū�� �� k�Lg��� �� �� �� Ι  ū�� �� ��Lg��� �� �� �� Κ  ū�� �� ��z�h`H�Z b���� �� �� �� �� ���  �� ���  ��� ͜ 0W͝ R�� ͞ 0J͟ E�� ͜ � �L��� ͝ � ?�L� 䪩��  ��� ���  �� ��� ���  ��ή �߭� ͜ 0͝ �� ͞ 0͟ 	 � ��L�� z�h`H�Z 䪜� ���  � Ͻ �� �� ��z�h`H�Z 䪩$�� ���  �� �� 7�� �� ک$��  �����  �� �� ک$��  �����  ��$��  ��z�h`H�Z b���� �� �� �� �� ���  �Ι ���  ��� ͜ 0W͝ R�� ͞ 0J͟ E�� ͜ � @�L9��� ͝ � j�L9� 䪩��  ��Ϊ ���  �� ��Ϊ ���  ��ή �߭� ͜ 0͝ �� ͞ 0͟  � ��ΰ z�h`H�Z 䪜� ���  �� �� �� �� Ͻ �� � ��z�h`H�Z 䪩'�� ���  �Ϊ  �Ϊ  7�Ϊ  �� ��z�h`H�Z b�Ο ��� �� �� �� �� ���  �Κ ���  ��� ͜ 0G͝ B�� ͞ 0:͟ 5 䪩��  ���� 8��� ���  �� ���� 8��� ���  ��ή �ӭ� ͜ 0͝ Ο �� ͞ 0͟  � ��α z�h`H�Z 䪜� ���  �� �� Ӿ �� �� �� �� ��z�h`H�Z 䪩|�� ���  ���� 8���  k��� 8���  Q��� 8���  �� ��z�h`H�Z b���� �� �� �� �� ���  �� ���  ��� ͜ 0`͝ [�� ͞ 0S͟ N�� ͞ � ]�LV�͟ � ��LV� 䪩��  ���� i�� ���  �� ���� i�� ���  ��ή �ӭ� ͜ 0͝ �� ͞ 0͟  � ��� z�h`H�Z 䪜� ���  �� �� �� Ӿ �� ��z�h`H�Z 䪩p�� ���  ���� i��  Q��� i�� �� Z�p��  ��z��  k��� i�� �� Z�p��  ��z��  ���p��  ��z�h`H�Z�� 8�

�� �� 8�



�� z�h`H�Z�� 
���썠 ��썡 �� �� �� �� �� �� �� �퍢 ��퍣 �� �Z�� ��-� � z��Υ �� � �Ȁ�Τ �� � ��� �� �� i�� �� i �� �L)�z�h`H�Z��� ��� �� �� ��  �z�h`H�Z��� ���  ��z�h`H� ��  ����� h`H�Z�� �� �� �� ���� z�h`H�Z�� �� ���� �� ���� z�h`H�Z�� �� �� �� �� ��z�h`H�Z�� �� ���� �� �� ��z�h`H�Z�z � �1��� 8��� �	�� 8��� ة�� ���� ��  |���� ��  |�z�h`H�Z�)�JJJJ��  ���)��  ��z�h`H�Z�� �a��$��b��%��c��&��d��'������ ����� ��� �� ��� ���� �� ��-� ���� Ȳ�-� ���� ��� ���� �� z�h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          H�Z������� ��  Oǭu ����v �	��*��v � ��  �ǭ� �� ���r ����� k���е����Шz�h`H�Z�� ��� �  Oǭu �� ���g��
�����V΀ �  O�� � �u ���  O�� �u �� ���.΀ �  O�� � �u ���  O�� �u �� r�� �z�h`H�Z�v �����M  �� =��� ��� ��u  ��� �v �u  �ǭi��  Oǭu �0��� �� �� ��� �  �ǭ ͊ 0$͋ �� ͌ 0͍ � ���v �u  cŭ͊ 0͋ �͌ 0͍  � ��z�h`H�Z�v �����M  �� =��� ��� ��u  ��� � �v �u  �ǭi�� �� �  Oǭu �0��� �� �� ��� � �� �  �ǭ ͊ 0*͋ %�� ͌ 0͍ �� ����v �u  cŭ͊ 0͋ �͌ 0͍  � ��z�h`H�Z�v �����M  �� =��� ��� ��u  ��� � �v �u  �ǭi�� �� �  Oǭu �0��� �� �� ��� � �� �  �ǭ ͊ 0*͋ %�� ͌ 0͍ �� ����v �u  cŭ͊ 0͋ �͌ 0͍  � ��z�h`H�Z��� �i
�� ��� �i�� z�h`H�Z��� �i
�� ��� �i�� z�h`H�Z��G���A��r  ˹���M  ���u  �� cũ��  �΂ ���8�� �ũ��  �΂ ��z�h`H�Z� �� �� �u ��� � �� ��� ���� ����zh`H�Z�� ��� � ��  ��z�h`H�Z�������u  �� c�z�h`H�Z�������  Yީ���  Yީ���  Yީ���  Yީ ���  Yީ����� �z�h`H�Z�� �0�������� 8���  Y��z�h`H�Z��� m� �� �� i �� �� i �� ة������  Yީ���  Yީ ���  Y�z�h`H�Z��z  �ݩ���� ީ���� Yީ��  Yީ"��  Yީ��<�� � <������ ީ���� Yީ��  Yީ"��  Yީ��<�� � <����x���u  cũ�i ��j �������h  �ܩ��s �  vީ��Z�� ީ��Z��w �  vީ2��  �΂ ��z�h`H�Z��z  �ݩ	��F��  ީ��Z���u  �� � � c� � ��u  �� � � cũ��  �΂ ��z�h`H�Z��z  �ݩ���� ީ���� Yީ��  Yީ"��  Yީ��<�� � <������� ީ��d�� ީ��d���u  cũ�� �   v�������* �ŭ�d���� cũ �� L涩d� cũ�� L����L�z�h`H�Z �ݩ���� ީ��2�� ީ��P�� ީ��n�� ީ����� ީ
��2���u  cŭ  ���� v���L�����, �ŭ� ��� �i� c�L����� �2� c�L����л �ŭ� �0�� �8�� c�L����� �n� c�L��z�h`H�Z���M  �� ˹��u  �� cũ
��<�� ީ2��  �΂ ��z�h`H�Z�� ��� � �u  �ǭ�������t ��t z�h`H�Z���M  ��r ��z  ���w  ��z�h`H�Zz�h`H�Z �ݩ��P���u  cũ�i ��j ���X���h  �ܩ��s �  vީ��(�� ީ��w �  vީ2��  �΂ ��z�h`H�Z������ �z�h`H�Z������
�j ��i  ��z�h`H�Z���<���  Yީ���  Yީ"���  Y�z�h`H�Z�
����� ��� ���� ��~ �~ �  O� c�� �i����
��� ��i�� ���z�h`H�Z�8�

��8�



�z�h`H�Z�8�

��8�



�z�h`H�Z�u �h ��} ��j  �z�h`H�Z�u �h ��} ��j  �z�h`H�Z�u �h ��} ��j  �z�h`H�Z�u �h � �} ��j  �z�h`H�Z�u �h � �} ��j  �z�h`H�Z�u �h � �} ��j  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} �
�i  �z�h`H�Z�u �h � �} �	�i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h �<�} ��i  �z�h`H�Z�u �h �8�} ��i  �z�h`H�Z�u �h �4�} ��i  �z�h`H�Z�u �h �0�} ��i  �z�h`H�Z�u �h �,�} ��i  �z�h`H�Z�u �h �(�} ��i  �z�h`H�Z�u �h �$�} ��i  �z�h`H�Z�u �h � �} ��i  �z�h`H�Z�u �h ��} �	�i  �z�h`H�Z�u �h ��} �
�i  �z�h`H�Z�u �h ��} ��i  �z�h`H�Z�u �h ��} ��i  �z�h`H�Z�u �h ��} ��i  �z�h`H�Z�u �h ��} ��i  �z�h`H�Z�u �h ��} ��i  �z�h`H�Z�� �� ��� ���  �z�h`H�Z�� �� ��� ���  �z�h`H�Z�� �� ��� ���  �z�h`H�Z�� �� � �� ���  �z�h`H�Z�� �� � �� ���  �z�h`H�Z�� �� � �� ���  �z�h`H�Z�� �� � �� ���  �z�h`H�Z�� �� � �� ���  �z�h`H�Z�� �� � �� ���  �z�h`H�Z�� �� �0�� ���  �z�h`H�Z�� �� � �� ���  �z�h`H�Z�� �� ��� ���  �z�h`                                                                                                                                                                                                                                                                                   ���ة��[ ���  ��� � �` � � �a � ��"  �� t ����T ��U �� � �T����U ��� ��X�ߍ&  ��L �H�Z�[ �[ �P0�[ �[ �] � ��] �^ � � ��� ��� �� � ��=��  =�z�(h@H�Z�' )���# �\ �\ ��  ��\ �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                    ���Z �� �� ��z  u� �� Gߩ�J  r� �ݭ   v�����(�# �\ �=�� � � � � � �� �� +���s  ��� �J  r�z  >� �� �� ڳ �� � 7� (� D���� ��� �� �� �� �� �r ��L�í  ���L������� � ��� L���	 v� � �Įz ��L�� ��� �� � � ��� Y�L���� ��L���� 3�L���� � ���� ��� L�¬� ��� ����  ��{ ���{  �͐ � �L�����	 �  �L�����	 A�  �L�����	 c�  �L����� (�  � �Ǭ�� ��� �� �� �� �� �  ��r � �#�r �s �s � � �LZ� b��� � �4 �L;­� � ��� � � �L�í� � � <��t �� q�LZ�L��LR�H�Z��w ��� �r �z �� �� �� ������) �� ))��z�h`H�Z�� �w ʊ


�� m� ���
��>��T �Y��U �T�� ȱT�� �w ��t��T ����U �T�� � �w �����T ����U �T�� z�h`H�Z�z � ���{ �Mz �z z�h`H�Z��j ��i �
�����n ��o ��p ��q �(��j ��i ������n � �o � �p �	�q z�h`H�Z�������������V ���W �V�u  c�ȭi�����i����z�h`H�Z��j ��i �} �u �h  �z�h`H�Z��j ��i  ��z�h`H�Z�w �� �� �� 
m� 


��� � ���� �j�V ���W �8�� ����T ���U �V�TȊm� ���ҩ �����z�h`H�Z�w �� �� �� ��,��T �5��U � �T�ȱT����V �#��W � �V�ȱV�z�h`H�Z�� �� �� �� �� �� �� �� �w �LK����� ��� LK����� ��� ��� ��� LK��!��� ��� ��� ��� ��� ��� LK��?��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� LK��P��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� z�h`H�Z�� ���T ���U � �T�u z�h`H�Z�� ���T ���U � �T�u z�h`H�Z�� ���T ���U � �T�� z�h`H�Z�� ���V ���W � �u �Vz�h`H�Z�� ���V ���W � �u �Vz�h`H�Z�� ��� �u  ��z�h`H�Z�� ���V ���W � �� �Vz�h`H�Z��n |��0u�� ���  Oǭu ����r L��� � �ȀP�����M  �� �� �� �Ȁ9�� ɀ0���  Oǭu �� 2ɀ ɀ�� �Ȁ�� �Ȁ ��z�h`H�Z�� ��� ��u  ��� ��u  �ǩ
�u  �� �� /� � j� D� � O� /� � 4�� D�� ���� ��� �
�u  ��z�h`H�Z � D� � � /� �z�h`H�Z�� ��� ��u  ��� ��u  �ǩ�u  ��� ��u  �� �� /� � j� D� � O� /� � 4�� D�� ���� ��� ��u  ��z�h`H�Z�� � ���  Oǭu ����r LG���p��g�����M  �� �� ���
�u  �� ��� ��u  �ǩ��  ˹ ����
�u  �� c� � �����u  �� c� �΂ �� � ���� Kʀ �z�h`H�Z� ���  Oǭu ��@�� ��u  ��� �
�u  �� ����� ��� �
�u  ��� ��u  �ǀ �z�h`H�Z���  ˹ ����
�u  �� cŭi� �����u  �� cŭ8�� � �����u  �� cŭi� �����u  �� cŭ8�� �΂ �� � Јz�h`H�Z ˹�
�u  �� c�z�h`H�Z ˹��u  �� c�z�h`H�Z��n  �� � j� � O� � 4� ݀ �z�h`H�Z�� �˩�� �˩'�� 8�z�h`H�Z�� ��� �� O� �����i�� L��z�h`H�Z�	������ ��~ �~ �~ �  O� cŭi�� ���	�� ���i����z�h`H�Z��� �i
� �� O� [��i�� ���z�h`H�Z�� �̩�� �̩&�� �z�h`H�Z�� ��� �� O� '�����i�� L��z�h`H�Z�	������ ��~ �~ �~ �  O� cŭi�� ���	�� ���i����z�h`H�Z��� �i
� �� O� u�� �i����z�h`H�Z�� uͩ�� �ͩ%�� �z�h`H�Z�� ��� �� O� A�����i�� L��z�h`H�Z�	������ ��~ �~ �~ �  O� c��i�� ���� �	����i����z�h`H�Z��� �i
� �� O� ��� �i����z�h`H�Z� �z�h`H�Z��o 0|��u�:� ���  Oǭu ����r L��� � �΀P�����M  �� �� �� �΀9�� >π0���  Oǭu �� ]π >π�� �΀�� �΀ ��z�h`H�Z�� ��� ��u  ��� ��u  �ǩ�u  �� �� Z� � �� o� � t� Z� � V�� o�� ���� ��� ��u  ��z�h`H�Z Z� � o� � Z� � o� �z�h`H�Z�� ��� ��u  ��� ��u  �ǩ�u  ��� ��u  �� �� Z� � �� o� � t� Z� � V�� o�� ���� ��� ��u  ��z�h`H�Z�� � ���  Oǭu ����r Lr���p��g�����M  �� �� ����u  �� ��� ��u  �ǩ��  ˹ �����u  �� c� � �����u  �� c� �΂ �� � ���� vЀ >�z�h`H�Z� ���  Oǭu ��@�� ��u  ��� ��u  �� ����� ��� �
�u  ��� ��u  �ǀ �z�h`H�Z���  ˹ �����u  �� cŭ8�� �����u  �� cŭi� � �����u  �� cŭ8�� �����u  �� cŭi� �΂ �� � Јz�h`H�Z ˹��u  �� c�z�h`H�Z ˹��u  �� c�z�h`H�Z��o 0 �� � �� � t� � V� ݀ �z�h`H�Z�� �ѩ�� ҩ%�� `�z�h`H�Z���� � ���  O� A�� ��i����z�h`H�Z�	�����~ ��� �~ �  O� c�� �i����� �	����i����z�h`H�Z����� �i	�  O� ��� �i����z�h`H�Z�� �ҩ�� �ҩ&�� B�z�h`H�Z���� � ���  O� '�� ��i����z�h`H�Z�	�����~ ��� �~ �  O� c�� �i����	�� ���i����z�h`H�Z����� �i	�  O� u�� �i����z�h`H�Z�� �ө�� �ө'�� $�z�h`H�Z���� � ���  O� �� ��i����z�h`H�Z�	�����~ ��� �~ �  O� c�� �i����	�� ���i����z�h`H�Z����� �i	�  O� [�� �i����z�h`H�Z� �z�h`H�Z��p 0e��� ΀ ��  Oǭu ����r L��� � �Ԁ>�����M  �� �� �� �Ԁ'�� IՀ�� IՀ�� �Ԁ�� �Ԁ h�z�h`H�Z�� ��� ��u  ��΀ ��u  �ǩ�u  �� _� 	� � �� � � �� 	� � �� �� ���� ��� ��u  ��z�h`H�Z 	� � � � 	� � � �z�h`H�Z�� ��� ΀  Oǭu ����r L���r��n�����M  �� �� ����u  �� ��� ��u  �ǩ��  ˹ �ŭ8����u  �� c� � �ŭ8����u  �� c� �΂ ���� I�z�h`H�Z ˹��u  �� c�z�h`H�Z ˹��u  �� c�z�h`H�Z��p 0 _� � �� � �� � � ݀ �z�h`H�Z�� �֩�� ��  �֩t�� ��z�h`H�Z�
��� ��� ΀  O� }��i�� ���z�h`H�Z i�z�h`H�Z�
��i�� ��  O� ��� �i����z�h`H�Z�� ש�� ��  Kשx�� U�z�h`H�Z�
��� ��� ΀  O� 弭i�� ���z�h`H�Z i�z�h`H�Z�
��i�� ��  O� _�� �i����z�h`H�Z�� �ש�� ��  �ש|�� ��z�h`H�Z�
��� ��� ΀  O� M��i�� ���z�h`H�Z i�z�h`H�Z�
��i�� ��  O� ǻ� �i����z�h`H�Z� �z�h`H�Z��q l��0e��� � ��  Oǭu ����r L��� � �؀>�����M  �� �� �� �؀'�� ـ�� ـ�� �؀�� �؀ 4�z�h`H�Z�� ��� ��u  ��� ��u  �ǩ�u  �� 0� �� � �� �� � ^� �� � ��� ��� ���� ��� ��u  ��z�h`H�Z �� � �� � �� � �� �z�h`H�Z�� ��� �  Oǭu ����r L����w��s�����M  �� �� ����u  �� ��΀ ��u  �ǩ��  ˹ �ŭi���u  �� c� � �ŭi��	�u  �� c� �΂ �� � ���� �z�h`H�Z ˹��u  �� c�z�h`H�Z ˹�	�u  �� c�z�h`H�Z��q  0� � �� � ^� � �� ݀ �z�h`H�Z�� Vک�� ��  �ک|�� ��z�h`H�Z�
��� ���  O� M�� �i����z�h`H�Z� i��z�h`H�Z�i�� �� �
� O� ǻ� �i����z�h`H�Z�� �ک�� ��  ۩x�� ,�z�h`H�Z�
��� ���  O� �� �i����z�h`H�Z� i��z�h`H�Z�i�� �� �
� O� _�� �i����z�h`H�Z�� �۩�� ��  �۩t�� ��z�h`H�Z�
��� ���  O� }�� �i����z�h`H�Z� i��z�h`H�Z�i�� �� �
� O� ��� �i����z�h`H�Z� �z�h`H�Z�h 
����T ���U �i ��j ���} �| ��V ���W ��Z�| �T-Z �| z�V��� �Ȁ���� ��j ��T i�T �U i �U �L&�z�h`H�Z�h 
����T ���U m� �U �i ��j ����V ���W ���T-Z �V�T i�T �U i �U ��� �Ȁ���� �
�j ��L��z�h`H� �Z  ܩ��Z h`H� �Z  �ܩ��Z h`H�Z�O���� ���� ��z�h`H�Z�/���� ���� ��z�h`H�Z�  �[ �� ��z�h`ڭ  �[ �� ���`H Y����� ��h`H Y�����h`H�[ h`Hڪ���




���)�& �h`H�Z�  ��
���썓 ��썔 � �� �@�� � � ������(���� i0�� �� i �� �� i(�� �� i �� ���Ωߍ& z�h`H�Z�T �@�U � � � �T����U ���z�h`H�Z
����X 轡�Y � �X�$��a��b��c��d�8�7�  v�Ȁ�z�h`H�Z�)�JJJJ�  vފ)�  v�z�h`xH�Z� �a��$��b��%��c��&��d��'�����T ����U �����V ���W ��T-Z �V�T ȲT-Z �V�T ������z�hX`H�Z������ Yީ��� Yީ�� ީ����� �z�hH�Z���M  �� ˹��u  �� cũ2��  �΂ ��z�h`H�Z� �ݩ��� ��j ��i � �� ���� �� ��� ���h  �ܭ� �r� /��� �i ����i �ө�� ����  /ݩ�� �� �� ��� ���i ��h  ���� �� �� ��� ��� �i ��h  �ܭ� �D0 /ݭ� ��� �� ����� �� /ݭ� ���i �� ���h  	ݭ� i�� ���h  �ܭ� ���h  	ݭ� 8��� ���h  �ܭ� �� /݀���^ ���M  ��(��  �΂ ��� ��z�h�� `� � � �  .� 2� � � � � � � � �* �G �O � ���H �S `� ���%�+ � .�$ � �% �  d��+ �+ �& � � ���%�8 � 2�1 � �2 �  ���8 �8 �3 � t� ���X� ���� � .� � �	 �  �� ���� � 2� � � �  ��� � �
 � ��� � � � ��S ��� B� ��`� �� ȱ�	 ȱ�
 ȱ� ȱ� )
���� 轰� � )0� ȭO �	�����H Ȍ � � �
 � �Ls�  ^�� �� � �� ��Ȍ � ���! �"�$ ȱ"�% ȱ"�& ȱ"�' ȱ"�( )
����) 轰�* �( )0�- ȱ"����H Ȍ! �+ �, �& � �� � � �M )����� �.  t�`�. �/�1 ȱ/�2 ȱ/�3 ȱ/�4 ȱ/�5 )
����6 轰�7 �5 )0�: ȱ/����H Ȍ. �8 �9 �3 � Ы� � � �M )��@К��� �!  ‍� �� ȱ� ȱ� ȱ� ȱ� )
���� 轰� � )0�  ȭO �	�����H Ȍ � � � � Х�  |�� �� � �� ��Ȍ � ���J 
��Z�K �Z�L �K� ȱK� `�J 
��d�K �d�L �K� ȱK� `H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; � �8�� �� )0� Ȍ ����� � � �; � z�h`H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; �  �8��  �� )0�  Ȍ ����� � � �; � z�h`H�Z�' )?	@�; �' I��-; �; �, �)��( )@��J��; �; �- �8��- ��( )0�- Ȍ, �)����, �( �, �; � z�h`H�Z�4 )?	@�; �4 I��-; �; �9 �6��5 )@��J��; �; �: �8��: ��5 )0�: Ȍ9 �6����9 �5 �9 �; � z�h`� `� `�H ���S  B�`H�Z�H ���%�I ���H �O �I )?
����Q ���R �P  �z�h`�O �* �G `�P �Q�C ȱQ�= ȱQ�> ȱQ�D )
����@ 轰�A �D )0�E ȌP �? �B �C � u�S `H�Z�O ���Ln�= �F �C I�F )��F �B �@��D )@��J��F �F �E �8��E ��D )0�E ȌB �@����B �D �B �C )�; �I )����
�@����; �; �F �( �; �G ��* �G �? �? �> � �z�h`H�Z�  ^�  |� � �� �  �� �� �� �� B��� z�h`H�Z� � �
� � ��N �M )?�N �Q�� �K�N 
����" ���/ 轔�# ���0 �! �. � � � �M )�����  t�M ���  � B�z�h` K�� _�� K�� _�� q�� _�� K�� _�� K�� _�� q�� _�� 8�� K�� _�� q�� q�� _�� K�� _�� q(��     � �
�!� �
�!� �
�!  q
�!� �
�!� �
�!� �(�!  �
�!� �
�!� �
�!  q
�!� �
�!� �
�!� �(�!  �
�!� �
�!� �
�!  q
�!� �
�!� �
�!� �(�!      � �
�!� �
�!� �
�!  q
�!� �
�!� �
�!� �(�! .
�!� �
�!� �
�!  �
�!� �
�!� �
�!� �(�!  �
�!� �
�!� �
�! .
�!� �
�!� �
�!� ��!� ��!        ?� � G� � K� � ?� � G� � K� � T� � K� � T� � _� �     � ?�!� 8�� ?�!� G�� ?�!� G�� K�!� G�� K�!� T�� K�!� T�� _�!�     � �(�� �(�� �(�� �(�� �(�� �(��     � ��� /2��     � KP���     � <��     � _ȧ �     � ȧ �     � ���� _���     � �� d�� T�� ?��     ������-�@�K�W�   � � � � � � � � � �      �J   �J      �   �     ( �
     ( �
    	

			�
	�	��













�





















�

		�
	�






	
	
		



	
	
				
	
			�n�x����r�|�����  �� �  @�  @�  ��  ��  ��  ��      j�|�������j��������V�a�n�u��������aGAMEaaOVERa$PAUSE$LEVEL$STAGE$END$TIME$CONTINUE$PRESSaaSLaKEY$PRESSaaSTaKEY$PRESSaaUPaKEY$PRESSaaDNaKEY$PRESSaSTARTaKEY$LIFE$OUTaOFaTIME$YOURaSCOREa$YOURaaSCOREaaIS$COPYRIGHT$BON$HIGHaSCOREa$LEVELaaSELECT$EASY$NORMAL$HARD$�������������������+�;�@�L�X�h�r�v����� �@����� �@����� �@����� �@�����З  � �P��� � � 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____^^^^^^____  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����������������������������������������������������������������������������������������������������������������������������������������������������  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`����  @`���� 
��������� "���������$&(*,.02468:<>@BDFHJLNPRTVX���������������������������Z[\]^_`abcdefghijklmnopqrst���������������������������uvwxyz{|}���������  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              Z� ���