L�H�Z�� �l������l���)�k��l����� � �l������l�e��j%����
���������� � ��j��� �����j���e��i �� �k�����ڢ������������e��i �� � ���Ȁ�� �k�����ڢ����������� ����Ȁ� =� !�������z�h`H�Z�:
��/���0��� ���H�
�hH)�JJJJ��h)���-���-e��i �z�h`N�\�#H�Z� ��������j���	���� p���� М} r�����z�h`H�Z�L��L��K� �mL��y����z����{�������:� Т ��m���������%i�i�� %�����4����%i�i�� %�λ������%�i�� %�κ�m���ͽ���L� ��Lz�h` H�Z�
��L���M��� ���ȱ���k
��僅�情� ����y���m���H)�JJJJ��h)��z�h`                                                                            H����������  ЭM��'��#��H���  �h���M����������
��������~h`H�j%�)���%���%��  ЭM��mI�M �h`ń-�������
�;�ڈA��������������Ӎ;��{���������T�[�-�7����%��������8�ш:���������������ύ3��s�����{�y�N�N��#������I����v�|���7�4�������������ߌ��΍-��m�����k�d�:�5������H�                       DDDAD   D@   @   @   @   @   D   DDDDADDDDD@  4@�  @�  @   D@   @  @  �DDDDDGc!1U!1UDDDD@  D@   @   @   @    @   D@  DDDDDDDDDN� �N���@ �@ �  �� �N���N� �DDDDD�3s5u3s5eDDDDD@   @    DD DDDAD@DDD@   @   @       @   @   @   DDDDDAD@DDD@  �@  D@  D@   @   @ D@D@ADDDDDD@   @ @@ @@ @@ @@ @@   4DD@DDDD@DD@   @���@� @� @�@� @ �DDDDD�08h`XPDDf"Df3v3f�D@DDD@   @   @ @@ @@ @@   @   DDDDDDA@AD@A  A�DD � @�@  @DDD@A@AD@DAD@  D  �� D@��D@  AD@DA@ADDDDD 4@ @@ @  @  DDDDDADDDD      DD� ADDA0X8P��v'fw3Uw3U"De#UDDDD  @   @   D@  @  @  @  DDDDDADODD@D@@  @   @   D   D@ ADD@H"Dfq3UrDDDAD   D@ D 4@ D @   @ D O D D   DDDDA"DUDDD@DM   M����C�� � ����@�� �@����@   DDDDDDD DDD      DDD DDDD DD� ��    DDD@A@A@A�px�"Df�CUDdaDDDA@  A@  A@  AD@ DD@  @  @  $DDDDDDDAD   D@� @   B  C   @ �D   DDDDA�3U"DfrUQPQPQUPUU      UU  Q  QUUQUUQPQUUP Q    QUUP QPQUUQ�D&URUUUP UP UP � P �P � UP UP UUUUUUQP  QP��QP  QUU UU  � UUUtW1c6EuUUQQ   QUUUQUUQ# Q�Q  QU QQUQ QU UQ  Q   QP UQP QUUQ@H!C%1#SAEUQ�QU UQQ   QUUQ QUQUUUUQP   QP   QU%U�QUU$%C3cUQU UP U U QU UP UPUPQUUUQPU U     PU UUUUQUQUUQ   QUUQUQ X�CECUUQUUS URP�  �PUPUUQUUUUQP QP Q_ QUUQ rD#sUUUUU   P _PU UP   %PU UP PP   UUUUUQPUUUUP   PPUP %P   P PPUP   UUUUUU  UU UUUUUQU�  U]���] ��]�  ] ���]� �U�� UUPUQPQPQPQUU Q   QUUUQ H�P@X��cACEC"R!QSPUUUUP   PU UPU UP   PU UPU UP   �UUUUUUPUUU] ��P ���] ��]� ��]� �]�� �]�� UUUPUUUU 5PP�UUP�  P���P���P   UUUUPQx0xACE3Uq6fUUUQU   UP �P�0�P   P� �P �U   UUUUQ1affff`f`&`   `� �`� �`   ` � `f`ffffffff```f``   `   `   `f`b`6ffff�SEtDqffff`   `  f`  ` ``  ``` `   ffffffff`   `�� `   ` ��`   `  ��`   �fff`ffffff`� 6 �  `�� ` � ` ��`  �`  �ffffffffff`   &n� ��`   ` � `   n� ��`   ffff( @Hx�q1dBBBfffff`   &`�  f   f � a   af  �fo   ffffffffff`   `   ff ff a aff ffb   6fffff�%Q#CQEffff`f`�`   f��f��a��af   f`f`6ffff"%RUfff` &`�`�ff`�`  �` ��f`  ffffffab a`�a`�fff`�  `�   `���`   fffffa a aff ff`   ` � `���`   &ffffffff  &ff  `  � ��`  �ff    �fffffffc  `�`�f`� `�� `   `  fffffa�@����QS5#6A4T3Ss!A4fffff`   `��`  ff ff a a a`af`f` fn �f`   ` � `   fn �f` `ff`a`a`a`f `f`a`a`afa` a`affa  XP8PX@1QC1QCQQQUQQ QUQQQUUUUUR   P �P �  P � P �P� ^  �UUUUUQQQQUUUUU  P   P����UUUUUQQQQUUUUUP    P��P  P�P P��R   UUUUUUUUQU  UP   P � P��P � P   U   UUUUQ ���T'!AaS!Aa!A3UUUU     UUUUUU�UU  %    UUUQ0QUUUUP �P�   P �UU  UUUQUUP%UUUP    UUUPPUU@H��c�E#CSs�wpwy�   ������ � �  �� �����   ��wpw|wwwww     wwwww�wwy�  (w���  ��w����  �ww|�|wy�   �����   8�www|�wwwy�   (���������   �w��|������ PX�X@���Q3r5Uu1Q�wwwy�   �  ��  ��  ��  ��  ��   �wpw|�wwwy�   (��w���w��   �   �   �   �ww|�pwwy�   ��  �� ��� ��  ��   �   8�www|�wpwy�   �� ��� ��   �� ��� ��   (�www|XP(0��A4TsAaCECEafffa/  a   a   a   a   afffaaf a`    a`      a` aff0a`    a`  aff ff`    ffffffffff     ff ff a`    a`      affffa` f   a    f   a`  af��"AWQ#Cc%2R$D2RDFA4T&2R$DU QP P Q QP    QUUUQUQ#QP    QP   P      QP UQUQR  QUU UUP    UUUUU Q   Q �  Q  QU�@A1At2RD62R4AACE`ffff`   �m����m����m�  m���` ��`   fffffba`` a` `  a`  `  afffffffff   `    `  `&ff&` ` `  0  ff`fffffff`  a`  `  a` ` a`bafX�`��1Qq41QqSrtvT1QUUUUUP   QP  P  QP P  QP  P  QUUUUUUUUUU�   P    P   P     UUUUUUUUUUP       P   P U PPPQ%UUQQUUPQ%PPP U P   P   P   UPUUUUUUU   QP  Q QQP  QUUUUU�8@w'��1Q1QqS1Qq6s1QEfwww��  �� ��| ��   �y �� ��   �www�ACEj�n�s�v�y�����������������ʙؙ             0

0

4

 4

                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           L/�L�L��L�L��                              D�H� �	������������ ǩo��� ��d���� � �� ��D�������	 � � ���i��8�� � ����T�ة���  �< �:��h`�H�H�H�H������������ �h�h�h�h�`H�Z�/���� ���� ��z�h`H�Z 7� �� A� ]��I�J�ろ�炍 y� � �ĩ������$ ũD�����' ŭ  ���
���K���s�敏��  �J����J ]��ろ�炍 y����� �I A��ろ�炍 y���������  �J����J ]��ろ�炍 y����������  � � �� � �ĩD�����$ ũ������' ŭ  ������"���������������J ]������ ������  � �� ��z�h`H� �	�<�����I q� ��h`H� �	�������J q� ��h`H �ĩ�	������ �h`H�Z� �	� �
��ろ�炍������ ����ߠ �
��낍�킍�������� ������z�h`ZZPPT��STAGE$LEVEL$H�Z 7ĩ �	� �� ��$���%������� �  �ȩ$��p������� �ũ�����( ũ(�� ����� �ũ@���������� �Š �A��1�� �	��  ��( ����� �� �.���/���ȭ0���1�� ǀ� �ĩ���  �z�h`BON TREASURE$1992$PRESS  START$H�Z 7ĩs��<������� �ũ��� �����	�� �Ţ � � �	�	����(���)������ �ȩ1������  �� ��󽁄�
��*���+�� ǀ� �ĩ���  �z�h` GOOD$GO ON PLEASE$H�Z 7ĩ �	� �� ��&���'������� �  �ȩ@��s��
����� �ũ���������� �Šȭ  �� ��� �ĩR��  � -��R��  �z�h`WIN$CONGRATULATE YOU$H�Z 7Ģ ��������ڊ
������� ������ݠȭ  �� ��� ��z�h`DESIGNER$MISS XIAOYING GAO$MUSIC$MR XUHUI HU$PICTURE$MR YOUG BAN$(@Xp�Hک�H�I
mJ�K�L��������K�腍��h`
 #N�@����  ȃՃڃ���������*���A�n�w���������2������(f������� � � � );Mcz�����+?Sex�����'?[{����#B\y����&Ig����1St���,Rv����;Yt�����	)	D	]	w	�	�	�	�	�	�	

5
G
Z
k
|
�
�
 ����� �������� � ������� �  ���? �� �  ������? �� � ��� ���� �� � ��� ���� �� � ��? ������ � ��  �
���� < < �� ��
����� < < �� ��	��? ��� ��?� �  ���	�� �� ��?�� �  ���	�� ���� �?��<  � ��
�	��  �����?�� �?�?�
���?  ���?��? ��� 
��� ���?��� �?�� �	��� �	��? ���� �  �	��� ����� �?  �	��� ������  �	����?������ 	���� ?����� 	��� � �����?�  	���? � � ���� �	���? ��?��� ���? �	���  ?����?<  ���?�? �	��� �  ��� ���� ? �����? ����? ����  � ������ �?���? �� �? ���� ���� ��? �  ��� ������ �� �� � ���?  ������ ��  ���? �����?  0����� �� ���� ����� �����??
 � ����� ���� � ��  �� � �������� �" ���? � ��
����� �  ������ ���� ����� � 
 �����? ���? �����* � �������?���? ��� ����?������ � ��� (
 �����<�� ���� ����  ����?�� ���� ����?  ����?��  ���� ����?  ����? ��� ����  �����  ���� ���� (	 � ���� �  ���� ���� � �
���� � ���� ����  �* �� �" ���<� ���� ����� ��0 � ���?�� ���� ���   �  �0� ������ ��� ���:      �0 �   ���� ����? �? ��> ��  �0 �����0 ���? ����> ��  �� � ����?������� ����? �|U�    *  ���?�� ��� �����? �WUU� �  ���?��  ��� �?��� ��U�u �����  ���� �?���� ��U�] ����  ���� �?���� �pU�]5 �U���� ���� ��뮪 �pU�}5 �@T����� ����  ����> �pU]Wu5 �U���+�� ����  �����> �\U]W��  @UU���8�? ����  �����; ��_�W�W� @U�����/ ����  �����? �0\�W�_WSTU��_���� ����  ���? �0\\_WU����?� ����?  ���? �0\??\_]U��&��?���� ��� �0\??\_]UUP��~���������� �P5_?\?\W]UTUZ��������j� �T�w_�UWUAUU_���?�����j� �TUw�W���UTUկ�W�� �	����  PU�wU��= PUU՗�����������  TUU��U�W� U���������� @UU���UU5 PU����
�
��� ���WUU�?  TU���
��� ���]UU�� �P���
���> �pu�U�wW ����_��� �\uW�uW ���������� �\UU\UU �����W�������� �\UU\UU ��<bU}�
��Z� �\UU\UU  �����z�
���� �������  ��[�j��
����: ���;���  �/�z
�
���Z� �軮���
  �K���	����� ����
  �P�U�	�
�����  ���
  �z�
�����  ��� ���{�
�
����n ��
  �����
����j � ���o������? ��� ������
����j� ���� ���������� ��
  ��
������ � �*  ���������� ���� ����    (�� ������? ��� ����� ����    ����? �  � ��    ������   �� ����
���; � ��
"""�(e� � � � � � �   8Pi�����)CZ{����8Wt����!:Sl������&@Ys�����9Xp�����1Om�����2Mj�����		2	G	[	n	�	�	�	�	�	�	�	�	�	�	� $ � �      � �     � � �  ��� � � �  � � �  �� �� �	 � �  ��    � � � �   ��   �7 � � �   ��  �7 �� � �   ��  �  ���U� � � � �   �
 ��pU5p � � � � �  � �\_U�p � �          �p_U�\ � �       � �pMU�� � � ,  �  ��T�� � � , � �< �5 � � � �� � � �  �� � �W3 � � � 	 �( � �W= � � �  �� �� �( �  �W� 0 � � , �<�? (	 �* �( �\5��? � �  ��T10 �* �� ��? �� � �  �U�C5 �* �� ��U � �  W�W5P5
 �*  � �� �� � � W�T �� �(( �ʯ ��� � �  \U @U
 �* �*�>  �? � �  \U�  ���� ��/��	 � �  pU� 
 � �����? � �  �U�� **��  �
 ���� � �   _UU*( ��  �:  ��� � �  ��� ���
  �
  � ��? � � �� ���*�*�
 ( �  �? � �  ��� ��
( ���� < � �  �� ��� ����� � �  �( ��
   ����� � �  ���  
  ����> � �  ���  � ���� � �  �� �
  ����� � �  �� �� ��	 ��
 � �  ��  ��  �?
 ��	 � �  �� �� ��:	 � �  �� �� ���	 � �  �� �< ���	 � �  � � � ���	 � �  � � �� ���	 � �  � , �� ���� � �  � , �< ���� � �  �>��� �� ���� � �  �:ךּ  ? ���*2 � �  �:묪�� ����2 � �  +��+��? ��*��2 � �  +�+��� ��*��: � � ���*�> ��*�� � � ������� ����� � � �*��*� �� ���: � � ��������?	 ��> ���8 � �   �� ���� ��� ���: � �  ��? ��
����(� � �  ���  0�꿊�(�� � �  ��� ,�
���*��� � �  �� ����**����� � �  ��> �����*���    �  �0� ��**��*��:�  ;  �  �0� ��*��*����  ;  �  ��� �< ����������:  �  ��� �� ����������:  �  ��� �� ���������:�:  �  �+�  � �𿨢��*:��  �  �/� �� ������(��� �  ��� �� �����꿪� �  ����� �����*� �  ������  � �𫪨�(� �  ����>��  � ������� �  ����:��  �
 ����  �� �  �����(? �	 �� � �   <+��Ⱚ�: +>� ��� � �   ���*Ⱚ� +��< ��? � �  �����갪�>���� �� � �  ������ê�:�"��� �� � �  �������*���"�(�� � �  ���������(��? � �   ���������"(�? � �   �(�������� � � ��*��������> � � �>�������� � � �ꬪ�*�*���? � � ���*�*�(��? � � ���*����� � � ���
����� � � ������� � � ̋������ � � �������? � � ����? � � ,��� � � ���� � � ����! � � �# � &�� $]� � � � � � � +<Obu������&@[w����#?_~���� A_{����1Rs����/Pq����5Qn����-Jg����	%	C	[	t	�	�	�	�	�	�	� � #���" �� �� �� ��\5 �� �|54 �� �\44 �� ��4 �� �\Q5 �� ���L �� �� �� �? ���_ �� ���� �\s= �� �|�� �� �� �\u� �u � �� �T7 �\}P� �� �\1� ��s�� �� ���S5 �p4? �� ��<5 �p5 �� �� ��5W �� �\� �� �p� �	 �\�� �� ��W1 � �<QQ �� ���� ���� ��P �� ��� �_�u= ����U� �� �? ��U�]� �pU�A� �� �� �\U� �p@}QW �� �\ �WU�5 �p ]�@ �� �� ��U�� �p�P �� �W� �pU� ��?@u �� �G}5 �\U� �_�t �� � ]4 �WU� �p3T5 �� �W�4 �WU�5 �_0� �� �|�@5 ��U�� ��5 �� ���_ ��UU�UU�� ��A]� �� ���� �pU� _U5�� ��Es� �� �p1S �pU5�U�� ��Ws� �� �\@E5 �\U�U�_ ���? �� �P4 �\U�U�_ ��� �� ��5 �\U�� �_ �_�U �� ��\= �WU�� �_ ��A �� �\5� �WU�� �_ �uQ �� �� �WU�� �_ �WT� ��	 ��WU � �_ �|��? ��	 �p5WU�� �_? ���P� ��	 �p�WU�� �_�� �|�� ��	 �p_WU�� �_}� �W� � ��	 �pwWU�u�W]� ��PC= �� � �pW_U5�}5�W�� ��tA �� W �pW_U� _s��U]� ���E ��?G �pWsUU�WsU�]� ��U ����E� �pW�U��pU�]� ��W ���QA_ �p]WUU5pU�]� �� ���@ ��]\UUpU��5  �? ���0 ���pU�pU�W �� ��_3P �W��? pU�W ���: ��p�� �� \ 33 pU�� ���� ���=4 ����3 ? pU�? ���� ��\�� ��� 0 �pUU�  ���� ��PQ  �: 0 �pUU� ����� ���  ���� � �\UU� �����> ��4G  ����� �WUU5 �:����3 ��5W �����>  �WUU5 �ꫪ�>0 ��W� ������  �U���ꯪ�� ��� �ê�:� <sU���ꬪ�?� �� ������� �_U���ꫪ�  �� �0�Ϊ���U������ �� �������_U����>� � �� �� ����_UUի���  W �� �? �������?�����  ?G �� ��? ��� ����� ��E� ��	 �����: �  �  �QA_ �� ���? ����? ��@ �� �  ��0 �� ��?� �� �_3P �� ���\5 �� �� �p�� �� �p�4 �\5 �W ��=4 �� �pP5  �4  ?G �\�� �� �pEE  \54 ��E� �PQ �� ��L� ��4��QA_ �� �� ��U P��W�@ �4G �� ���  @�S�0 �5W �� �p�P \U� _3P �W� �� �\ 5� ��Pp�� �� �� �@4 �\�L��=4 �� �P_� ��@? \�� �� �\�p�  �T@ PQ �� ��?p�  �tA � �� ��?  ��5 4G �� ���4 5W �� ��E5 W� �� �W\ � �� �� � �1                 ���          _�u=         �U�]�        \UUUU        WUUUU5       �UUUUU�       pUUUUUU      \UUUUUU      WUUUUUU      WUUUUUU5     �UUUUUUU�     �UU�UU��     pU� _U5��     pU5�U��     \U�U�_    \U�U�_    \U�� �_    WU�� �_    WU�� �_    WU�� �_  �WU � �_  p5WU�� �_? p�WU�� �_�� p_WU�� �_}� pwWU�u�W]� pW_U5�}5�W�� pW_U� _s��U]� pWsUU�WsUUU]� pW�UUU�pUUU]� p]WUU5pUUU]� �]\UUpUUU�5 ��pU�pUUUW  W��? pUUUW  \ 33 pUUU� ��3 ? pUUU? � 0    pUU�  �: 0    pUU� ��� �    \UU� ����    WUU5 �:�>    WUU5 ����  �UUU���:� <sUUU������� �_UUU��ꫪΪ���UUU���������_UUUU����������_UUի���� �������?����? ���    ����1      �0           ���          |]��         �Wu�U        pUUUU5        \UUUU�        WUUUUU      �UUUUUU      pUUUUUU5      pUUUUUU�      \UUUUUU�      WUUUUUUU     W�WUU�UU     W\U� _U     �pU�\U    ��pU�pU5    ��?�U�pU5    ��?� ��U5    ��?� ��U�    p�?� ��U�    p�� ��U�    p�� � �U�� �p�� ��U�\ Ws�?� ��U�W W}�?0 �pU�� �u�p]�pU�� ww�\}�\U�� wuU�W�� WU�� wuUUU���UU�� �uUUUWUUU�� �uUUU\UU�pu \UUUpUU5pu p�UUU�WU�_ ��UUU ��p�  �UUU �� p5 : �UUU �� ���  WUU     �� WUU     �� WUU5     ��: \UU�    ���� \UU�   � �����_UUU�  ����:��zUUU�< 0��ꫪ�UUU�3 ﯯ�����_UUU����������zUUUU����������WUU����������:������� ���?    ��: � ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              )��������������������        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        ���������������������
(                                    ?        ��        #�       �"2      ���8      ���2      ��_;     �|Ug    �3sUg    0��U�    ���U�6   0~�U6   &���U5   &�]�W}  �&�uWW]5  ���uW^�5 �� WUz�5  � WU~�5 HZ�e�����Zre��Zv5V��p���Y]5T��\}��Z]5�  Wϥåu�  �U��ZU�  p� �åU�  p����Z]U pժ��UuU� �����UU�*  �
� W��       ��                                                                       
(                                                             " �      ���      hb�     Xb	�     ��%�     ��%�    �����   �����   XYUi�   hVUe�   Xv�g� � ��U_�Y
 � j�U_��&�������
 �ꎪ*      <;       ��      ���0     �����   ����,""  ���8���+��"">��
 ����("�� �
""���m�"��� �~��� ""  ��ꮺ>�  ������ �ϫ��>�� �����     ����� �  0����  �]�o�    ������    ��ݪ��    �����
'                                 �       �3�     �3���?    <�<33�   ��0����  0��17�<  �puq_�  <_u�w=�  �\��w�� <WWWU=? ��U5?W��� �uU=?�W]3�uU??U��<s]U�?�U]?3]����W]�<p]�?��_}�3�u����uU?�u�����U3�u����uW?pw����uW3pw�����uW?p]U����]W�]U����]]�uU����W]�uU����W]\�U����Wu\WW����Wu\]]����W�5\]u����V��\u� ��U�W]�   �UW�?0�   ��_= 33  3 � ��  33    0�   0           
(                                                      ���      ����    ������    ������  �������  �������?  ��������  �������� �������������������������������������������U���������������WU�����������������������?"""�������������   �����   �������������    �� ��    �? �������� �    ��      ��       �?   ������                                                              (e� �  � � � � � �� � � � � � &8L`t�������"5H[o������6Oi������������*BZu������)[>Qdw��������*>PZdnx��� � � � �'��* ���  ����
  ��  �  �
  �  �� �
  �� �(  �( �   � ��  �
 ��  ���  �� �*  ����*  �����  �� � ��*  *  �( �
 ���  �  �
 �( ��� ��  �� �� ��* �
  �� �� ��
 �  �  ��
 �� �(  �( �
 �� �   � �* �� ��  � �* �� ��  � �� �� ��  � ��  �� ��  � �
*  �� ��  � �
� *� ��  � �
���� ��  �( �   � �   �( ��   � �(  �� ��    
 �(  �� �� �  
 �
  �� �( �  ( ��  �
 �* �  � ��  ��  �� �  �
  (  ���
 �     � ��� 
 ����
    � ���

 
 ��  � �      ��  �
 
 �
  �  ���
 �
  �	 	 �� �
  � �
  � �
	 	 �� �(  � �  � �(	 	 �( �   � �  ( � 	 	 � ��  � �   ��	 	 �
 ��  � �  
 ��	 	 � �� � �   �� 	 � ��� ���� �� 	 �
 ��  � �  
 ��	 	 �( ��  � �  ( ��	 	 �( �(  � �
  ( �(	 	 �� �
  ���
  � �
	 	 ��  �  �   ,  �  �	 
 �*  � �8   � �*  �
 
 �� ��    � �� *
 
 ����*�    ���
  �� �� �  ,*  *  �� �* �  �  �  �
 �( �    ��  �� �� �  ( �
  �� �� �  
 �  �  ��     �(  � �
 �� � ��  � �
���
� ��  � �
�  �� ��  � �

  �� ��  � �� �� ��  � �� �� ��  �( ��
 �� �(  �� �� ��
 �(  �� �� ��
 �
  �� �( ��* ��  �
 �
 ��� ��  ��  �   ��
  (  ��
 �  ��� �
  ���
  �����  �
 ��  �( ��  �( �(  �� �
  ��  �  �*  �  �� *  ���� !  0       �0     0�0     �0      �0      �?     �U�   0_UU   �UUU5   WWUU%  �UWUU�  ��WUU�  ��U]W�  puU]WU p]�W�W? \]�W�W� ]__� W_��_� W_��_� W]�_�_�]uW�}uu�U��]�wUUU�] �U�_uu �UUuu5 ��WUU�? pwWUUw7 \�}U��� W���_�UWUUWUUWUUWUUWUUWUU������!    0     �0     00     �0     0     ��     _U=    �UU�3   pUUU�   `UUUW  \UUUW  \UUU_  \U�U]  WU�Uu5 �W�U��5 W�U��� �������W���W����U�]�W�w��]�U�uu�]UUUu uu��U�  puuUU  ��UUU� pwWUUw7 \�}U��� W���_�UWUUWUUWUUWUUWUUWUU������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          πӀ؀ۀހ��������#�/�=�7�y�����?���K���ρ�S���ׂ�[���߃!�c����)�k����1�s�����9�{�����A���ň�I���͉�Q���Պ���������#���'�)�+�-�/�1�3�5�Ø���\���L�G���?���Þ���˟�O�����ͣ������Ӣ��¦��Ld�             0

0

4

 4

 UUUU                                           @@@@    @@@@    @@@@    @@@@  ����  �3���ì:�3�����3ϳ3�γγγγγ3����3�3���ì:�3���  ���������ê��ÿ��ð������0���0���0��0��0��0��0��0��0��0��������?�����|�~U��~U�5|U��|U��U��?V��w��w��w_���U�_��?_����� �  0  0  � � 0(0��0;�:�������:�:��� ��  �:  �  �   � �� 0�: ��� <<��?��1���à��� �3 ��<���0��:��� � 0000����    �������Ã��Ã��Ã�������WW]�������U�����    0000������0��03��3��� �� �0��03���3�� �� ��0�03���3��� �  �� 0000���0   �����0� 0�00�0��������]� ���0W��0��� ���� 3�� 000���3   3��� �������3���3��� �]�����W3��3�  ��0 ����0��3�� 3��� 33��� W]u����UW3���3    00 3���03�0 �������<,� ,,�0,,�0,,������uu� ���0WW�0����   �000 ��� ����ԃ���kii飠��[ZZڃ���kii駠��[ZZڃ���kii駠��[ZZڃ�����������(�(�*�*�������������������""���*��*���*�*���"��������������(     ����  ��  �0  �  �����WU��W������;Wu�:W��WU�WU�WU���� �?  0�� ?  �;  �;  �� �;3 �� �;  �;  �;  �;  ��? ����������������\UU\�W;���� ����E��RZ찦b�()�����Wu�:WU�:WU�WU�WU����      ����  �0  �  �����WU��������������W}�:���:wU����WU���� ����            � �� � �
(                  �  �  �  � ���?O���?��7��7��7>���883���p�����     @  �  �  � @@��G�����G@@ �  
  �  
  ��  �'  @	  � l5��=��    �"�(>0B�0B�0B�0 B��B�Z� �� L:�? �  ��� ��� �         �  4 �C��_��W��\P5\UU5pUU�UU �� ?  ��?�7p�W�UU0_�0��0  00�?��: �� �� �33�0��3�  ��    �?��|�W=�UU0_��0��  �  00  �� ���00������  �  ����_�?�������\5�<W�<��_�?�03�0����?�3����?�  �   �    ����_�?��?��?�\5?<W�<��W���0��0����?���?� ��  ��    �?  _�  W� ������������?w�W���W����\�5��W�_� �����?  �� �?  _�  W� ������������?wUU��UU�����\�5��W _����?����  ���0  �003��3� �� �UU�W����3�\�5p��p��W�?<�?�0���?      ����003��3� �� �UU?\�5��7\�35p���UU�W��?<�?�  �� �  �  �?  p <p<�_��UU�5\ 7� ��T��WpUU��?��00  �? �  �  �?  p  p �_���UU�p � �W��WpUU����00�?�   �  0 ��p5\����p3��3��3�0<�<��p5\>���:�^������   �  0 ��p5\p�S��?|�W=\�W5\�W5���?���5\����^�:����  �� �? ���  0  0<<0?�0?�0��   �� ��� �����:�����?��  �� �? ���  0  0<<0?�0?�0��   ��  �� �����:����:���?��� ���? ��������:����몪������� 3���� ������ ��� �0?���<�  ��<� 0�? �<����?<���  ��<��  �><��������>  ���������  ���?  ������������몪��������? ����� ��ê��� ��� �0?�� �  �� � 0�? � �����? ������� ���?�> ����������>  ���������          ���    ����   𪪪�  �����:  �ê��� �� �� ��:<<0��00���������������:�������?�������:�������:�������0333333  ���    ����   𪪪�  �����:  ������ ��0��:�;0��� ;� �����ê:�������:�������:��?  ���;      쫪��������������3333333�  �� �  0  ���3<<�����<<�  �  �����0��0�30�30�30��?�ϳ<<�������<<��<<���?����?0��0��������:�������� ���  ��  �� �  0  ���3<<�����<<�  �  �����0��0�30��?��33��30�30�������<<�3<<�3�?�����?0  00�?�0�?�� ��������? �                �  0 �?���3����+�3��0���3�?�3�?�3�?�����  �3���2�׿0ޯ���O����_����?p��p��pUU�UU�UU0W���?33��3��  �  0  �  0  �? �����3���+�3��0��?3�?�3�?�3�?�����  �3���2�׿0ޯ���O����_����?p��p��p��p����{0w��\533���3�� ��    �   � 0�?  0�ó�0  �γ����êγ�?  ����:    ��    �00    ��      �      0  �  0  <�  �  �< ?���<�WU�� �UU � pUU5 � p}�5 � p}�5 �pUU5 ��UU���3<WU�03����<�0<� �00�?���?� ��� �    �>�:    ���    �����������    ��          �  �� �   0 0�?  ������0�?  �;0;    �0    �00    ��      �      0  ��  0  WU ��UU�< UU�<�|}��� p}�5 � pUU5 �0�UU=0�0�WU;0����:<�0�:?3�0<�:�000 �� 0����00 ?��� �  �� � �� �>�:    ���    �����������    ��               �?      ��    �7p=    |p�  �W�U=  |U�U���_U W<<p�  W���  �3��?  _3��� �U�pUpU�?�_UpUU�UUpU��sWUpUuW�]U�UuW�]U _UW�U�  pU�_U  pU��U  |ժ�W= �׵��^��յ�^Wpյ��^W|5����\=\����p5\�����5�ܪ�70?0p���33�UU���?�����  0      �      p  �  p  p  p5  \  p�  W  pU�U  p���_  p<<p  p��  ��3�  _�3�� �U�pU\U�?�_U5WUU�UU�WU��sWU�\UuW�]U5�UuW�]U _UW�U�  p�UUW  p�u]W  |�u]W= ���u]W���5�\Wp���[_W|5����\=\����p5\�����5�̪�30?00���33�  ���?�����   � �   �p�  � � � �: �5 ���������U�UU��^U�UU���������WU�uU� ��]�� ���uW�_������_�����_:�����W:��4��:�V4p�:�Z34̥���W��|?�0�7\�  �5\=���p5W=���:|�W����?w�W]���u�W�  ��W�U��U�����UU��װ������ê���۫�(�(��3�0���������?   �   �  p  �;  �  �;  �5  �� ���� ��U�UU�:�^U�UU�:��������WU�uU� ��]�� ���uW�_������_���4�_:���4�W:��4��:�V4p�:�Z34̥���W��|?�0�7\�  �5\=���p5W�  ��W]���_u�W]UTUu�WU�WU��W�UUUU�����UU��װ������ê���۫�(�(��3�0���������? ��    �pU  �UpU�  _Up�_��Wp5p5\\�5��W3\ 7�5\3�  �����  �?  �?      � �      0            0      0      0�������?�������0      0      0      0      �      �           � ��    �\U  �U5\U5  \U5WU���WU�WU�  WU�WU�  WU�ww�  �����  033 ��  ���U=  |U�U��WU��_p�W�5p5\\�5��W3\ 7�5\3�  �����  �?  ��      � �      0 ��� ���0<�;<0���;�?�ꬳ�:�0������0�����:0�����:0�����0����:� �:� � <�:<  ���� ��    �\U  �U5\U5  \U5WU���WU�WU�  WU�WU�  WU�ww�  �����  033 ��     �  0�  0�  0�0 0� 0�0 0�  0�  0� ��� �� �� �� � � 0 0 �         0? 3    0 �0���� ��: ��?  �?  � �  0  0  0  ?  �3  �3  �<  <0  �  �?����:�:����� �?  � �  0  0  0  ?0�30�3�0�<�<0  �������:�:�����         �?  � �  �  �  �0?�03��03���  ����:�����?��             �?  � �  �  �  �� ���  �<<��  �� ��?�0� � ��������  �  �  �  �  �  �  �  �  �  �  �  �  ���������	����������������      �      �      �      �      �      �      �      �      �      �      �      �      �����������������!��������  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ���������	!����������������      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �      �����������������)��������������������        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        �        ���������������������  ��    ���   �  �     � �    �    < <    0     �     �     �    �    �    �    �    �    �    �     � <    � <    < �     �  �  ?  �   � ?   ���           @           @A @@A@@AQ@A&PQiPV�@�a �i d       �   "  �  �   �	� �%`�$&`�$� �$�H��Hb@%H@%ET	�UU ��             �� ���?���������������?�  �?  �  �  �      ����?<<�������������������3<��<��?��� ��  <<  �  �  �  0 � � ��7�?��3= �� �� � W�2 �? � \�Y�jU����  �?  ?� �[�VT��3�UU?�VUů_iի�Vլ�U1�^�:�Z����쫪�����   �  
? �� �2� ��
 h H  H  J  J. �H.  �# �# �� `= �  � ��� �  0  �3 ���?333�����333����� 0  0  <<  3� ��3�?�            �       � � � ��$��$ �$	H�	Hb@	H@	ET�U�  �
               �  �  "  �$ ��	�`"	(b&�`&�X�	P	V ThU� ��
       �      �"                   H      B      B   �  B    * B    �	     	%  � $�  �(� �  ���`@  ��`@
 H���@� Hb��P� Bb��P"���`P"	��$� 	�$$�	`� %PI	`P�@ 	`PT @	`A  @�   P�    �  V   T%  X  U)   UP�  �RUU*    ���      *       �             �       �!      ��      ��      ��     �� �    `��"    X�`    $�
 �$( �	F� ��	F�   �F�! ���! ���� `�	$`$$` $$`a�X	` �	` PT	�  PA	�   @ V    P X   �  hU  @%  �VPU   �UU�    ��*     �   �   �����
���������������*��   �   �   �   �   �       �       �       �       �       �       �       �       �       �       �       �  �*� �  
�
 �  �
 
 �   (� �   (*  �  
�
 �  ���
 �       �       �       �       �       �       �       �       �       �       �       �       �       �   � �� �� �� �� �� �� �� �� ��   � �� �� ��   �      �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �       �   �  �   �  �   �  �       �   �   �   � �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*� �*�   �   � �*� �*� �*� �*� �*�   �   �   �       �       �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �   �  �       �       �   �  �   �  �   �  �   �  �   �  �       �       �       �6 @ I S [ c k r y        y � � � � � � � �  � ���� � ���* � � �� � ( �
 � 
 �( �� �� �� �� �  ���( �� �
�( ���� ���� �� �� �( � 
 �
 � � �� � �
 ��  ��
 (d��� ��� � � '>Uk������,B[x�����*CZp������.Hb}����9Yz���.Qt�����(@Yu����5Tr����	)	D	_	x	�	�	�	�	�	�	�	�	�	�	�	�	�	�	��� � �� �3 � �7 �0 �́3 � �7 � �́3 � ��5 � �́3 �0 ��5 � � �́3 �0 �7p5 \   �́3 �� ��p5 p   �́3 �  \�5 � �  �́3 �  \�� �5 0  0 �́3 �  \����5 0  0 �́3 �0  W�p�5   3 �́3 ��  W��u�  �? �́3 �� �� W�U�  � �́3 ��� WsU�  0 �́3 ��U�U]U� �0 �́3	 �� �0�U}U�5 � �́3
 �  0�U�5  �́3
 �<  � WU� ��  �́3
 �� �WU� �<  ��  ́3
 �  \U�� �� �|  ́3
 �00 �pU�= �� �W  ́3
 �0�  �WU� 0 ��� �́3
 ��  ���?  0 ��� �́3 �� �0 �p� �́3 �  �0 �pU  ́3 �����? < �0 �pU  ́3 �0 �� �3 ��U  ́3 � � �3 �W5  ́3 �� �3	 ��? W5� ́3	 �
 �3	 ���\5\́3 ����?	 �Wp5p5́3 �	 ��_]w� �\p5�5́3 ��	 �|UUuU= �\5p5�5��3 �0	 �WU�� �p5\5�5́3 ��	 ��U� �p�\5��́3 ��	 �pU�5 �p�W�p�́3 ��5	 �\U�� �pUU�\�́3 ��50 �WU� �pU�W5́3 �?�5< �WU� �pU�5́3 ��5�53 ��U� �pU�̋3  �<p��� ��U� ��U�́3 �\pU� �pU��U�5 ��WUU� ́3 �WpU� �pU��WU�UU5 �_UU= ́3 �WpU� �pU5�_U�Uu5 ���� ́3 �Wp� 7 ��\U \U�U�� �́3 �W5\��5 ��U5\U pUWW�� �́3 �W�W�p5 ��U�\U ��WW�� �́3 �WU�_ �pUU_U ��U]�\
 �́3 �WU� �p�WWU �U�\W �? �́3 �WU� �pu]W� �WUU\w ��� �́3 �\U� �p]uU�  �WU�\ ���  ́3 �pU�� �p]WU�  �WU�\w ���́3 ��U�5 �p]WU�  �_U�\w ��́3 �WUU ��uUU�  �U�\ ���  ́3 ��U� ���]U� ��U�\W �� �́3 �� W��  ��U�\] ��� �́3 �\UW�  ��U�\� �� �́3 ���WU �U�\� �� �́3 ��UU �WU� \5 � �́3 �pUU |UU�W5 �< �́3 �pUU��WUU�W5 �� �́3 �pU��U5 �< �́3 �pU����UU5 �� �́3 ��UU�U��_U � �́3	 � ���U�_U�U �< �́3 �� ��UUW�WU�}U= �� �́3 � �\UU]�U�_U�  ��  �́3 �� ��WU���WU��U=  ��� �́3 �� �pUU? �WU��U� �< ��  ́3 �� �\U�  |U��UU  � �́3 �� �WU  �WU�WU  � �́3 ����  �U� �|U�� |U5	 �́3 ��? pU5 ���_U��? �U5	 �́3	 � \�  ��������� W�	 �́3 ��  \U  ��:  �����U �́3 �  WU �ꪯ�  ����|U= �́3 �� �WU �����  ����:pU5 �́3 ���  W�������  �����p�� �́3 �wv��ꬪ� �����sv� �́3 �|W��ﯪ� ���~�� �́3 �������� �����5 �́3 ������ ����� �́3 ������ ���
 �́3 ����?  0 �
 �́3 �0 ��  ���
 �́3 ��� �́3& �́�&���(d��� ��� � � '>Uk������,B[x�����*CZp������.Hb}����9Yz���.Qt�����(@Yu����5Tr����	)	D	_	x	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�� � �0 ���3 �� �� �� �́3 ��0 �� �� �́3 ��0 �\ �0 �́3 ��0 �? \� � �́3 ���  �5 \� � �́3 ���  p \� � �́3 ��  p \�5  � �́3 � �  \ W�5  0 �́3 � �  \�W�5  0 �́3 �� � 0 \s���   �́3 ��� 0 W]���   �́3 �0� � WU�� W  �́3 ��� � WU�� W� �́3 ��� �WUuU�U0 �́3 ���� �\U�}U �	 �́3 � �\U�  �
 �́3 �� � �pU��   <
 �̅3  � �� < ��U��� ��
 �̅3  p= ��� �WU�50  �0
 �̅3  �� �� �|U� �
 �́3 �W � �WU�  �
 �́3 �W �  ��? �0 
 �́3 �W �0 �� �̆3  �U �0 �� � �̆3  pU �0 �< �?�� �̆3  pU ��0 �� � �̅3  \� ��0 �0 �� �̈3 ?\� �	 ��0 � �̈3�5\5�W�	 ��0
 �0	 �̇3\\p�	 ���� �̇3\\p5 ��W�u�	 �0 �̇?\\\5 �|U]UU=	 �� �̇3\\5\ �WU��	 �� �̇3W\5W ��U�	 �7 �̇3W_�W �\U�	 �� �̇3W5WUU �WU�5	 �\ �̃3\�U� ��U�� �\ �̂3\U� ��U�� �<\� �̂3pU� �pU� ��\\ �̂3�U� �pU� �p_p<�  ̇3 WUU� �\U��_U �pUp5 �̆3 |UU� �\UU�U��WU �pUp� �̆3 ��� �\]U�U�\U �7�Up� �́3 �WsU�U5 pU5�� �� Wp� �́3 �Ws��U pU5\U �\W5\� �́3 ��p��W �U5WU �\W�W� �́3
 ��5�puU_ �U�UU �p�U�� �́3 �� ���5�U� �U��W �pU�� �́3 ��� ���5�UU� �W�u] �pU�� �̆3  ��? ���5�WU�  WU]u ��U�5 �̄3�� ���5�WU�  WU�u �WU� �̃3�� ���5�_U�  WU�u �\U� �̅3  �? ���5�_U�  WUU] ��UU� �́3 ��� ���5�U� �WUuW �U? �́3 ��� ��u5�U�  W� ��� �́3 �? �w5�U�?  W�U5 �́3 � �_5�_U�? �U�W �́3 �� �\5 _U�? �UU� �́3 �< �\��_UU= pUU �́3 �� �\��WUU��_UU �́3 �< �\UU� �́3 � �\UU��U� �́3 �� �pU�_U��UU� �́3 �< �pU�U��WUW� �0	 �́3 �� �|U}U��_�UU �� �́3 �0 ��?  ��U�U�_uUU5 �� �́3 ��?�  |UWU��_�WU� �� �̈3  ��? < �WUWU��� �UU �? �́3 ��  �UU_U�=  _U5 �� �́3 ��?  pU��U��  �U� �� �́3	 �\U= WU�= �WU  ��� �́3	 �\U �U���� �\U � �́3	 �W� ��������  pW5 �	 �́3 ��U7����  ���  �U5   �́3 �|U=����  ���� pU�  � �́3 �\U����  ���� pU� � �́3 �__��Ϊ  ��ꪯpW�  �? �́3 �_�ͪ��� ���:��p�� �́3 ����� ���������= �́3 �\f��� ���:��� �́3 ������ ���ꫪ �́3
 ���� ����� �́3
 �0 � � ��� �́3
 ����  � � �́3 �� �́3& �́�&���H��� � 7ĩm�� ��������� �ũ~��,��������� �ũ���8��������� �� ���P��  ��� Ј�� �����R��  �h`TRY AGAIN$GAME IS OVER$PLEASE$ٺ��HZک �	��������ʀ��ˀ����Ȁ��ɀ������ �  ���zh`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���آ t ���d���� � �����������  ��� � �� � �� �ύ& ��"  7ĩ�� d
�� ��L`�       ^�n�~�������������������.�>�N�^�n�~®¾�����������.�>�N�^�n�~ÎÞ�  ��$�                                                                                                                                                                            �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  HZ�H�@��m��������8��HJJH

�zh8����m�� ����ɪ�8��i0��i ����h�zh`H�i0��i ��_�����8������h`H�H�H�H�H������ k�h�h�h�h�h`�H�Z�ڮڦڦ� ��8��JJ�8���� � ����� ����h�h�h�h�z�h(`Hڭ  �� �������%���h`������������{}~���������������������H�  ����h`H�Z�ڦڦڦڮ	�
��`���a�� �Ü	� �  q�-  y���� �����iɠ���iɠ������h�	h�h�h�h�z�h(`   Hڪ)�JJJJ Ŋ) ��h`HZ� ��$�#�0i��:8�0��A08�7�i �Ȁ�zh`�H����� L��Z�H�H�H�H�H�H�H��H��Hi�H�i �H ��8��JJ�8�����m��i ��������?������6� ��ȭ��h�h�� �������� ��m��i ���hh� h�h��0�� �����������ݬ�������
�h���h�	��h�h�h�h�h�h�h�zh(`�� �2��.HZ�Z�Z� ���������
������� �h�h�zh`�H�Z�H�H�H�H�H�H �à �ȍ���-�i��i �� � y�����m��i � ����h�h�h�h�h�h�z�h(`� �#��H���hH�Z�ڦڠ �������Lv�L�L~���� �Ȁ����LYȥH�H�Z�
�������������	8������	�� ��������*�e��i ��e��	i �	� �������	���8����	��������
�8����������������8h���h������
�������	��������h�h�z�h`ڦ
����	��.������`H�� �� h`�  � `H�Z�H�H� H�H�H�H�H�H�H�H�H �Ì�JJ�NN� ����:����:�ȱ���:����:��8�����h�Hڭɀ�
��8�
���Hȱ�����he��e������� ��h�+� � � qʍ �� �3� m������ q�ڮ� y�����
������P��r� m�����m ����8� � �8� �	� �m ��H q� y�h��,���� qʍ �� �� � q�ڢ ��� �� ������ �L.�h�h�h�h�h�h�h�h�h� h�h�(z�h`Z���z�`Hڦ��	���Q����h`�ڮڮڍZ�)���=%ˑȱ�=(ˑ8����Z�JJ�����

������	��
�M��z�

�����JJ����z��ȭ�h�h�h��h`?���H�Z�H�H�H�F�H� �

�ȱ�z��Z�H��hHڍ ǭm����m����hhh�h�h�h�z�h`��d % 4 O B 
 z  0 
7 p 
   � � ���7�kĺ���ŀŕ������vǀȗȦȭ�q�y�,�                                                                                                                          �L��L��L��L��Li�L��x�d�# X � Ω�)��& ���X � �ĩ�� � ;Ωύ& ��� � "Ω���� � O��H� -Щ( Щ���  � f΀� �� �ͥ�
�	�����ѭ��
 �ĭ���d
��L��.ͅ�/ͅ   *Э���
 Ѐ �� �ͥ�����N�O�P�T�V�V�V�V�\�g�r�}�PAUSE$F�`` !�`�` �`�`H�� �h`H�� �h`H�� �h`H�� �h`H iΥ����� � $�dh`H�  ��	�J�IL���������������h@�Ѝ&  ��h�
h�h�h��H(L}�H�Z�' )������ � 	褐�# �$ �% z�h@H��)	 �&   ��ύ& h`H��)	 �&  ��ύ& ��Hh`H��)	 �&  ��ύ& h`H��)	��&   ��ύ&  �h`L̀H�Z� �	�����$���%�� � �Ω���I
��R���S�� ǩ4���� 'Щ������ �ũ �z�h`H������H �� ��h`ڮHڢ ��
��
H��i�h��H�mH��H�(` 0 < �� <        � ���?�?  �0��3�3��3�  L>ѭ �΍L>ѭ �΍L>ѭ�0	� �΅�� �΅L>ѭ�0	� �΅�� �΅L>ѭ�0	� �΅�	� ��)�L�͠ ��	� �Α�ȱ �ΑL>Ѡ���ݠ�٠�ՠ
�Ѡ�͠��L�έ���H�H�Z��0� ��kh�h�` �L\�L�L��L��LB�L��L0�L��L
�L��LG�L-�L��L��L4�LX�Hڦ���d:����h`�Z��Z����m����z��z�`H�Z��:
���Ѕ��Ѕ���
 B�m����Mz�h`N�\�#Hک �	���� \ЭM
��*���+�� �� ��h`H�	���� ��������������� G� 
՜������� k� n�h`H��



���



�h`H�Z��:
���Ѕ��Ѕ���
 B�m���M�z�h`H�Z�H��



��� �

���͌�
��͌�&�H����@��)�JJJJ����)�������+������)�JJJJ����)������������ �� ��h�z�h`H�Z���L�ӭ�������� �ԭ��L�� 5ծ������,�����~�	�(�,� �~� 0�ʀ��~��Ȁ��~� 0� 7�L7ӈ�� �ԭ��<�������� \ЭM��c�$�� �'�����+��*��������=L7�L5�L%�Lӎ��� c�,LM� �� �ێ������������M � �Ѐ����� ���� �ԭ��`�	���� �ԭ��K� ���� �ԭ��6��2��� �Ԁ$�����H����  �������� �Հ�T 
խ��H�( 0Э���������� \ЭM�$���� \ЭM������M � �М�� u֜�z�h`�������  �H8�� �HLb�H�Z�Y�#�����G0E:� BШ������)?�(������!���#��  Ԁ Ԁ AԀ gԘi����z�h`H�Z����������M �z�h`H�Z����������M �����M �z�h`H�Z����������M �����M �z�h`H�Z����������M �����M ����	�M �����M �z�h`H�Z��������� \ЮM��ԍ��#�8��ԍ��8� Ս� �


��� ��z�h`               Hڭ������� �Щ �	�~
������� ��h`H�������� ��h`H�Z��� �	���T0R:� BЪ�������� �н�)?�8�

��}��Z���[����Ȁ� Ǌi���­}��}��}z�h`H�Z�����;09:� BЪ��)?�!�������� ���� ���� ���� �Њi����z�h`Hک�	��)�:
����������������� �� ��h`H�Z �ĭ����������� \ЭM����� �� eـL1� �ک���  �� ��z�h`H�Z����)�JJJi���:� BЪ����)?ͺ���ݔ���ݕ��i��٩����D��������8���0�������������� r� ؜� �� Gս������  �z�h`����������� \ЮM��8��ԍ��8� Ս�����:� BЪ��)?����������i����߀
��)?8��� `H � �� �ש���  �< 0� � �� �ש���  �( 0�h`Hڭ�):
����������������� �Щ�	 ��h`H�Z�������� �Э�):��y؍�y؍� �	�� q� ��z�h`  H�Z��):

����}A؍���}Q؍� �����z�h`                          Hک �	�$����$���%�� ǭI
��R���S���T��� ǩ<����H q� �ũl� ���h`H�� q� �ũ& ŭ� q� ��h`H�Z 7� a؜�2�� � �������& �-���.�� �ȩύ& �  ���	��z�h`H�Z��)�� ��)
����������Sٍ�\ٍ �z�h`$-D[d[D-ZC:CZqzqH(1H_h_H1^^G>G^u~uH�Z �ĭ  ������� �Ģ��)����	��LYک�	���������Bٍ�Jٍ ǽ�)
����������Sٍ�\ٍ� �	 ǭ  ���G���a���	���� dڀt����  � �ĩ�	 ǩ�	���������Bٍ�Jٍ ǜ�Lk٩���  � �� ����
��)���L�٢	�既��  � �� ����	�
��)���L�٢ ����  �z�h`H�Z��)���0�)��%������ ?܀ �܀ J݀ �݀ �݀ ހ �z�h`H�Z�H��



��� �

���͌�
��͌�&�H����@��)�JJJJ����)�������+������)�JJJJ����)������������ �� ��h�z�h`�������  ��c����Lb̢������  � �� �J���J��)	��&  	��ύ& Le̩�)	��&  ��ύ& ��JLh�H�)	���h`H�Z �ة���  ��	� �����  ���� 0�κ�� و��)� �轱)��	������.������ ٩���  � �Ġ(��� 0Э  ���񩂅�  �z�h`H�Z�`�����
��������� �z�h`H �� ܩ���������� �� �� �ĭ����m �� �� �Հ� �ĭ�́���͂�ԩ���������� \ЭMл���� \ЭM��
������ 
խ������� 
՞�����  h`H�Z�H �� ܩ 0� �՞���:� BЪ����")?8���	��)�	�)?���)����i���� �ө 0� Gթ���  �h�z�h`HZ� �� ܩ���������� �� �� �ĭ����d �� �� �Հ� �ĭ�́���͂�ԩ���������� \ЭMл���� \ЭM�
��������M � �О�����  �zh`H �� ܞ����Hi��H
�(��(�H� 0Щ���  � k�h`HZ� �� ܩ���������� �� �� �ĭ����> �� �� �Հ� �ĩ���������� \ЭM�˞� �� ׽�8����0�������   �՞� �� G՜��zh`4HZ� ׽������� �Ќ��

��� �	������������������������ ǩ���  � 0���Ȭ��
����À� ǩ( 0� G��zh`HZ� �� ܩ���������� �� �� �ĭ����j �� �� �Հ� �ĭ�́���͂�ԩ���������� \ЭMл���� \ЭM��
��
������� �M � �О�����  �zh`H�Z�������X�������J�� �������� ���	��	���� �ĭ��� \ЭM�������������  �z�h`HZ� ���0]�[:�)HZ���	�O��)?���!��#�����}��	�/������ �!��)?�!��� �����:�����zh`HZ� ���0]�[:�!HZ����O��)?�!�����}���7������ �)��)?���!��#��� �����:�����zh`H��� \ЭM����� \ЭM���������8�-��ͺ�$��



�����



�ͼ������h`HZ��H)�JJJJJJ�h)?{ᝓzh`��@ H�H���� �� `� `��h�h`H�H���� � `���h�h`H�Z�H:�����  ����� ������ `���h�z�h`H�Z�H:�����  ����� ������ `���h�z�h`H�Z�H��



����



��i���8����i��	�8������������^���*��������������:�ｕ���������:���� \ЭM����� \ЭM���������h�z�h`H�H���� �� `��h�h`H��)��ɀ�� ��� ��� &�� 6�h`H�Z���s �խ�H���j�� �ө���:� BЪ��"��)?��8�
��L�������   �ӊi����Ό �ӭ�еh�� �� Gխ����� �H0� 
Հ
����  � 5�z�h`�������:���������������HZ��)?8�
�� ���������ȱ��zh`H�Z����������� ��H8��0�H��H r� 
թ 0ЭH�����  ����z�h`H��~ 
�h`Hک���  סּ���������� \ЮI����M�'�M � �� 
���4���� �ح�Ͱ� ���h`H�������������0 \ЭM��U��Q�������	� \ЭM��:��6�������0� \ЭM������������ \ЭM������M � ��h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   L�L��L`�LI�L�L�� �P�Q�R �� �� � � � � � � � �* d�d�� ����d�`�Q����y� ��r� �s�  D��y�y�t� R�R������ ��� ���  ��憥�Ł� ��P���J�Q����]� ��V� �W�  ��R����k� ��d� �e�  ���]�]�X� ���k�k�f� ���� �� `�`�S�T�VȱT�WȱT�XȱT�YȱT�Z)
�����[����\�Z)0�`ȱT�����ȄSd]d^�X� �L��_ l�� �
�T� �d_��Ȅ_dS���o�p�rȱp�sȱp�tȱp�uȱp�v)
�����w����x�v)0�{ȱp�����Ȅodydz�t� �� �Q� ��)��	���Rd| ��`�|�}�ȱ}��ȱ}��ȱ}��ȱ}��)
�������������)0��ȱ}�����Ȅ|d�d���� к� �R� ��)��@Ы���Qdo R����a�b�dȱb�eȱb�fȱb�gȱb�h)
�����i����j�h)0�nȱb�����Ȅadkdl�f� й�m ��� �
�b� �dm��Ȅmda����
������轐������Tȱ��U`��
������轘������bȱ��c`H�Z�Y)?	@���Y;��%����^�[��Z)@��J������`�8��`��Z)0�`Ȅ^�[����^�Zd^��� z�h`H�Z�g)?	@���g;��%����l�i��h)@��J������n�8��n��h)0�nȄl�i����l�hdl��� z�h`H�Z�u)?	@���u;��%����z�w��v)@��J������{�8��{��v)0�{Ȅz�w����z�vdz��� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ƈ��d���� z�h`� `� `H�Z���������������)?
������轓���d� %�z�h`d��* d�`������ȱ���ȱ���ȱ���)
�������������)0��Ȅ�d�d���� �d�`H�Z�����L�󥋅���;��)����������)@��J��������8������)0��Ȅ������Ɛ��d���)����)����
�@����������( ��ŕ��* ��捥�Ō� %�z�h`H�Z�  l�  ��dSda��_�m �� � �� �� ����Pz�h`H�Z�Q� ��R� �d���)?Ŝ�D�� �>��
�����p����}����q����~dod|� �Q�R��)�����R �����Q R� ��z�h` ��b� ��b� �H�b� ��b� ��b� ��b� �<�b� �b� q�b� �H�b� ��b� ��b� ��b� �<�b� ��b� ��b� ��b� �<�b� ��b� ��b� �<�b�     � ��b� ��b� �H�b� ��b� ��b� �H�b� ��b� �b� �b� <�b� �b� _�b� q�b� �<�b� ��b� q�b� �<�b� ��b� �0�b� ��b� ��b� �`�b�     ���"���"�}�"�.�"���"�.$�"���"���"�T�"���"�T�"�.$�"�}�"�T�"�.�"��"�.�"���"���"�T�"��"���"�     �T$�"���"�}�"�.�"���"�}�"��$�"���"���"���"���"���"��$�"���"���"�T�"���"�T�"�T$�"���"�.�"�}�"�.�"�     �T�"�}$�"���"���"�\�"���"�}�"���"���"���"�\�"���"���"���"���"���"�:�"�\�"���"���"�\�"���"�T�"�}�"�T�"�T�"�}�"��0�"��`�"�     � q��� q��� ���� q��� ���� ���� �(��� q��� q��� w��� d��� qP���     � ���� ���� ���� ���� ���� ���� �(��� �
��� ���� �
��� �
��� �
��� ���� �P���     ��(���.(���}(���.(���.(����(����(��� �(����(���}(���.(���}(����(����(����P���     � �,�D� ��D� ��D� ��D� ��D�.,�D� ��D� ��D� ��D� ��D� �X�D� q,�D� ��D� ��D� ��D� �B�D�     �.�D� ��D� ��D� ��D� �X�D� ��D� ��A�  ,�D� ��D� ��D�  ,�D� ��D� ��D�  ,�D� ��D� ��D�  ,�D� ��D� ��D�  ,�D�     ��,�3��,�3�\,�3�\,�3��,�3��,�3�\,�3�}�3�T�3�.�3��,�3��,�3�\,�3�\,�3�     ��,�3��,�3�\�3���3��,�3��,�3�  ,�3��,�3�  ,�3��,�3�  ,�3��,�3�  ,�3��,�3�  ,�3�     �\�3��$�3�\	�3�\Q�3���3�\�3���3��6�3�\	�3��	�3�O~�3��	�3�O	�3�\�3�     ��~�3��	�3��	�3��l�3��	�3�O	�3�\�3��~�3��	�3��	�3��$�3�     �����$������$��:��\���������$�����O��  $�����\	��:��\	������	���$���$�����:��     �\�����  $���l��  $���$�����:��\�����  $���$��     � ��� /(��     � %w� #w� %w� %u� #u� %u� %s� #s� %s� %q� #q� %q�     � w�"�     ��"�     �����T�������T�������T���     �  H �� �� �� �� �� �� ����.�@�T�h�}�������     � *��� *"���     � �x� � _� x� �z� �|� �     �  � � � � � � �. �} �� �\ �� �� �� �� �� �     � �{� �{� �{� �{��{��{��{�}{� {� q{� d{� _{�     �����/�B�]�h�s�������������o  �?  �O  �   OMLKJIGFECAOMLKJIHGFECA/    o  �O  �   O  �?  �/  �   o  (�   O  (�   _  �_  �   �o
5��o
5��o
5�   �o   �/�  ��_�  ��_�  �   �/�  ��O�  �   �O�  ��/�  �   �?�  �   ��0�@�E�J�����	�
	�
	�
�
�				


�
	 � �����������������W���  ��  _���  C���  {���  �����  ��W�  ��)�  w�������=�����E�w�������������E�          �� ���