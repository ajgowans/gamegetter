UUUUUUU TUUUUUUUUUUUUUUU    @UUUTUUU UUUUUUUUPUUU PUUUUUUUUU    UUTUUUU UUUUUUUUUUUU   UUUUUUUUUP   UU UUUUUUUUUUUUUPUUPA  PUUUUUUUUU   UUUUUUUUUEUUUUUUUU   PUU  UUUUUUU   @UUUUUUUUUUU���UUU   TUUU DUUUUUU    UUUUUUUUUUU ��_U @UUUUUUUUUUUUUQ   @QPUUUUUUUUUU5 �O�UUUUUUUUUUUUUUUUU      @UUUUUUUUUU5 ? �WUUUUUUUUUUUUUUUU  P@UUUUUUUUUUU5 � �WUUUUUUUU@U @U    TUUUUTUUUUUUUUU� �J�_UUUUUUUUUU      UUUUUUUUUUUUUUUUU����_UUUUUUUA       UUUUUUUUU�WUUUUUUU�  ��UUUUUUUUU@    QUUUUUUUUU�UUUUUUUUU# ��UUUUUUUUUU  TUUUUUUUUUU�WUUUUUUUU�  �UUUUUUUUUUUPUUUUUUUUUUUUU�UUUUUUUUU= ��UUUUUUUUUUTUUUUUUUUUUUUU�UUUUUUUUU�� ��WUUUUUUUUUQUUUUUUUUUUUUUU�WUUUUUUUU�3��_UUUUUUUUTUUUUUUUUUWUUUW�}UUUUUUUUU0��UUUUUUUUUUUUUUUUUU�wUU���WUUUUUUUU��UUUUUUUUUUUUUUUUU���UU�����UUUU���� ������������������������������������� }�������������������������������������D�U���������ꪪ����ꪪ�����������ꪪ���D�_������������������������������������.D�_���������������������ꪪ�����������>UU�������������������������������������:UUի�����������ꫪ����������������������TQԯ
�����������������ꪪ�����������뮮�PAU} ������������������������ꪪ�������CTU�U����������������ꯪ�������ꪪ���T�U 𮪪�����������ꯪ����몮����ꪪ�/U�W����������ꪮ���꭮����������������DU�[����ꪪ��������������ꪪ����ꪪ�ꪾpUAm ���������������z����������������UA}@կ��������������ݪ��������ꪫꪺ���VU��U��������ꪪ������ꪺ������������ UU?T?�������������jժ�꺪�ꮫ������� �oU>T� �������������������몮��뮪���  �U<T� �.���������^ߪ����������몪�?   ��@�P�/�+�����ꫫ��V�����ꪯ������CUU�P� ����
C���������֪��몮����ꮪ>PUUU�/W� �����CU𪪺���֪������������TUUU�W�  ���� T������gݮ������������� @UU�W�  ����@ ��ꪪ�g�����몪�����/  @UU�W�  ��0 ��������g����������ꪪ�   PE�W� ��?���������v�ꪪ���ꪪ���P   �W� ��?���ꪺ��U����꾪������;TP   �W�> �����������]^�꾪��������UU   ��U�� ���ꪪ���^y������������ UUU ������<���ꪺ����_m������������:PU ����  �8�𯪪�����[u��_�jU�V�> ����  �>��� ������WU��jU�UU���  �����>  �:���  �ꪪ��u��U�jVPe���  �����:  �����������������U��jU ԯ� �������  �����������꺪����yU��V @�ꪪ�����������������ꪫ몫�����^U�*  Ծ�������ꫪ�=����������������e�WU�j��������������������﫺�������UVVUj���@�����꫺��TU������ꪺ����zUYUeU�j E������������?TU�����«��������[ZUUU�j
  ������ꪪꪮ ����������������oUUUU�j�
`�������ꪺ�� �����0��������UUUUU�jV������������ ������  �����WUUUUU�jVUկ�뮫������ ���?��? ������UUUUUU�jV��������������??��* �����_UUUUUU�jVU������������﮺��è�  �����U��U�V�jVU�����ꮺ���������� �*�𺪪UUUUUi�jVU�������뮮�������� �. ���WUUUUUU�jVi��������������
 �� ����UUUUUUU�jVU�����������������
 ��  ��_UUUUUUU�jV����몪���ꪮ������
 �
  ��UUUUUUUU��jV�����������������
  �/ �~UUUUUUUe��jV������몿������*  �23,\UUUUUUUU��jV������������/�� �TUUUUU�VU�������������������몯��  (�
 HUUUUUUUU���������믯��몺�����/���� TU�UU�UU�������꾻��������������#  �� PUUUUUUU������������������������:b TUUUUUU��������﫯���ﺪ���������("��A TUUUUUU�z��������������������?��UD UUUjUU��V����������������꿪��請2 �pEDUUUUUeiV�����������뫺����몪��È�\UUUUUi�������������������ﺺ��GU UUUUU�U����꿮�����������������.UQEATUU�V�U���������﫪ꪻ���������3HUDQTUUU�����������������������꾪�.�TUAUUU���������������������� EUU@QU�����������﮻�������꫾�����rDQUQT��������������������뾪��뺪�NUUQTA���������������������껺���PTT@������������������������������Q UUD������������������������������STUU����������������>���������������*�ETUU#��뫫�꿪��������������뿮�������<UT �����������������������ﾪ���.�0PP�?� ������﫯����(��������뾻���������*�,���������������뿫�����������
����+��������������������������������������� ����������,����﾿�����������"� #��*������������������������������*����.���ϸ����������/����������������������������꺿�������������ﻺ�����������￪���Ȩ����������������������������ʠ����*�"������>������������뮺ﮯ���*�8Ϗ/���8�*�．���?�����������������������"���((���"/;/�����뿾��������꿪���<�,����+�������������������������뫺ﯮ�
ʪ������������;�������뿮�����������?�����?��ȿ���������������������������Ͼ���̸ྫྷ��>�(��������������������������;�����>�����������������������������������;���������������������������������?������:����������﮾��������﫿���?��?����.˪ο������������������������������ϼ�󫈊?������������������������������������������?������������������������������?����/�������������������������������?���������Ͽ��������������������������������������?������������������������������������>�����������������������������������������?�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ﯿ��������������������������������������������������ﯿ�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������￿���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������￿��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������￿����������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 P                                     PUU                               @UU PUUU                               UUUUUUUUU                              UUUUUUUUU                              UUUUUUUUU                              PUUUUUUUU                              PUUUAUUU                                UUU  @U                                                                                                                                                                                                            @UUUUQ                                 @TUUUUU                                PUUUUUUU    UUU                       @UUUUUUUU  PUUU                       @UUUUUUUU TUUUU                      PUUUUUUUU QUUUUUUU                    PUUUUUUUUUUUUUUUUUU                  @UUUUUUUUAUUUUUUUUUUU                 PUUUUUUUUUTUUUUUUUUUUU                 PUUUUUUUUUTUUUUUUUUUUU                 TUUUUUUUUUTUUUUUUUUUUU                 UUUUUUUUUUUUUUUUUUUUU                 QUUUUUUUUQUUUUUUUUUUUU                 TUUUUUUUUPUUUUUUUUUUUU                 UUUUUUUUUUUUUUUUUUUUU                 UUUUUUUUUUUUUUUUUUUUUU                 UUUUUUUUUUUUUUUUUUUUU                 UUUUUUUUTUUUUUUUUUUUU                 PUUUUUUU@UUUUUUUUUUUE                   UUUUUUU QUUUUUUUUU                    PUUUUUD  PUUUUUUUU                       PUE@   @UUUUUUU                                PUUUUU                                   PUU                                                                                                                                                                                                                                                                                                                                                                                                                                  @UU                                    @UUUU                                @UUUUUUUU                              PUUUUUUUUU                             TUUUUUUUUU                      U  P @UUUUUUUUUU                     TU@U PUUUUUUUUUU                     UUUQU PUUUUUUUUU                     @UUUUU @UUUUUUU                       PUUUUU @UUUUUUU                        PUUUUU  TUUUUU                        @UUUU   PUUUUU                          UUUU     UUU                           TUU      TU             @UU           TU                     @UUUU                                   @UU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUQUUUTUUEUUUTUUEUUEUUQUUUEUUUTUUUQUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUQDEUUQDUTQTEUUTQTEUEUUQDUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUPUTTUUQUPUTTUUEUAUQQUUEUAUQQUUQUPUTTUEUQQUUEUQQUUUEUDUUAUEUDUUAEUQQUUUUUUUUUUUUUTUTETUTUTETUUUUUTUUUUUUUTUUUUUUUQUUUUUUUQUUUUUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDUUUUUUDUUUUUTUUUUUUTUUUUUUUDUUUUUDUUUUDUUTTUUUTTUUUUUDUPA@TAQUPA@TAQUE@QEUE@QEUPA@TAQUUUTAUUTATTUPUTTUPUUUTAUUTQUUUUUTQUUUUUUPEUUUUUUPEUUUUUTQUUUUUUUTUUUUUUTUUUUUUUPUUUUUUUPUUUUUUTUUTUUUUUUTUUUUUUPUUUUUUPUUUUUUTUUUUUUPUTUUPUTUUA@UPUATA@UPUATPUTUUTAP@DQTAP@DQQ@EQ@ETAP@DQUU@UQ@UU@UQ@UUUUDU UUUUDU UU@UQ@UDUUUUUDUUUUUUUUUUUUUUUDUUUUUTUUUUUUUTUUUUUUUQUUUUUUUQUUUUUUUTUUUUUUUUU@PUUUU@PUUUU @UUUU @UUUU@PUTPPPTPPPUP@@@UP@@@TPPP  T @A  T @A  PU    PU    T @APTUUTPTUUTAPUUUPU@PUUUPUPTUUTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�������������������������������������������������������������������������������ꫪ�������������������������������������ꫪ�������������������������������������ꫪ�������������������������������������ꫪ��������������������������������������
                                    ��
                                    ��
UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��
UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��
UUUUUUUUU��VUU��������ZUUUUUUUUUUUUU��
UUUU��UUUeUYUUYUUUUUUUeUUUUUUUUUUUUU��
UUUUYUVUUe�YUUZUUUUUUU�UUU��ZUU��ZUU��
UUUUVZYUUeUYUUZUUUYUUU�UUU��YUU��YUU��
UUU��jeUU��VUUZYUUfUUe�UUU��YUU��YUU��
UU������UUUUUUZfUUYUU��UUU��YUU��YUU��
UU�UUUU�U��VUUZYUUUUUe�UUU��YUU��YUU��
UU������UeUYUUZUUUUUUU�UUU��YUU��YUU��
UUU��jeUUe�YUUZUUUUUUU�UUU��YUU��YUU��
UUUUVZYUUeUYUUZU����ZU�UUU��ZUU��ZUU��
UUUUYUVUU��VUUZUYUUUeU�UUU��ZUU��ZUU��
UUUU��UUUUUUUUZUYUUUeU�UUUUUUUUUUUUU��
UUUUUUUUU��VUUZUV����U�UUUUUUUUUUUUU��
UUUUUUUUUeUYUUZUV����U�UUUUUUUUUUUUU��
UUUUUUUUUe�YUUZ�����VV�UUUUUUUUUUUUU��
UUUUUUUUUeUYUUZ�����VV�UUUUUUUUUUUUU��
UUUUUUUUU��VUUZe����ZY�UUUUUUUUUUUUU��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������������������������
��������`UUUUUUUUUUUUUUUUUUUUUUUUUUUUU(��������
`������������������������������ ������
`������������������������������(������
`������������������������������(������
`������������������������������ �(
`�����������������������������蠨"�*�""
`�����������������������������蠨"�(""
`�����������������������������蠨"*�(""
`�����������������������������蠨� "
`�����������������������������蠪������
`�����������������������������萪������`������������������������������`UUUUUUU	`�����������������������������耪������`������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `��������������������������������       `��������������������������������       `�������������������������������< ?     `������������������������������        `�������������������������������3 ?     `��������������������������������       `��������������������������������       `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `�������������������������������       `�������������������������������       `������������������������������� ?     `������������������������������ �       `������������������������������ < ?     `������������������������������ <       `������������������������������ <       `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `�������������������������������       `������������������������������� ?     `�������������������������������       `������������������������������� ?     `�������������������������������       `�������������������������������       `��������������������������������      `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `������������������������������         `�����������������������������耪����� `������������������������������YUUUUe
 `������������������������������`������	 `������������������������������    �
 `������������������������������`���*�	 `������������������������������`�VUU��	 `������������������������������`bUUUU�	 `������������������������������`bUUUU�	 `������������������������������`�VUU��	 `������������������������������`�����	 `������������������������������`�*���	 `������������������������������`�*���	 `������������������������������`������	 `������������������������������`�ZUU��	 `������������������������������`������	 `������������������������������`�UUUU�	 `������������������������������`�UUUU�	 `������������������������������`�eeYY�	 `������������������������������`��Z�V�	 `������������������������������`�UUUU�	 `������������������������������`�UUUU�	 `������������������������������`V�Z��	 `������������������������������`XUU%�	 `������������������������������`�U�
�	 `������������������������������` �* �	 `������������������������������` `	 �	 `������������������������������` � �	 `������������������������������` � �	 `������������������������������` `
 �	 `������������������������������` �	 �	 `������������������������������` h& �	 `������������������������������` �) �	 `������������������������������` h& �	 `������������������������������` �) �	 `������������������������������` h& �	 `������������������������������` �	 �	 `������������������������������` � �	                               �    �
 �������������������������������`������	 �������������������������������YUUUUe
  �������������������������������������                                                                                                                                                                     �������
                               �ZUUUUUU�                               ���������                               �
      �                                                                       <<��                                 <<?��                                 <<?��                                 <<���                                 <<���                                 �?���                                 ���                                                                       �
      �                               ���������                               �ZUUUUUU�                                �������
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    H�@�� �d��� ��� � �t ���u �u �s �t �r  �ʭu �r� ��u �� ���� �� ѩ�� ���� ��� �u �u �s �t �r �d���  ��Θ Θ �� �s �� �r �� �� �f �ʭ� �D0 ѭ� �� � ����� �� ѭu �s ��� �t �r �d �ʭt i�t �r  �ʭ� �r �f �ʭ� 8��� �r  �ʭ� �� р����b  �ܩ( 9�h é�y �� ��w ��b  �ܹ�ꍃ ȹ�ꍅ ȹ��r ȹ��s  � ��ȹ�� 9� ��� ��w �����y и�
 9� �ũ��h ��\  i�H��{ ���h � �\  i۩� �  é�y �\�r �\�s ��� ���  ��ڢ` ����\�r �\�s ��� ��� ڢb ��� ���y з �ҭ j�� � П�{ І���h ��\  i� Ü� h� �� �@�� �  �� �ũ 9� d© Ll� �( 9�H�@�� ��� ��� ��r �o�s ��y �h�z �  (ɩ�� ��� ��r ���s ��y �j�z  (�h� 9�L4ԩ@��  é�r �s ��� ���� �* � �ӭ� �r �� �s ��� ��� �p �ʩ 9Ѯ� ���͗ 
Η �Щ 9ѭ� � �%��r ���s �� i Щ�r �x�s � � �©d 9ќ� L.©@��  é<�s ��r �!�� �� �x ��� �t �ʩ< 9ѩ�� �t 1˩ 9� ��r 8�(�r � �	�!ݍ� �ة( 9� �� �ө�r ��s � Щ�r �2�s � Щ�r �K�s � Щ�r �_�s � Щ�r �x�s � Щ�r ���s � Э  ��� �ϩ� 9ѭ  ��� �ϩ(��  �� d© Q�L� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              � ?�       �  ��_�� ��ޭ�
  �     �      �=     �W�   �]]�� ��������   **        ?         ��         pU       ����      ��W��   �o���f�3 ��������������������?    ��       ����        ��           0              �              W            �U            �U�           �W�W?         �������      �������Z��  ����*����j����꺮�����꺮����ꪮ�����ꪮ����������������?      ���           �����          ���?           �?                                                          �                    p5                    |�                    \�                    �_                  ���                  |���                  ת�^               �������             ���
�����         ���Z����������     ���z��  �
  ���j��   ��z�����������������������������������>����ꪪ����Z��������꼪��ꪪ����ꪪ����������������������������        ������                 ����                  ���z                �����?                \�����                ������                ������               �����                ���:                  �?�          �  p  \5 ����eY�eY�����f�Z�p�f���pYep��pYe�W� �?       � ������>;�����)�b�/���Z�<�������0�� � ; < <     ��   �� ��� ��_�������?/�����/����+$ 
�%h�
��?
 ��� ��=��?�� �?�� ��� ��+� �����/�� �, P�,�����¯>����� ? �  TUUUUUUUUUUUUUUtUUUUUUUUUUUUUUTUUUUUUUUUUUUUUT           T @   @     T @    T   @  T U       @   TU          T     @      T     P       T        @   T        P    T            T    @       T    @        T            TU          T PUU        T            @T            T            T           @T        @   P T        @    T        @    T        @    T        @  @  T        @  @  TU       @   T          �T @         T          �T  @         T  @     @   (T       @   T       @   �T       @   (T       @   �T   @    T   �T          T         ��TUUUUUUUUUUUUUUT      @   ��T    P     ��T    @ T   ��T    U    ��T          ��TP         ��T         @��T         @ ��T         @  �T         @  �T @        @  �T     PU  @  �T      @  �T
   P  @  �T
      @  �T*   �
 @ �T*  P �"@   �T"   ��@    T"   (�@  P T(   ��@   TT* @ ��*@    T� P ��(@    T(@  �"
@    T�B  "�
@    T�@ ���@    T*@ ���@    T(@ ��"     T*@U  �
     T*        PU PT*        @  T*      P @ T
       @   T
       P   T PU       T  @U      TU    P   T       U   T            TUUUUUUUUUUUUUUT            P T PU @      @ T  @  @UU@T   T     T   @    TTU   T�@ T  �
  *  T  (�  �
  T ���  �
  T ��� P�*  T �*�B  ��
  T ���   �� @ T�"�TU �� @  T "
@�� @  T �BQ ��   T  P  P��   T   �@ (   T  ��J  @T@UU�*
   T    �"
   T    P �PP T    @��@ T TUU�� TT@ATP      @ U T   PP       T �*@A  �   T ��  ��  PT *�T�� T *
 �*
 T@��
  �
 T �� ��
@T P��
 ��
P T @ � P��B T @ � @!�@ PT     ��P@T   U��T TP  @P @T@  P @UP TUUUUUUUUUUUUUUT   @ @ �T @A  U@ �T @@  � @�T*@@  � �T�@@@ ��
P �T�@@@ �*
@ �T�@P@P ��
@�T�B@U���( P�T�B  ���* @�T�B P��*� @@�T�
 @���� @@�T�
 @����@@�T�
TU����
@ Q�T�* ����( A T�* ���� UT�"P@���� E T*� T����D PT��
@@���E T��
P  �*�A �T��
��T���A@�T�**��B���A�T��*��B���BP�T��*��*
��B�T*�*���
���T��*��*��*E�T��
�*��@  AA��T�
P����@@AP�*T�����@��T�����@ ��T�
U����@@(�T�
@��*@@���T�( �� TT���T�* �* ���T�
  UD�*�T
 QP PE����T PATUP A����T@    P@����TUUUUUUUUUUUUUUtUUUUUUUUUUUUUUTUUUUUUUUUUUUUU� ��> �� �� �  �? ��  ��  �
 �?  ��@� �� �  ���� � ?��@� ��? ������ �����p� ��? � ����   � ����� p+ �� � ���  @��� |^�� |?  ��7 �W�? �?  � ���; |  ��7 ���? �?  � ���* �����= �?� _��� �� ���� �= �� ����  � ��W� �}   � �� � �= ��  � ��   ������������������������������������������������_U��W�U�_UU�WU�W��U��WUU��  �> �    ? ��  �� ��
 �    � ܿ �� �� �� |� |? �� ��� �� �� |� |; �� ��?  �� � W W �/  �?  ߿��? �? ���?  �� �?  ������� ��� �?  ����������0 ������� ����  �������  @  �   � � � �� �?  p @������������������������������������������������VUU�W�U�W��W��UU�_U��������������������� ��� �? � ���?   ���? � ����?  ����� �: ����   ���� �: �����𪪪�� �� ����  ����ê� �:��������>����ê��� �����ê��:��j�:��j�ꬩ������� �����ê��9k�V�:��V�ꬩg���eU�  ��eU����g9[�UYꫥ��֬�g�s�e�?  p�e�?��e�e5[f]Y֫UUU�lY�UUs�U   p�U �eUUe5WVsU�WUUU�\UUUUsUU�  pUU��UUUU5WU�U�WUUU�\UUUUsUUU  pUUU�UUUU5WU�U�\UUU5\UUUUsUUU  pUUU�UUUU5WU�U��_U�\UUUUsUUU  pUUU�UUUU5WU�U� pU5 \UUUUsUU�  pUU��UUUU5WU}U� pU5 \U�UUsUU   pUU �U�UU5\UUU� \U5 \UWUsUU�?  pUU�?�U5WU5\UUU5 \U5 \UWUsUUU� pUUU��U5WU5\UUU pU5 \UWU�UUUU �UUUU�U5\U5\UU� pU5 \U\U�UUUU �UUUU�UpU5\UU5  �W pUp� _UUU  _UUUW�U\U�   � ���? ����  �����  ���  �����������������������������?�������� �?��� ��?����<����3?�����������������?>�3;�����3/â��������������/??��?����<;3���� ��<��� ��?� ������3/�������� ��������?�?���<����3;�����<�����������?������.�������������ˏ ����/ �����������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ===============================  %&#  ===   ==============  $  = &#  ============  >>+   >)  ============  /(   >>(  =============  /*    !>'  ==============   -  =  )  ==============  ====  '  ====================  >>+  ====================  !>>*  ====================  >.  ===  ================   ,-  ====# =================   ===  >)  ===============   ==== >*  ================     ==  -  =============  !>>* =====================  >.  ======================   -   ==========)  ========= %&#  ========  (  =======  )  ======   '   ======  >'  ======  )   =====  >>$  ====  >'  ======  >>)  ==== >$  ======  />'  ===  >>%#   ====   ">)  ==  />)  =====   !>>'  ===  !>*  =======  /)  ==   >+  =========  /'  ===  >(  ====  ====   -   ===  >>*  ===    ====     ===  >>+   ==  #  ====  ==== = >>'   =  $  =========  >>>)  =  >>)  ========  >>*  = *  =======   >>.  == .  =======  >+  ====  ,-  =======  >>(  =======   =======  >(  =================  >*  ===============  >.  ===============  >>-  ================  >>  =================  >> =================== >>>==================== >>>>===================>>>>>>========================= =========================  ========================= /   ======================== !%#  =========================)  ========================*  ========================.  =========================(  =======   ==============='   ====  %# =============)  ==== )  ==========='   ==  >>(  ===========>)  ===  !>* ============>'  === >>+  ============>>)  =  ( =============>>*    * =============>>>.  =  . ==============>>+   ===  ,-  ==============>>(   =====  ================>(   =======================>*  ========================.  =========================-   =========================   ====================================================  ========================   =======================  >======================  >======================  >>======================   />=======================    ========================   "========================    @  PU TA  U PUUUPUUU     @ D  @QU TUU PUPUU  U Z�Z���Z��f�U�VU�VUj�VZ��fj��Uj�UZ�UYZ�YUUU�Z�U�ZZ��Zj�V�j���j�Z�     �  |�  p5  �  � ���\ee�|ee��ee� gf l�  p6  �  �     �   p  \  �  g6 �f� pff\�eWVe5W_}5�\�5?\? [9 �Y� ��  �   �  \5  \5  �6  �6  �6  \5  \5  \5  \5  \5  \5  p  p  �  �?  �  \5  W�  ��  ��  g�  �� �Ye�Ye��j�Z���f [�  ��  W�  �?  �  |=  W� ��V�eY�eY��Z�Z�p�fpYe�f�����j��UU _�  �  �  p  \5 ����eY�eY�����f�Z�p�f���pYep��pYe�W� �?  �?  �  p  p  \5  \5  \5  \5  \5  \5  �6  �6  �6  \5  \5  �  �?  W�  ��  [� ��f�Z���j�Ye�Ye ��  g�  ��  ��  W�  \5  �  �  _� �UU�j�����f�pYep�f�Z���Z�eY�eY��V W�  |=  �  �? �W�pYep��pYe���p�f�Z���f����eY�eY��� \5  p  � UUUUUTQUUUU�VUUUUQ�UYVUUQUUU����jUUUU������VET��������UU�����������UUUU� @p@\@�@�@=@=@=@@@@�>@�?@<@UUUUUUUU  @  @�@��C�:�Nq5\M�:�N�:�N�:�N�:�N�?�O��C  @  @UUUUUUUU�@�7@p@��@��@S�@S�@S�@S�@S�@S�@S�@\5@�@UUUUUUUU�@L5@�:@�:@L5@L5@L5@L5@L5@L5@�?@�@�;@<<@UUUUUUUU�@p@�@p@�@p@p@p@|=@|=@w�@w�@��@�@UUUUUUUU  @  @  @  @  @  @  @  @  @  @  @  @  @  @UUUU � p \ \ W�W����  � �< 0  0   �  � �� � �? � �0              � �� �5 � �0                         � h��                      0 �   00�� �  0�<������<3���0��<3 0���0�0�<3 �� ��< �0 00� 0  0��   0  ����l90��Ss4�\�5L14pt������������������������������������������������������������������������������������*��*��*��*��*��*��������������������       �       �       �       �       �<<     �<<     �0    ��     �0    �<<     �<8     �       �       �0     �0     �0    ��     ��    ��     ��     �       �       �       �������������������*��*��*��*��*��*��������������������    �        �         �         �         �?       ��6 ��  ����    �]�Z�?� �������? �UWuU�� ��������� �������������������갪�����������������:      � ��   \ ]�? _���W���_UUUUU� �WU���  �W��7   �_� �   ��     �W     ��  �?������������ ��?  �  �  �   �   � 0����� ��?  �?  ����������?��� �����?���?��         3  0�  �� ��������?������             ���* �VUU�`UUUU	�����
 Z�V�  �*��  �*��  ���� �ZUU��fUU�����V�UUUU�UUUU�eeYY��Z�V�UUUU�UUUU V�Z�  XUU%  �V�
   �*    `	    �    �    `
    �	    h&    �)    h&    �)    h&    �	    �         ���  hUU) �VUU�`UUUU	`U�ZU	`�*�j	��*�� ����  VUU� �YUUe����Z�UUUU��Z�V�%c�X�%`	X��Z�V�UUUU�UYeU V�Z�  XUU%  �UU
   ��    `	    �    �    `
    �	    h&    �)    h&    �)    h&    �	    �  UUUUUUUUUUUTUUUQUUUUUUUUUUUUUUUUEUUQDUUUUUUUUUUUUUUUUUQUPUTTUEUQQUUUUUUUTUUUUUUUUUUUUUUUUUUUDUUUUUDUPA@TAQUUUTAUUTQUUUUUUUTUUTUUUUUUPUTUUTAP@DQUU@UQ@UDUUUUUTUUUUUUUUU@PUTPPP  T @APTUUTUUUUUUUUUUUUUUUUUUUUUUUUAD ��
Db@D*E*��R"DFU$)�������@Q PE��PbAD ��
Db@D*E*��R U  "  UPD EQ��@Q PE��PbAD �������Ϊ������� ��� ���>����:���;���;���;���;���?���?�?��;�:��;�?��;���;����:���>���� ��� ��� ��� ���� � �?����� ������ �묿��� ;����� ;���? � ;����� ;��ï� ;� ��� ;�<����?��쯳��:���곪�?�?����        �        0       �       0        �       �#       2                        ?               
       �       �       	                �        /       
      �       �                       �                
        �        �                  4        �        �         �        �       �#        `                 ~        �        �        �       ��@P����������*(�*��������*��*(����������            �������������
           &         &�         "&         &           &  �
�*   &  �" "    &  "" "    &  " �
   &  " "    &  " �     &  �
 �*   &           &           &           &  ��*��
�  &     "&      &     � &  � �* &     "&     �  &           &           &           &  ��*��*�*&   " &   " &  � �
&   � &    &  � ��
&           &           &           &  ��
��*   &  "      &  "      &  �  ��
   &  �*     &         &    ��
   &           &           &           &         &�         "&         &           &������������&XUUUUUUUUUUU%������������*               � PA� Q�U T�PEh�P ��h��j�U@�UYP�YUPU�Z�U�ZQ��Z`�V�h���h�Z�      @� UP @�TU�UU��  ��T�UZ@YZ�YUUU�Z�U�ZZ��Zj�V�j���j�Z� X� PX�T�U T�@Eh�P��U@��`�U �UY �YU@U�Z�U�ZX��Zh�V�h���j�Z�  P   E AU  P  U @UUU PU � �UY �YUT�Z U�ZP��Zh�V�h���h�Z�  Z�  Z� @�U AU�  j�P��UU��P�U  TY �YUU�Z U�ZE��ZE�V�`���h�Z�  X�  Z� d�UVU�@Uj�@Z��Ej��Ej�U �UY  YU�Z  �Z �ZU�V�T���@�Z�   � PA� Q�U P�PE`�P ��h��j�U@�UY@�YU@U�ZT�Z �ZUV�P�� Z� �Z� �Z�`�U TU� Tj� X��Uh��Uh�UP�UY �YU   Z   ZU XU �PUU� UU Z�Z���Z��f�U�VU�QUj�PZ��Aj��Ej�U@�UY �  @   PU TU UPUU UU X�Z%��Z��f�U�VU�QUj�@Z��Aj�� �U@@YTPU  �Z A�Z��ZU�V�U��PZ�Z�Z���Z��f�U�VU�VUj�UZ��ej�� `�U �UY  YU�Z  �ZUZU� U� @    @   T  U   TfjTUUj UZ� Z� UU�
�U�
Z��j�Vj��%j�Z� @�B�FU�P VUBVZ
fj
UUj)TZ�U Z�Y UU��U�Z��@j�VEj��j�Z% U �A �P� VTVZPUfj  Uj@Z�YZ�YUUU�Z�U�ZZ��Zj�V�j���j�Z�  P    @P  @Q PUUdBUU @Z* YZ�YUUU�Z�U�ZZ��Zj�V�j���j�Z�Z�@���fT�VVU VZBfj
UUj)PZ�U Z�Y UU��U�Z��
j�Vj��%j�Z�Z���RD�fQ�VVU VZJfjJUUjUZ� Z�  UU�TZ%DUj)PUj�P j� 
 @���U�R VT VZPfj@UUj TZ�  Z� UUA�UEZ�Uj�@Uj�Pj�P Z� ���fA�VVUR VZ f
TU
 PZ
 Z	T UE�P @U
 PU@UU PU Z�Z���Z�f��VU%VUj	VZ�Afj�PUj)PZ* Z) U�UQZ�BUj�Uj�j� X�Z���Z��f�U�VU�VUj�VZ��fj��@jT �P �  U  PU AUUPUTUU  T Z�Z���Z�f��VU@VU* VZfjBUUjIPP� P�	 AU UA PUU TUPUU  U Z�Z���Z�f��VUVUj	VZ�Ifj�EUj�Z�UZ�YU��� Z P*@UUJTU T X�Z���Z��f�U�VU�TUj�PZ��Aj�� �U  PY  PUD@�Z @�ZU �ZU�TU�@U PUUPTT  U TP  @U @UTPTUU  @  @  TU@UUUU PU  @ VUYUUZV��jiY%��U	��V
(�Z�U��V��Z��(j��j* �j	��Z%������VU�ZUH�Z� �� �΋ ���� ��z�h`H�Z� ���� �s 08�s �0
�r ͮ "�
�r ͮ ��r �i�r ���r ��r �08��r ��r �~ )�0��s �����r ��z�h`ڭ� H�� H� ��� �L^��� �s 0"8�s �0 ��L^��r ͮ 0 ��L^� ��L^� ���h�� h�� �r ��ȭs ���`�Z����� �ǀ ��z�`�s  u�����s �r  u�����r �r  u�����r `�s  u�����s �r  u�����r �r  u�����r `����r Hȱ��s H�ȱ�H)�� h*�LУ�� ڬ� Z J��  �z�� ��� �Z�   J�������LQ����LQ����LQ� �����4�s � �L��s  ������ � �΋ L�� ΋ ��s ���b  �����4�s ��L��s  ������ ��΋ L�� ΋ ��s ���b  �����1�r � �^�r  ������ � �΋ L�� ΋ ��r ���b  �����0�r ��)�r  ������ ��΋ �� ΋ ��r ���b  ��z�� ��� �Z��r H��ȭs H���� H�m� �w  %�h�� h�s h�r  ���� � �L
�z�� ��� �Z�   J������������������b  �܀ܭ� H �����#h�� z�� ��� h�s h�r ��r ��ȭs ���Fh�� z�� ��� ���)͋ ����)��hh�#hh��r ��s ��� �7�� ��y �$ ��L�� �� �L���r H�s H�r � 058� �r �
*r r �s � 08� �s �
s s s s �. .�h�s h�r `H�Z�r �0�0�� �8�� �� �s �0�0�� �8�� �� �r 8� � �s 8� � � z�h`��ꍠ ��ꍡ � ���� ȱ��r ȱ��s ȱ��)�� ȱ�)�� `� ��ꍠ ��ꍡ � ��� �ȱ��͍ ���͎ � K��F��ѭ   J������ �ϩ 9� �é l� �� 0Ţ" mɩ �r �]�s ��� �#�� � ��`�#�r �D�s � �� '� �Щ�r ���s ���)�� J Щ �r �\�s ��� �#�� � �ʭ   J������L�� �� ѩ�r ��s ��� �7�� ��y �$ mɩ�r ��V�s �c�o  ^Ю   J�����
 9ѩa�o  ^Ј��$�� ����
 9ѩa�o  ^����
������h�V�s �c�o  ^��� �����Ф �� ����m� �w Lڡ�� ̧�-�� � D��!��L٥ Q� � �� *� �� �� �ϩ
 ѩ l� �� 0Ţ" m�`�r  u�����r �s  u�����s �s  u�����s `�r  u�����r �s  u�����s �s  u�����s `H�Z�u JJ:�� �t �� �#�r ��s  '� �Т#�r �.�s ��  '� �� '� פ �� ��z�h`�  ���� � ����**����� g�`H�Z��r ��s � Щ�r �(�s � �� '� �Щ�r �<�s ���) '� �Щ�r �<�s � Щ�r �L�s �	 Р��)���r �n�s  �ȭ   J��� ���� �ϩ �z�h`�Z���**�Lg��� ڬ� Z�y ����r Hȱ��s H J�� �m� �w  %�h�s h�r  ��z�� ��� �Z ^Ţ ��  (��   J����Lb����� � (�ʀ0 (��� �(���� � (�� (�� ����������з� �ώ�  (��
 9р� ��� � �� ���v�v  j� ȩ�
 9ѭ   J�������L@����L@����L��v J8������y 
���b  �܀ǭ   J����� � ��  ȩ�H���� �	��  ȩ�5z�� ��� L٧���� � ��  j�����L��� �	�L���  j��y L�� �ϩ l� ��z�� ��� ���)?��� 9р ��z�z�`HZ�� H�� H� �� � �� � �0� �� � �m� �w  %ĭ 

�r � 



�s �v  ��h�� h�� zh`HZ�� H�� H� �� � �� � ��0� �� � �m� �w  %ĭ 

�r � 



�s �v  ��h�� h�� zh`Hڭ� 

�r ���s ���� ���  ��h`  �  �U U   �S? ��     �  p1  p� T L? \�  �        �����?WUUUU5����4����4�3���4�����4����4����4WUUUU5�����?  W5    W5    W5    W5    W5    W5    W5    W5    W5    W5    W5    \    p    �    ��    �WU�    \U   �W�V   pU5  �_U��@�   pU� �UUU��_  �UU�UUUUUUU�  �UUUUUUUUUUUU �UUUUUUUUUUUU= �UUUUUUU  VUU �UUUUU����ZU�  ���WU���j�X�  p��UU]UUտ�?   𪶪�WUU��    �j���UUU      �� �UU�       �?  pUU=           \U�           ��?                                          ���           �UU�           �UU���         _�ժ�   ��?  �_U}U��   pU� �UUM R]  �UU�UUU��W�  �UU]UUUU��UU �UUUUUUUUUUUU=  WUUUUUUUUUUU  WUUUUU TUU�  ���UU���_]U�  p�zUU����s�?   𪦪�WUU��?    �j���WUU�?     �� �UU�       �?  pUU=           \U�           ���              @D                      W           @UUU                     �Z           TUUUU                     ��           UUUUU                    ��          TUUUUU                   ��          TUUUU                    p�         TDD                         p�                   U                 p5                  UU            ���� �5  U             EU          ��������: PUU                       ����������: TUUU                       ���������UPUEQ                        �������U                             ��������U                            ��������U                           ������������>                         ���������ꮾ���                         �����뻾�������                         ��������������     UUUUUUUUUUUUUUUUUUU���������������WUUUUUUUUUUUUUUUUUUUUUUU���������������_UUUUUUUUUUUUUUUUAUAPUU���몪����������^UTAAP@DUAUEUQEUTQժ��������������^TQEUUUUUTUUUUEE�����������������EUQTUUUUUUUUUUEUUEUUQ�����������������TEEUTUUUUATUUUUE@TU�����ﯾ����������E@TDU ETTE QQUUUUUU뿪������������UUUUUUUUUUUUUUUUAUEP��������﫾��������WUQUUUUATUUUAUUEUU�������������������WUEUUUUUUUUUUUUUDT�������������ﯮ���GUDPQ@UDQ UUUTU��������������������WUUUQUUDEUUAU UP@��������������������CTUUUUUUUUUATEUUQU�������������������UUTUEUUUUUUUTUUEUUQ�����������������WUTUEUDQQUUEEUUEEPDQ����������������UDADDUQUUUUEUUUTDTU����������������WEEUDPUUAUUEUUEAUUUUUUU��������UUQUAQTUUPQQTUAUQTTUDU�UU��������_UPEEQT@UUTUUUQUEUAUEPU���WUUU������WUUUUQUEUUUUUUUUEUUUUAQ��UUEUUUUUUUUUTUUUUUET@@QUETDUET@@QE QDUUETATQPUETATUUUETATQPUDD@UEUU@ TU  UU@ @UUU@PTU@QUD EUQTUEQUTUQTUUUEAUQTUEQUTEUQPUUUQPTUEAEUUQPQ@UUTUUQPTUEAPUQQUT@EUQ QUT@ETUPQUT@EUQ UEU @DDTUEQUDDTUEUUQ@DTEQDDUPAP  A @AP  P@  AP  A   @QPUEUUTUTQUEUUTUQAUEUUTUTQUTEPET @UQ U AUE PU @UQ  UEQ T @UU @UU QTUU @UU EUU @UU QTU DQDUPATUADUPADQTDUPATUAQATQUUUUTUUUUPUUUUTUUUUUUUUTUUUUPUUUUAUTUUUPUUUUTUUUUUUUUTUUUPUUUU@UUUU  PT @  P@ T PT @P U@@ TU@P QUATU@P U@TU@P QUADUPU@UTUP@UTPUAU@UTUPTUP@EUTPUUPPAUTPUATUTPUUPPAUUAAU @U@UUUUUUUEU@UUUQPUUUU@UUUUUUUUTUU  @UU   UUP @UU  PU  @UU   UU  TU PUETTQUET AUUETTQA@PUD@@@ @   P@ @  @@ @     P EA U T TP U T A  U T TP@P EQU  TA  PU  TA  U  TA  PP @UQPUQAUAUEUPUQAUTUTPUPUQAUAUEUUTDUTUTUQUPUTUTUUUUUTUTUQUPUEUU@U UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUAUUUUUUUUUUUUUUUUUUUUTU    �?      ��     �YU    |]�U   �_UU�   �UUVU5   |U�WU�  �W�uUU�  �UYU�W� �_VUUU?  |eUUuU�  \YuU�U� �WUuW��� ��_U^U�� p�\uzU�  p\}�U�  �W]��� ��U]?�W ���]�� ������   �����5   �??��   �< ��   �0  �  � 0  �    �  |       p5       �5       ��        �        W       W       \       �       �       \       \       \       \       l       �       �       �       W       W                                  @      P       P U      P             @@     P @     PP     PP     @T     PT     PT     PP     TP     T@U     TE T     DU@         PET    @TT   P PT   @  @Q%   @  A�      �             	   P @Q	   @b  E    � U	     YP	     `P     �*      U�      �U�      `��      ���      @�     ? �    �� Z
    ��p    �]�	    �U5�    �U5     �U5 (    �U5 ,    �U50    �W�0   �UW�    _U_U?   WU]U�    \UuUU#   ��UU     \UU�     pUU}�    �UUu�     WUU�     \UU�     |UU�    ��U[�    �����           @            @      @@            AE      PP      P     @P     PP     P     PP     PP     TD     T@     TP     TU     TU     TUT     PU@    PT     PQEU    �QUT    EUT    HAQ�     EA�     @U   P PU     PT	   `@@Q	   �  E   � E    VU@    �@P     V	      U%     @�U�      `Z�      ��        �     ? �    �� Z    ���
    �]�	    �U5�	    �U5 +    �U5 &    �U5 ,    �U5     �W�    �UW�    _U_U?    WU]U�    \UuUU   ��UU     \UU�     pUU}�    �UUu�     WUU�     \UU�     |UU�    ��U[�    �����          �����
 ���������j�ZU���
�V� �Z�
�T PP*�     @*h     @)h���<@)h���?<@)`��<<@	h���<<@)h����<@)Z���<@�Z�<�<�C�Z�<�<��Z       �Z     P�hUP @U)�V�UUUV�*�j�ZU�Z�*�������� �*����*  �
��*�                                                                                                                                                                                                                                                                                                   ���ة��  ��� � �� � � �� � �ύ& ��" � t ����k ��l �� � �k����l ��� �XL �H�Z�~ � � �� (z�h@H�Z�' )��h ��� �� ���~ ��# �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                                                                               W© Qќ� �(��  é��  �� d©x��# � Q�L � �ϩ Q� � �© �^  �ܩ l� �� z� �� �휨 �� �� �� `�� �� �� �� ��� ��� �� �(�� � �b�� �����$��  ��`�  ���� � � ,�`� �w � ��ꍠ ��ꍡ �ڮw �A둠������w �� ��`ک'�r �^�s �	�� �$�� � ��`� ���� � � Xâ��� Q�L}�`H�Z�k �@�l � � � �k����l ���z�h`��^  �� � T� �ϩ
 9ќ�  � �֜� �� �� Lx�`��^  �� � U� �ϩ 9ќ� � �� ������ Q�L�� �  �� �`H�Z�� � �[�  ���� J�	����
� ��� �  	����
� � �� �  	����
� � �� �  ��$��� 	����
� ��� �	�w ���b  �� %ĭ  �����L�� �ϩ
 9�z�h`H�Z Ѯ �� �s  f�� �s i�s ɐ0� f� y�z�h`�Z�  �����	�����0�z�`ک�� ��� �  ���`H�Z��t �<�u  0Ţ" m� ⦭  ���� J�	�����u �� 0� ��8��u �R�  	�����u �x� 0� ��i�u �4�  	�����t � � 0� ���t ��  	���Ж�t ��� 0� ���t  0Ţ" mɩ 9ѩ��h ��\  i� � ��L��z�h`�t �r �u �s ��� ��� �y `H�Z�  ���� L	�z�h`H�Z���JJJJ
��덢 �덣 � � H

�r ���s ���v�� ���hi����� �h�� θ z�h`H�Z �ŭ� � ��� ��� �ϩ
 9� ��LR�z�h`�  ������ �����`� m � � m � � ���� � ��r � ��s � ��� ����$��� 0ѩ��  9� �� 0Ҁ Ǹ �̀ �`�� � � �� �ҩ lѩ 9�`H�Z� 8�� �&J��� ���	�� � ���	8��鍈 ��z�h`ڜw � ����� ȱ���  ���� � ��r ͙ ��s ͚ ��w �� 0ݭw �0���� �`�Z���)�0 �ƀ V�z�`�� 
���덶 轹덷 �s 
����� ȱ��� �r ���=�� �>����8�6��2� ��ꍠ ��ꍡ � ��� �����r �ȱ��s �
�� 0ԩ ���`�� 
���덶 轹덷 �s 
����� ȱ��� �r ���>�C� ��ꍠ ��ꍡ � ��� �"����r �ȱ��s �ȱ�)������
�� 0é ���`�� 
���덶 轹덷 �s 
����� ȱ��� �r ���>�2� ��ꍠ ��ꍡ � ��� �����r �ȱ��s �
�� 0ԩ ���`�x )�JJJJ�y �x )�x �
08�
�x i�x ��y � ��x i�x �y ��حx `H�Z�� 
���덶 轹덷 �r �� 
����k ȱ��l � � ��k i�k �l i �l ��� �k
� ���r �r �r �r ��
0�z�h`H��� ��� ����4 Qʢ8 .ʀ���2 Qʢ6 .ʀ� �ʀ�h`H�Z�x  �ʢ � ��- ���̃ ��
 9� U��� ��z�h`�x ��썄 ڮz  1� ������h ��\  i��x m� �x �r m� �r ��� 9� ����y п`H�Z�x  �ʩ�q my �q � �p � � ���p���y � ���1�������̃ �� U��p i0�p �q i �q �� ��z�h`H�Z�  �ʩ�q my �q � �p � � �p���̃ �� U��p i0�p �q i �q �� ��z�h`H�Z tʢ � ��Q����̃ �� U��� ��z�h`H�Z tʢ � ������̃ �� U��� ��z�h`H�Z tʢ � ��1����̃ �� U��� ��z�h`�Xꍞ �X�m� �� �x  ��`��鍞 ��鍟 m� ��  ��`�� mx �� �� i �� �@�� � �� �s � ��� i0�� �� i �� �� ���r m� �� �� i �� `H�� �� �x  1�h`H� �  �ʩ�� h`H�Z�� �� �x   ˀ��ꍞ 轠ꍟ  ��`H�Z �ʢ � ��- ���̄ �� U��� ��z�h`�� i0�� �� i �� �� m� �� �� i �� `H�Z�  ��譈 � �Q�r � 0I8� �r �
>r r �s � 008� �s �
%s s s s ڮ� ��	�� �Ȁ�� �����w Пz�h`HZ ̩�z �	�y �; -̢; -̢� -��y �� ��z ��zh`ک(�r �f�s ��� ��� �n ���`꩐�� �X�� �w �x �/��)





�w ��JJx ���w �x �����8�� �0�� �� � �� �����`��r �2�s �  Щ�r �F�s � Щ�r � �V�s �c�o  ^Э   J����� �,�5���� �"�+������ ��� �: â�� �֩ Q�L��a�o  ^�Ȁ	�a�o  ^Ј�V�s �c�o  ^Щ
 9р� �� ѩ Q�L}��g�s ��r ��� �
�� � �� �ͭ� �&� 0Ҁ	 �� G� ��`�I�s �&�r ��� ��� �l �� �� �ͭ� �* �� G� �р 0�`H�Z�&�r �W�s �
�� ��� � �� � �� �ͭ� �,0�� 9� 0Ҁ�&�� :π t� G� ��z�h`H�Z� 9Ѭ� ���� �,0�.�L�Ω��b  �ܜb � 9�L���(�}�*�=� � ���h ��\  i۹��r ȹ��s ȩ�� ���  ʩ 9� ����0�L�΢@����h ��\  i۹��r ȹ��s ȩ�� ���  ʩ 9� ����H�׀v�����r ȹ��s ȩ	�� ���  ʩ��h ��\  i۩ 9� ����0ʀ:�����h ��\  i۹��r ȹ��s ȩ�� ���  ʩ 9� ����0ש 9�z�h`��r �F�s ���� ���  ����  �ө��h � �\  i۩ 9� � _�`��r �S�s ��� ��� � ʩ��  �ө��h � �\  i۩ 9� � _�`��r �\�s ��� ��� � ʩ��  �ө��h � �\  i۩ 9� � _�`��r �f�s ��� ��� � ʩ��  �ө��h � �\  i۩ 9� � _�`H�  ���� �h`H�~ �  ����~ �0�h`��� � Q� �֩ Q�L�H�Z
����| 轲�} � �|�$�#H�x ��� h�a��b�8�7�o  ^��r �r Ȁ�z�h`H�Z�o �a��$L���b��%L���c��&L���d��'����k ��l ��w �s � �m �@�n �m i0�m �n i �n ���r �k- �m�k Ȳk- �m�k �s �w п8�s ��s z�h`� �  ^Щ�� `H�Z�)�JJJJ�o  ^��r �r �)�o  ^��r �r z�h`ڢ '�����`H�Z���������z�h`ڪ ѭ  �������� ���`Hڪ���




�y ��)y �& �h`H�Z Q�
���獞 轧獟 � �� �@�� � � ��- ����(���� i0�� �� i �� �� i(�� �� i �� ���˩ύ& z�h� �� Q�L%�`H�Z���b  �ܜb ��y ��w �d�s �
�r ��� ��� �  m� ��s �w �� mҩ 9Ѣ  mҩ 9��y ��z�h`H�Z���b  �ܜb ��w �d�s ��r �	�� ��� � mҩ 9��s �w ��z�h`H�Z��鍞 ��鍟 �@�� � �� �s � ��� i0�� �� i �� �� ���r m� �� �� i �� � � �� �S��- ���̃ �� U��� ��z�h`H�Z��w � �� �@�� �  �� ��w ��z�h`� ��I�����(���� i0�� �� i �� ����`H�Z��� ��r �Z�s �� )�o  ^��r �r ��  �Э�  �� X�z�h`��� ��r �#�s �� )�o  ^��r �r ��  �Э�  ��`H�Z��r �
�s � Щ�r ��s � Щ�r �7�s � Щ�r �B�s � � �� "�z�h`�� � � ��Ϋ �� ��`��� iP�� �� i �� �� i )�� �`H�Z�� ͪ 0&��� ͩ 0��� ͨ 0�� �� �� �� �� �� z�h`��r ���s ��� �	�� �x �ʩd 9� é�r �2�s � Щ�r �F�s � Щ�r � �V�s �c�o  ^Э  ���� �!�*���� �� ������� �2 �� �LQթa�o  ^�Ȁ	�a�o  ^Ј�V�s �c�o  ^Щ
 9р� �� ѩ Q�L}�� �N鍠 �N鍡 � �P鍶 �P鍷 � ��Ѡ����	����0߀�J�� 
i(�� ���r �x�s � Щ( 9� Ü� L.¢��L}���r �(�s � Т �I�r �F�s � Т  � �ϽI�r  �� � � ^� � ѭ  ������� �� 3� �Հ���� �� ^� �Հ������ ��L�Ԁ'��� ��� ���� ���� ������  �Lx��Z� �N鍶 ȹN鍷 ���o i7��z �`H�Z� �N鍶 ȹN鍷 �����b�8�7�o z�h`H�Z8�7�y �o �a�
�y �o ��A8�7�o ��a�o h`H�A8�7�y �o �a�
�y ��o ��Z8�7�o ��a�o h`H�Z�	�w �  ��譈 � ��s �s s s �r  h��w ��z�h`� � � �  a� eۜ � � � � � � � �* �[ �d � ���\ �h `H�Z� ���%�? � aۭ8 � �9 �  ���? �? �: � 4ح ���%�L � eۭE � �F �  ���L �L �G � �ح ���X� ����# � aۭ � � �  �٭ ����1 � eۭ* � �+ �  2��# �# � � ���1 �1 �, � � i� ��z�h`� �� ȱ� ȱ� ȱ� ȱ�  )
��o�! �o�" �  )0�& ȱ����\ �h Ȍ �# �$ � � �L�ج%  ��� �� � ��% ��Ȍ% � ���5 �6�8 ȱ6�9 ȱ6�: ȱ6�; ȱ6�< )
��o�= �o�> �< )0�A ȱ6����\ �h Ȍ5 �? �@ �: � �� � � �b )����� �B  ��`�B �C�E ȱC�F ȱC�G ȱC�H ȱC�I )
��o�J �o�K �I )0�N ȱC����\ �h ȌB �L �M �G � Ш� � � �b )��@З��� �5  4؀��' �(�* ȱ(�+ ȱ(�, ȱ(�- ȱ(�. )
��o�/ �o�0 �. )0�4 ȱ(����\ �h Ȍ' �1 �2 �, � Ч�3  ��� ��( � ��3 ��Ȍ3 �' ���^ 
��7�` �7�a �`� ȱ`� `�^ 
��?�` �?�a �`�( ȱ`�) `H�Z� )?	@�O � I��-O �O �$ �!��  )@��J��O �O �& �8��& ��  )0�& Ȍ$ �!����$ �  �$ �O � z�h`H�Z�- )?	@�O �- I��-O �O �2 �/��. )@��J��O �O �4 �8��4 ��. )0�4 Ȍ2 �/����2 �. �2 �O � z�h`H�Z�; )?	@�O �; I��-O �O �@ �=��< )@��J��O �O �A �8��A ��< )0�A Ȍ@ �=����@ �< �@ �O � z�h`H�Z�H )?	@�O �H I��-O �O �M �J��I )@��J��O �O �N �8��N ��I )0�N ȌM �J����M �I �M �O � z�h`� `� `H�Z�\ ���%�] ���\ �d �] )?
����f 轧�g �e  ��z�h`�d �* �[ `�e �f�W ȱf�Q ȱf�R ȱf�X )
��o�T �o�U �X )0�Y Ȍe �S �V �W � �ۜh `H�Z�d ���L�ܭQ �Z �W I�Z )��Z �V �T��X )@��J��Z �Z �Y �8��Y ��X )0�Y ȌV �T����V �X �V �W )�O �] )����
�@����O �O �Z �( �O �[ ��* �[ �S �S �R � ��z�h`H�Z�  �٠  �ٜ �' ��% �3  �� � �� 2� i۩�� z�h`H�Z� � �
� � ��c �b )?�c �Q�� �K�c 
����6 ���C 轇�7 ���D �5 �B � � � �b )�����  �حb ���  4� i�z�h` ��� �(�� �(�� ɠ�� ɠ�� �(�� �(�� �(�� �(�� �(�� �(��(�� �(���� �(��(��.��.(��(��@(���������� d(�� Y(�� d(�� q(�� w(�� �(�� �(�� w(�� d�� P��     � �(�� �(�� �(��P��@(��.(��(��@(���(��.(�� �(��(�� �(�� �(��(��.(��@(��.(��ȧ�(�� �(��(�� ���� ���� �P�� �P�� �P��(��@P��.(��(��@(��     ��(�� P��(�� �(�� �(�� �(�� �(�� �(��(�� �(��(��.���.���     ��x�	�(���x��(���x��(���x��(���x��(���x��(���x��(���x�	�(���x��(���x��(���x��(���x��(��Rx��(��Rx��(��Rx��(��Rx��(��     � �(�� ��� ���  � ��� ��� ��� �(�� ��� ��� �� ��� ��� ���(�� ����� ���� ��� ���(�� ��� �(�� ��� ��� ��� �P�� P�� _P�� T�� _�� ��� ��� ��� �(��     ���	���������!����!������������������	���!�����!����������     � �(��Tx�� �(��Tx�� �(�� ��� ��� �(�� �x�� ��� �� ��� ����� ��� ��� ����� ��� ��� ��� �(��Tx��     � (�� (�� �x�� �(�� �(��Tx�� ?(�� ?(�� Tx�� (�� (�� �x��     ��(�	�(���(��(��!(��(��!(�	�(���(��(���(��(���(�	�(��!(��(��!(��(���(��(��     � q<�� j<�� q��� �<�� <�� �<�� �<�� ��� ��� ��� �<�� ��� ��� j��� _<�� j<�� q�� �� qx�� ��� q�� �x�� �<�� �<�� ���     � �<�� <�� ���� �<�� ��� ��� �<�� �x�� �x�� ���� �<�� ���� q<�� ��� �x�� �x�� �x�� �x�� �x�� �x�� ���     � ��� _���     �     � �
�� /d��     � /n��     � ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �(��     � ���     � d�� �� ��� ��� ��� ���.��T��������\�����!��     ���� ��� ��� T�� 2�� �� (��     �!��\��     � �� � _� � �� � G� � 8� � /� � %� � � � ��� ��� ��     � 0# 1#� 3#� 4#� 5#� 6#� 8#�     � �
	�
�
	�
�
��



		�

		�
	�			�
�G�S�[�g�O�W�c�k�?����  �  ��  ��  A�A���  �  ��  9�  U�X�w����������2�����;���������%������G������%�����������-�@�G�V����� ��    p/   �O�   �   G G G G  &� &   w &� &W J   ����   �O�   ������   G G G G G G G G    o<   /�    � � �������)�4�?�J�W�_�s�y����������� ������������� �'�.�5�?�CONTINUEa$END$aaaaaaaaaa$aFIGHTERaa$SUBMARINEa$DESTROYERa$BATTLESHIP$FLAGSHIPaa$CURRENTaLIFE$ALLOWED$SEARCHINGaTHEaENEMY$MOVES$bPASSWORDb$HIGH$YOUR$PASSWORD$aaINPUTaPASSWORD$SCORE$PASSWORD$aaPASSWORDaWRONG$NEW$PROGRAMaBY$ZHANGbXIAObMING$GRAPHaBY$ZHANGbLI$MUSICaBY$XIAObLIbWEI$TRAVE$WORLD$HEART$STAGEd$SCOREd$TURNSd$CbNUMBERd$PbNUMBERd$
� ���2F%/9"1<
P bd�x
1<!P
b#d�x
7B#Fnd��"
1
<P!bd �x	 xg]Snnnnyso xtni���:�ֈ�V���։�V���֊�V���֋4���t� �$�H��\����܌�S���Ӛ�S���ӛ�S���Ӝ�S���ӝ�S���Ӟ�S���ӟ^j�j�c�d.u�vʐF�j��w��~z�S���������c���c�,�>�b����������e�ef3f�f�g.kQ�\�~z"�b���V�      ���������4���I�e���ƻ�usnkb
[	G<0# %*/49>CHMRW\afkp(�-�2�7�<�&*,.v&(*vv(,.vv*.vvv&(*vvZ�<�2*�2*�28�28�(F�(F�(F�Z < < <222 2(
(((((	(���=�y�a7 � � ��:�W�t�����ˀ��"�?�\�y����:�W�t�������Ё� � � � � � � �
�'�D�a�~�����Ղ��,�I�f�������ڃ���1�N�k�����߄���6�S�p� � �����ǅ���;�X�u�����̆��#�@�]�z����� � � � � � � � � � � � � � � � � � � � � � � � � �ч��(�E�b������(  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  ������������������������������������������������������������������� � �� 9ѩ(�r �r ��s ��� ��� � ˩ 9ѭr �B0ݩ�� ��� � ˩�� ���  ���w �
�y ��r �
�s ��� ��� �y  ˩ 9�8��y ��w �� í� �r �� �s �s ��� ��� � � ���r ��s ��� �� �x ��� �r 1˩ 9��r 8�(�r � ����� �ۜw  ��w �w �(�  ��`����` � ���y �A�{  ��L�� �� 9�8��y �y �  ��`����`��r �/�s �	�� �@�� �y  �`�� �Z �s �� �r ��� ��� � � � ���`�\�s �r �(�� �D�� �, .ʩ�r �/�s �	�� �-�� � �`� �z ��w �r �{ �� �{ ��L{�	�� ��� 8�A� �s � ˭w � � c�� B�ͭ� �{ � ���w  X�`�A8� � ��`�� �z 0Ί ��{ N{ N{ �{ �{ �{ �w  X�`�� �	��������`H� �� ��^  �ܜ� ��r �(�s �
 Т����� s� �� ���r �� �s �� �� � � G��� ���+�r �i�s � ��� ����� 4ڀ�� ��  '� �Щ+�r �r�s ��  '� �Щ$�y �( -��y ��L�� �©��y �( -��y ���
 9� é
�r ��s � Щ�r �� )�o  ^Щ
�r �2�s �  Щ�r �� )�o  ^��r �r ��  �Э�  �Щ
�r �P�s �! Щ�r ��  '� �Щ
�r �n�s �" Э�  '� �Щ
�r ���s �# � ��r ���s �� )�o  ^Щ� 9ѩ� 9ѩ �^  ���h`�� �  ���� � �� ����`� ��ꍠ ��ꍡ ����� ȱ��� `H�Z��w �  ���� � �< ���	5���h �
�\  i��w �*� 8���0����� �����h � �\  i� ������z�h`ڭr ͔ 8�� �r �� �8� �� �s ͕ �� 8�s �� �8� �� m� �`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �<?�<<<<���������?�< < �?  �?�< <�� <<� �0�?  �? �< < <<��< �<<��?<< �����<<�<0<��<<<�? <<��<<�?<<<  �<<�<<�  �<   <�  �<<<<<�  �?  �  �?  �?  �     �< ?<<�?  <<<�?<<<  �������  �?    �  �� ? � �        �?  <??�?�<<<<  <?<�<�?�??<  �<<<<<�  �<<�     �<<<?<�?  �<<�<<  �< � <<�  �?������  <<<<<<�  <<<<<<<<<<0�  <�<�<�<�<�<<  <<<0�0<<?<  <<<<�����  �?< �� <�?                        �?�?      � �
�	**�	�
�     ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            O� �e�