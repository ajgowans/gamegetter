�5
����-���.l- ��=�}�������Ӄ_�()*./0+,-������������ԩ ���� !����#��+�0�����Y��[� 	� �憥���� *� �� o� ���5`� � �������F !����)�<8�
����'���(�}����~���� ������+� �'�-���. 5�� �)�! È 	� �� �)� �
�ͦ<ʼ寥 8�
�����)�+Ȅ,� 8�

e,����-���.е�5 ��`�;�@���L����@���� ���`�0�0� �<�  �����e<�� ��੅�:��0��@�� �F�� �L��@�S����X���� �`���� �#��p���e<
��^��-�_��.���0�-�  �������`��)������0 k�` ����`�`�
�ݩ �`�0���K�O k��5�<�@�� ��` �� *� ۍ M� �� `� �� � ^� (�`�F�}�G�F���G��o� �G� ��F�F��� �F�;8��;0���; �� !��̅+�8�)�i�-�?8�)�i�. 5�� �!���! Y�����-���.�� È 	� �`��)�E����;�:��5��6� ���@�;�:�%��<�	������ �J�=�
������4`��4`��_���`��)�/�;�,�@�;���
��� ��`�5� �s�� ��`��5 ��� �s`���; ��� ��!������" щ ��`     �E
��p��-�q��.l- z�����z����Y�� �� �J������(���� �  ���E`��)��J 6��J���E`�0�` =���5� �E�<�@�� ��`�#��6 ��<�<��� �<�̓�������4��`��4`                                                                            2(��0�D�Z�m����]��� �� ��` ���0����� k��_I�_ ׅ � l� �� 1�`� ���M�N�)�:� ��4� )��� )� � )��� )� � ���% ���)E � �
� ��� ��`����悥 J�3J�ZJ�L����)����`�)��έ?��� ݈� ��� ��`��)����`�?)�Ф�ɒ�� � � ��`��)����`�?)����� 	�� �� ��`L􄭟)��4��`�)���?�z�� �� �٩4 ��`��� ��;���; ��`   Ȇ� �2�-H�.H 1���0h�.h�- 5�� �!���A���� �� � ���`ɐ���!)�� �P�!�+�i�ÆH !� È 	� �h�' r���`)�ɀ�̱!ɀ���Ɂ��5�5�s� � � ��)�� ���!�+ !� È 	� ����� h����
�6��@���� ���`�0�0� �<� �5��慩�5���� � � `
� � ��)���)��)�?� �'�)��2��)��?)�#���?)����}υ�-�?}Ӆ�.� `��%�ƅ&`� �"�:8��!�
��
�!�"�� !����Y��"i�+ 	� ��Y����!i�+ 	� �`� �"�<�!�
��
�!�"�� !��̅�[��"i�+ 	� ��΅�[��!i�+ 	� �` !�� ������Y���i����Z����<i�+ 	� �Ɔ�����`������������� ���;�� !����燅�+�[�������� 	� �憥����`�����+�� 	� ����燅�[����� �©��C��-��. �����燅�[����� �¦�����C��-��. ��� ��� �C���-���.� �  ��` 5�� � �!���0���!��� `�@��-JJ����.�� ���`�0� i�-� 8��. ��`�0� i�.� i
�- ��`�0� i�.� 8��- ��`�0� i�-� i
�. ��`� �!��"�-8�JJJe!�!��"�.8�JJJ���!i�!��"���`���'���'� ��!�����'�
��
�'�$��'�# щ ��`	 	 	    	� �!u=�=�
��
�=�>����q�Bٳ����Aٕ���q�: *�`� �D�;�����D�D��)�������`���5� �E� � �� ��`�F��)0��;���F� �G`� ������`          � ��P������)�� �d��X�����`�5`�0����	�@I�@`�@I�@`�0� �M�N��J�,J�OJ�r� ��
���� ��`� )�� ݈� ����N`� ɒ�
���� ��`� )�� � ���M`� ��
����4 ��`� )�� 	�� ����M`� �z�
���� ��`� )�� �� ���N`�eM��?eN�?`�0� )�� y���� i�`              � �L��0�@0&�`�`�`��� �`�P�����
�0��L ���0�0��ͥL�	 � 1� ��` /��0����� k��0�@I�@� eM� � eN�  �� ��`� �M�N�0� )����)���M`����� )����)���N`�����p� ����J�&J�DJ�c r��0� �z�p��憽�/�k�i ��Le� ���0� ��pН憽��� ��LG�LU� ���0� ���p��憽������ ��LL� ���0� ��p��憽�/� ��L`� ������ ��� �� ��` ��� ���� ��� ���� ��� ���ۦ0�����p����Le���I<��` ����/� r�� ��Ш ��� ��4Н ��� �	�� r�� ��0�����p����LL�LG���I��`�0� )��)� )�� � i�-� i�. 5�� �0�!����0`��0�P�"i�Pɀ�)� �P�� ����� k�L�� �i��� � �0�iɴ�� �0�0�0���`��0��H�@���	�0�0���` ʏ�-e.�������� �� � ���`�����0H��0 k�h�0�0��к�� k�L@���H�@����P� ���H�H���`4��0�@0�0�0���`�H�� ʏ�-e.����� �0� ���P�H� �ש�P`�0�H��=�)�KJ�J�)J�4�4� � � �� ��`� ��`�� � � ���� � � �ڐީ� � � �̰� P��H��)J������`����5�
�_� ���`� � � �� ݈`� � � ɒ� �`� � � �� 	�`� � � �z� �`����)� � 



e ��U��p`� �-�.�0�H��8������@������������-�-�-�8������������������.�.�.`� �-�.`��)�e� �P�Z���T���-i�����.i����@0��8�������8��
�%���!�� �ڊH 5�� ��!�+ !� È 	� �h��P����`� ����� ��`�����Ȑ� ���H��i����i����0�@���
�0�0� ��.��8�������8��
����ڽ���ө�� k�Lϐh�H���-���. 5�� � �!�+ !� È 	� �h�L��12345`�Y��J�

i��/��+ !���!�" 	��!�܅#�"�$�-�+��)��*��&� �/�%�(�� %&�' ��'/�/�%�%��� �%�/� �© �/�#�� %&�' �L���#�''L��&&�!�#�(�(�������+�
��&� �(�)��*� ���$��8�-���L_��.�LU�`�(8�%��	0F'F'���`''���`��0�@0����� k��0�0���`
 #(-4<>IKQ_din�O�K�:����)� ��P �֤<��


e �� ��-��. 5�� �!�j�-i���.i����@0��8�������8��
�=���9�� �ڦ �P�-���.���h)�� i��!� �X�i iͅ+ È !� 	� ��O�h`���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5
����-���.l- �D�u�������ץJ�

i��I����+ I��J�J��� �J�5`�J

i��O��8�J��
i�+ I��J�J��ک �J���5`�0��
���4��6`�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5
����-���.l- )�f�𘸙()*./0�������ԩ ���� !������+�!�����Y��[� 	� �憥���� *� �� ���5`�@���G��0�J��V�?��_������� � ����@���� ���`�0�0� �<�  ��`��)������0 k�` ����`�`��ݩ �s�`�0�� k��� ���5` �� t�`��0������ �� ��` ������ k��_I�_ 8� l� ��`
 Ȇ� �4 5�� �!�+)�ɐ�%�!)��3�H� �!�+ !� È 	� �h�' r���`��-�� ��;� ��` ���5� ��� � ���`�0��@����0� �<� ���`�����4��6�@�;�`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5
����-���.l- �>���@� �����0�H� �e� ��� ���5��6`e}�)��>&������6��4�t�:� �=�>�?�@�A�B�q �` ������I����<�� ���)���ߩ �0 k���6`�����6`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������DTl\l|�4\\4,�lD\�ld$,\,|$,TTlD|\�dD<<T�<4��L$$|Tl4T$D\\|T|<4�\$$l4<4|d4|,�\l\T4�T4t�,TdD$��Ld<�tLTt4\4T4|t4dDttl�T<4D�,tTt\\tt|�$d$lD4T|L,d\$
L4���d4$dd,l$|T,�4d\|\ll�,4<\d,$$lt4DTTt,,\L<<LlDDd|D<Dlll$\dDT$4$<TTDl,,Dt<,4l,Dt4T\4D$TDDd$d,\D$,ttD\t,d|4t|dl44\dT4DlL,,$|\dD,L4TtL<TdT4td$,l|D,T4D|dD$4LD$$Dl4Dllt$$T,<ttT$$,,ll<DT4d\�4,|T<\<|lt,$D,dDL\4T$4|LJB^^BPVzzz44 	�������"�%�'�*�-�0�3�6�9�<�@�D�H�K�O�S�W�[�_�b�f�j�n�r�u�x�{�~�������������������������������������«ƫʫΫҫի٫ݫ�������������	������!�%�)�-�1�5�9�=�A�E�I�M�Q�  			

					
	

	
		




	



    
								
			
		


		

	


									Q�[�e�o�y���������������ɭӭݭ�������#�-�7�A�K�U�_�i�s�T$|\tdD�L\�$d$l\4�<�$dT\�<d���Tt$D�l$|��<l�4Tt,dd4�T\$L�t|$lT$|d�l$�|�|DD|,d,T�$�,d\l,Dl�LL|4��4�|�$t4lDT|\$T|�|Lt$�<d,�\t$�\l<�t,l,�d�$��|T�l$�D�t$<dt�L�|4�lDT$�t$Lt�dD$t�,lT��4d\l<�,�|�dd�td$l<L�t�d<�tD|4��\<�4l��<t|,|T��îͮ׮������	���'�1�;�E�O�Y�c�m�w���������������ǯѯۯ4|<TdtL4<Dl|D,4<dl|,D$,4<Tdtl$,T\|tT,4<\d|t$4T\l|$|$4<Ll|$<DLT\d,\$4Tt|,$D\dllt,4DLTltd$$L\tdd$$44DD\$<<L\|t$4LdltL|<<Ll|,l$,<T\lL4$,Ddtt$\$TTlt|$$4DTltt$,<\dlLD<\\t|l,4<dltD$$Ldll|l,,,4TdlD$$LTllT4<T\l|<$4\l||,$$\ddl 	").7<CHIJQV[dkpwx}��D4\tdD�$\T\4�T  D�<<d|4�Dl$$$t||�L�d�tDdT�L,T\l$t\  dd�t�<$\D\�dl�t4,TD4D,D,tdt |<lt�,dL,,\4,4tD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �5
����-���.l- ��=�}�������Ӄ_�()*./0+,-������������ԩ ���� !����#��+�0�����Y��[� 	� �憥���� *� �� o� ���5`� � �������F !����)�<8�
����'���(�}����~���� ������+� �'�-���. 5�� �)�! È 	� �� �)� �
�ͦ<ʼ寥 8�
�����)�+Ȅ,� 8�

e,����-���.е�5 ��`�;�@���L����@���� ���`�0�0� �<�  �����e<�� ��੅�:��0��@�� �F�� �L��@�S����X���� �`���� �#��p���e<
��^��-�_��.���0�-�  �������`��)������0 k�` ����`�`�
�ݩ �`�0���K�O k��5�<�@�� ��` �� *� ۍ M� �� `� �� � ^� (�`�F�}�G�F���G��o� �G� ��F�F��� �F�;8��;0���; �� !��̅+�8�)�i�-�?8�)�i�. 5�� �!���! Y�����-���.�� È 	� �`��)�E����;�:��5��6� ���@�;�:�%��<�	������ �J�=�
������4`��4`��_���`��)�/�;�,�@�;���
��� ��`�5� �s�� ��`��5 ��� �s`���; ��� ��!������" щ ��`     �E
��p��-�q��.l- z�����z����Y�� �� �J������(���� �  ���E`��)��J 6��J���E`�0�` =���5� �E�<�@�� ��`�#��6 ��<�<��� �<�̓�������4��`��4`                                                                            2(��0�D�Z�m����]��� �� ��` ���0����� k��_I�_ ׅ � l� �� 1�`� ���M�N�)�:� ��4� )��� )� � )��� )� � ���% ���)E � �
� ��� ��`����悥 J�3J�ZJ�L����)����`�)��έ?��� ݈� ��� ��`��)����`�?)�Ф�ɒ�� � � ��`��)����`�?)����� 	�� �� ��`L􄭟)��4��`�)���?�z�� �� �٩4 ��`��� ��;���; ��`   Ȇ� �2�-H�.H 1���0h�.h�- 5�� �!���A���� �� � ���`ɐ���!)�� �P�!�+�i�ÆH !� È 	� �h�' r���`)�ɀ�̱!ɀ���Ɂ��5�5�s� � � ��)�� ���!�+ !� È 	� ����� h����
�6��@���� ���`�0�0� �<� �5��慩�5���� � � `
� � ��)���)��)�?� �'�)��2��)��?)�#���?)����}υ�-�?}Ӆ�.� `��%�ƅ&`� �"�:8��!�
��
�!�"�� !����Y��"i�+ 	� ��Y����!i�+ 	� �`� �"�<�!�
��
�!�"�� !��̅�[��"i�+ 	� ��΅�[��!i�+ 	� �` !�� ������Y���i����Z����<i�+ 	� �Ɔ�����`������������� ���;�� !����燅�+�[�������� 	� �憥����`�����+�� 	� ����燅�[����� �©��C��-��. �����燅�[����� �¦�����C��-��. ��� ��� �C���-���.� �  ��` 5�� � �!���0���!��� `�@��-JJ����.�� ���`�0� i�-� 8��. ��`�0� i�.� i
�- ��`�0� i�.� 8��- ��`�0� i�-� i
�. ��`� �!��"�-8�JJJe!�!��"�.8�JJJ���!i�!��"���`���'���'� ��!�����'�
��
�'�$��'�# щ ��`	 	 	    	� �!u=�=�
��
�=�>����q�Bٳ����Aٕ���q�: *�`� �D�;�����D�D��)�������`���5� �E� � �� ��`�F��)0��;���F� �G`� ������`          � ��P������)�� �d��X�����`�5`�0����	�@I�@`�@I�@`�0� �M�N��J�,J�OJ�r� ��
���� ��`� )�� ݈� ����N`� ɒ�
���� ��`� )�� � ���M`� ��
����4 ��`� )�� 	�� ����M`� �z�
���� ��`� )�� �� ���N`�eM��?eN�?`�0� )�� y���� i�`              � �L��0�@0&�`�`�`��� �`�P�����
�0��L ���0�0��ͥL�	 � 1� ��` /��0����� k��0�@I�@� eM� � eN�  �� ��`� �M�N�0� )����)���M`����� )����)���N`�����p� ����J�&J�DJ�c r��0� �z�p��憽�/�k�i ��Le� ���0� ��pН憽��� ��LG�LU� ���0� ���p��憽������ ��LL� ���0� ��p��憽�/� ��L`� ������ ��� �� ��` ��� ���� ��� ���� ��� ���ۦ0�����p����Le���I<��` ����/� r�� ��Ш ��� ��4Н ��� �	�� r�� ��0�����p����LL�LG���I��`�0� )��)� )�� � i�-� i�. 5�� �0�!����0`��0�P�"i�Pɀ�)� �P�� ����� k�L�� �i��� � �0�iɴ�� �0�0�0���`��0��H�@���	�0�0���` ʏ�-e.�������� �� � ���`�����0H��0 k�h�0�0��к�� k�L@���H�@����P� ���H�H���`4��0�@0�0�0���`�H�� ʏ�-e.����� �0� ���P�H� �ש�P`�0�H��=�)�KJ�J�)J�4�4� � � �� ��`� ��`�� � � ���� � � �ڐީ� � � �̰� P��H��)J������`����5�
�_� ���`� � � �� ݈`� � � ɒ� �`� � � �� 	�`� � � �z� �`����)� � 



e ��U��p`� �-�.�0�H��8������@������������-�-�-�8������������������.�.�.`� �-�.`��)�e� �P�Z���T���-i�����.i����@0��8�������8��
�%���!�� �ڊH 5�� ��!�+ !� È 	� �h��P����`� ����� ��`�����Ȑ� ���H��i����i����0�@���
�0�0� ��.��8�������8��
����ڽ���ө�� k�Lϐh�H���-���. 5�� � �!�+ !� È 	� �h�L��12345`�Y��J�

i��/��+ !���!�" 	��!�܅#�"�$�-�+��)��*��&� �/�%�(�� %&�' ��'/�/�%�%��� �%�/� �© �/�#�� %&�' �L���#�''L��&&�!�#�(�(�������+�
��&� �(�)��*� ���$��8�-���L_��.�LU�`�(8�%��	0F'F'���`''���`��0�@0����� k��0�0���`
 #(-4<>IKQ_din�O�K�:����)� ��P �֤<��


e �� ��-��. 5�� �!�j�-i���.i����@0��8�������8��
�=���9�� �ڦ �P�-���.���h)�� i��!� �X�i iͅ+ È !� 	� ��O�h`���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5
����-���.l- �D�u�������ץJ�

i��I����+ I��J�J��� �J�5`�J

i��O��8�J��
i�+ I��J�J��ک �J���5`�0��
���4��6`�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5
����-���.l- )�f�𘸙()*./0�������ԩ ���� !������+�!�����Y��[� 	� �憥���� *� �� ���5`�@���G��0�J��V�?��_������� � ����@���� ���`�0�0� �<�  ��`��)������0 k�` ����`�`��ݩ �s�`�0�� k��� ���5` �� t�`��0������ �� ��` ������ k��_I�_ 8� l� ��`
 Ȇ� �4 5�� �!�+)�ɐ�%�!)��3�H� �!�+ !� È 	� �h�' r���`��-�� ��;� ��` ���5� ��� � ���`�0��@����0� �<� ���`�����4��6�@�;�`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5
����-���.l- �>���@� �����0�H� �e� ��� ���5��6`e}�)��>&������6��4�t�:� �=�>�?�@�A�B�q �` ������I����<�� ���)���ߩ �0 k���6`�����6`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������DTl\l|�4\\4,�lD\�ld$,\,|$,TTlD|\�dD<<T�<4��L$$|Tl4T$D\\|T|<4�\$$l4<4|d4|,�\l\T4�T4t�,TdD$��Ld<�tLTt4\4T4|t4dDttl�T<4D�,tTt\\tt|�$d$lD4T|L,d\$
L4���d4$dd,l$|T,�4d\|\ll�,4<\d,$$lt4DTTt,,\L<<LlDDd|D<Dlll$\dDT$4$<TTDl,,Dt<,4l,Dt4T\4D$TDDd$d,\D$,ttD\t,d|4t|dl44\dT4DlL,,$|\dD,L4TtL<TdT4td$,l|D,T4D|dD$4LD$$Dl4Dllt$$T,<ttT$$,,ll<DT4d\�4,|T<\<|lt,$D,dDL\4T$4|LJB^^BPVzzz44 	�������"�%�'�*�-�0�3�6�9�<�@�D�H�K�O�S�W�[�_�b�f�j�n�r�u�x�{�~�������������������������������������«ƫʫΫҫի٫ݫ�������������	������!�%�)�-�1�5�9�=�A�E�I�M�Q�  			

					
	

	
		




	



    
								
			
		


		

	


									Q�[�e�o�y���������������ɭӭݭ�������#�-�7�A�K�U�_�i�s�T$|\tdD�L\�$d$l\4�<�$dT\�<d���Tt$D�l$|��<l�4Tt,dd4�T\$L�t|$lT$|d�l$�|�|DD|,d,T�$�,d\l,Dl�LL|4��4�|�$t4lDT|\$T|�|Lt$�<d,�\t$�\l<�t,l,�d�$��|T�l$�D�t$<dt�L�|4�lDT$�t$Lt�dD$t�,lT��4d\l<�,�|�dd�td$l<L�t�d<�tD|4��\<�4l��<t|,|T��îͮ׮������	���'�1�;�E�O�Y�c�m�w���������������ǯѯۯ4|<TdtL4<Dl|D,4<dl|,D$,4<Tdtl$,T\|tT,4<\d|t$4T\l|$|$4<Ll|$<DLT\d,\$4Tt|,$D\dllt,4DLTltd$$L\tdd$$44DD\$<<L\|t$4LdltL|<<Ll|,l$,<T\lL4$,Ddtt$\$TTlt|$$4DTltt$,<\dlLD<\\t|l,4<dltD$$Ldll|l,,,4TdlD$$LTllT4<T\l|<$4\l||,$$\ddl 	").7<CHIJQV[dkpwx}��D4\tdD�$\T\4�T  D�<<d|4�Dl$$$t||�L�d�tDdT�L,T\l$t\  dd�t�<$\D\�dl�t4,TD4D,D,tdt |<lt�,dL,,\4,4tD���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �5
����-���.l- �&�� ���u�5`  0@�02�G�u0C�)����u�7�u�� ����u�u��&��6�<��4��t`�4��6�<�u���
���t` ��`bkt� tPY�P          ���#�M�$�	�%���&��)���)�
�'�
�(��6�'�w��)  ��(��'�#i�#���$��`�5
��䀅-�倅.��6l- ��m�� �@����0�0� �@� ��� ���5`@Xp��)�������� �0 k��)�/)����
����� �� �0 k����� ����`�)�����5�� ��`����@� ���4��6� �=�>�?�@�A�B�q�t�:�@�; �`����������������������������������������������������������������������������������������������������5
����-���.��6l- �e���߂��'���%�Յ&�J�$���#�5�'�	i��)  ��'�	�#i�#��`T�X�^�����������������
��N��-�O��.�b��'���%�Յ&�R�$��#�5� �(�(�-�)  ��'��(�#i�#��`��'���%�Յ&�Y�$���#�5�'�< i��)  ��'�	�#i�#�� ��`�0����4��6`���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������5
����-���.l- 1�4�ȅ��f������������
��6���%�Յ&�F�$� �'�J�L���'���)�&��#  ��'�'����5`������������������˄Մ���������������� �������������� ���� ������������������������ ��������� ������������� ������������ŉ��� ���������Ħ��� ���� �������	

 











	��)�` y��M�$���#� �(�*�����'�
��e��!�f��"�(�!��)�L�
����i}�)  ��'��#�#�(���*�*)���6�R�$�J����#Ф�
�#О�L�	�����`�5�LI�L�J�J� ��`�L��J���)�����`� �J�����5`�5� ����`VX���)�� y�� �(�*����$����#����'�
��e��!�f��"�(�!��)����i}�)  ��'��#�#�(���*�*�����6�����`�5� ��`����)����
���`���%�Յ&�J�*`�5
�����-����.l- ��?�n����������� � �� ����%�Յ&�M�$���#� �(�(����)  ��(�#�#�(���X�$��#� �(�(�����)  ��(�#�#�(����5��6���%�Յ&�P�$���#� �"�<�!�
��
�!�"���"i��)  ��#�#�!i��)  �`���%�Յ&�^�$��#� �(�(�����)  ��(�#�#�(����5`�03)�� � ��)�/�)0�))��<���<L���<�<�����<L����4�6� � `�������������������������������������������������������������������������������� �'��(�4����<8�
i���λ��!�É�"�����%��&� �!�$� ሱ!�#� ሱ!�) ሤ4���� �*�ǻ�/� �!�����)�+Lv� ሱ!�+ ሱ!��+��,�4����� �+���' � 	� �� ��/�8�*� �$�#i��#��$�#��$���$��*8� 
e#����,Щ �L^�`�!��"`�'��(`LNPRT� �'��(����!�É�"��%��&� �!�$� ሱ!�#� ሱ!�) ሩ� �*��/� �!�����)��LR� ሱ!�� ሱ!�����,� ���� �L��i��' 舥�iͅ+ 	� �� ��/�8�*� �$�#i��#��$�#��$���$��*8� 
e#����,Ф �L:�`�9���`�#���|�5�����Y��ڒw��ߔ��M��×��K��Қ���E��ݞ��i�)��ߢ~�@�����Z�N�O�E�D�C�@  �	$-6?HQZclu~���
%.7@.R[.mv���&/8AJS\enw����'09BKT]fox����(1:CLU^gpy���   )2.DM._hqz���  !*3<ENW`ir{���#  "+4=FOXajs|���,  5>Gbkt� tPY�P� ���������	����������������������������������������������������������������� �����������  ������ �����������@  �@��}�� t����P��V  V�V  V�V  V��Yt��V  V�V  V�V  V��d�IY��V  V�V  V�V  V��Y�;�V  V�V  V�V  �V�)@� �� 
     ��         	   	  �� �	�'
   
   � � � �	��  
� �          �  	  	    ��@� �
           � 	 �  ��   	     	��  
 ���     
   	    �  	 �
�   �
   �  �� �  �@� �
  �  � �
    �  	 	  	 
   �� �
 � �����
 � �	 	  �� �
�      �      ���@� �� � ���      ��      	�	  �	���  �  �   ����
�  ���  �  � �@� ��     ��    
��	��  ��	      
����     
   �� � ���  � � ��  ���  @� ��     � � �� 	 �  	 ����� 
    � �	� ��
  �	  �  �  �   	�  ��	�   � �@� �     �      ���
  
 	  ��	     �
�	 
 
� � ��   �     �	  � ����� 	��@� �� �   �      ������ 	   �  �   ���  ��� �       	� �	 �  �	�@� �   �    	  	� 	 	� �  �
�
   
   � �
  ��� � 
  �	  �� �  �    �� ��      ��@� ��     ��
  
�    	   �     �    �  ��    �    
�	      �	�   
�  ��    ��	      	�      ��	�@� �6�7�6��67 8 7�6�8�8�7�
6 6  8  6 6�
9�	6 6 9 6 6�9 9 9 6 9 9 9�77 7 7�7 7 77  88 8 8�8 8 88�	6�	6 6�6 6�@� �7�6 6 �6 8 9�	7�9�6 777 8 �6 9�888 9  7�6�9 97 8 6 6�7 7  8�	6 8 8 6 �6��6 9 9�9 6�6 9�6�9 6�6 7�6�8�@� �9�	6 6 6 9  9�79�
9  9�8  9779 9 9 9  7�9�889 9�9  8�7 7�9 9 9 9 6  98 8�	9�9 779 977 9 6 6 88�88 9�9�9�7 6 9�9 6 9�8�9�9 7 9 9 9 9 9 9�7 8�	7 9�8 6 9 9 9 98 9�@� �9 9 9 7�7 9 9 9�8 9 8�9 9 9�9�9 9 9�7 9 7�9 9 9 8 9 8 9 9 9�
9�
9 9 9 9 9 9 9 9 9�
9�
9 9 9 9 9 9 9 9 9�9 9 9 9�9 9 9 9�9 9 9 9 9 9 9 9 9�9 9 9 9�9 9 9  9@� �9�9 7 9 6 97 7 7 9�8�8 8 8�9�9 9 7�9�9�8 6�9�9 6 7�6�9�8 9 6  9�9 6�9�9�
6�9�9  6�	9�7�7 7 79  9�9  9�8 8 8�9�6  7�7 6 6�86 8�99 6�9�@� �7�9  7 8 6 6 6�8�9�7�7�9 7�7 8 6 8  7�8 7 8�
86 9 8�7�7 8  77 9  9 6 6 8�88�9�7 6 9 6 9  77 8�9�9  88�99 9 7�9�9  9�8�97 9 99 6�9 77  98 9�7 9 88�9�8 9�@�   7�6�8�9  6�9�6�6 7�9�7  9  9 8 7  9 6 8 6 9 998  9 7�8 9 6 9 9 7 9  7�9 7�8�899 9 8  6 9 99�9�9 99�6 999�6 6 6�9 6 �
6��6 6�@� �97 76 9 6 6�8 8�9�9�9�7 9 9 6 6 9 7 798�9 8 8�9 6 9 7 9 9�6�8��9 6�6 9 9 7�9�8  9 9 9 6 9 9 9�
7�9�9 9  9 9 9 8�9 7�6 8 9 7  7 7 7 7�	8  8 8 8 867 7 6�8 8�@� �7 6 6 7 9 9 9  8�	8�
9 9 9 7 9  6 96�8�7�9 9 9 9 6 8 6  6��6 9 9 6 76�9�98�79 97 9 9 9�97 8�8�9�9  8 9�9 677�7�88�8 99 6 6 99�9 9�	9 7�9�9�9�8  @� �9�6 9 9 7 6 9 7  9�8�9�8  9 9 6�7�7�6 68 9  8 6 7�7 8 9 9 99 9 9 68�9�	6�6 9 9 9  9�9�9 9 9�6 9 9  9�7�7�7�9 9 89 6 8 68  7�89 9 7 6 6 6�8�@� �:�:  ; A>>? =>>? =?  ;  < ;�<�; =>? =�>�: ;�=>? ; < =>? A? : @�;�;  ;�=? < @ =>>>B =B =>�@A>>? A>>>C =>>>?�;�;�;�:  @ ; A>>B�D>>C ; @  ; <�@�< ;�@;�: =>? :�;@�<  =B�D?  <  @�@� �:�:�@ ; : : : : : ; @�< ; ; ; ; ; <�:�; ; ; ; ;�:  < : ; ; ; ; ; : <�; ; ; ; ; ; ;�A>B < ; ; ; < D>C  <�; ; ;�<�A>? ; ; ; =>C�A>B�< < <�D>C  <�:�:�<�: ;�; :�AB ; =>>>? ; DC�;  ;�;  ;�< =B =>>>? D? <�@� �:�: : :  =? ; : >>>C < ; ;@�; ;�;�; D>>C =B <  : D?  ;�=B�<�; :�=>>�@�< ; : =?�:  =C�; <�@�DC  <�<�@ =>?�D?�@�@�:�: : @�AC <�< ;�DB�@�@�D>?�:�:�@ =>B =>>>? ; =>?�;�@� �: A>C : AC : @ :�< < ; < DB <�< :�;�:�;>>?  < @ =? @ < @ <�=? =C�=>C�; A�>C�<�AC  ; ;�DC�DB  ; ; =?  D�>�; ;�:�A>? =B ;�< =>? @ <�DC :�
: =C  < D>>>C =?  =B  <�@<�@�@�=?>@� @�@ : A? : @ : =>C  @  < ; AB�;�<�@  ; <  : < :�=?  =B�@;�D>?�:�:  ; :�=>>B  =B  ; < =>C�AB�; @ @ @  :  <  =>? <�; =>C�;�; =>>>? @ =>>? <�<�
:�	=? =C  : ; =>? :  @�;  < <�D?�=>>B�@� �: :�A>? :  : @  < < =? ;�D? <�<�
=>? @ @�A�>? :  :�: ;�;  ; A>>? < ;�: ;  < <�< =>>B <�A>?�:�@ =? <�=>>? < :�	:�; : =>? : ;�: : @; ;�; D? =B ;  ; < : : ;�DC ;�< ; < =>>?�< D?�;�@�@� �=>? =>>? :>C @ :�:�<�;  >>C : ; =>?�: ;�< < <�A>? < <�
: ;�	@ =>>? < < =?  AC�:�
DB >>>? ; A�>?�; ;�: =>?�@ =>B <�;�=>>�; =?�A�>? @ <�=?  ;�@ @�< =>? : =>C�@�;�;�@� �: : : =>>? @ : @�< < ;�;�	; A>>? A>B :  >C A>B <�<�;�< ;�A?�=>B�;  AC ;  :�=>B  DB < =B =�>�>? A>? A>>>C  A>>?�;�;�<  ;�: ; @ ;�; AC  < ;�DC =>>>B DB�; :  ;�@�@ < < AB =? @ =>?�;�@� �>C A�>? A>C A>>?  < ;�; < <�; =>>? ;�:�: <�< =>? D>>@;�=?�< =>?�=>>C�@�=>>?  @ <  A? @ =C�@�;�D? =C :�:  < @ @�< < A>B�:�<�=? =C D? =? :�
;�; A>>> =>? D>C  =>>B <�
;�@� �: @ =C @  =>C : @  <�;  @�< ;�=? D?  @ @  <  : @�@�@  =B�: =?�:  @  @�: <�=>B :  @�;�
; @  :  < A>? =C : <�@;�<�< <�=B�@  =>?�=? :�@  @�	; AC @  @  @ @ =? @; DB�@  AC�;�@  AB; @ @ : D? @�AB@;�;�@  ������ FHJKNOR TUXY\]`a �� GILMPQS VWZ[^_bc ������z{����|��� �������� ���}��� �������� ���~����y �����������y��������y��������dgjmpsv��������ehknqtw��������filorux������������ ���� ��������@� �E �E �E EEE  E E�E E�E E  E E �E �E E E  E E�E E  E E �E �E E  E E E�E�E �E	 E  �E�EEE E��E�E  �E E�EEE EEE  E�E��E �E EEE�E  �E�@� ��E EEE E E E  E�E E E�E E E  EEE E E E �E E�E E E E�E E E  EEE E �E E E E�E �E �E EEE E�E E E E  E E E �E E�E E E E��E E E E E E�E�E E E E E��E E E E �E	�E E E �E	 �E�@� ��E
�E E�
�E  E �E �E�EE E EE �E EEE �E E�E�
�E EE  �E EE�E  E  E��E EE E  E �E�E��E �E  E EEE E�E�E  E�E E�E EEE E EE E E�E�E�E �E	 E E  EEE�EEE��E	�@� ��E EEE �E  E�E E E��E E E E �E�	E E E E  E  EEE EE E E E EE E�E E E�E  �E E E �E E  E�E E  E EEE  E EEE EE EE E�E�E �E �E E�E�E �E �E  �E�
EE  �E
 �E�@� ��E EEE �E  E�EEE E�E  E �E EEE �E EE�E EEE E�E��E E E EEE E E��E  �E �E�E��E  �E EEE E E�
E E�E E E E  EEE�E�E E  �E��E E E�EEE�E E  �E EEE �E E�@�           �� �        ��          � �           �	 �   �   �    ���   �   ���          �  @�          ��         ��          ��          ���          �    ��     ���	   �	 �        @� �
          ���       � � �       � �      � �         � ��     �  �    �	  �     �   �	   @�    ���     ��  �     ��   � �  ��    ���   �
 �    @����  �   ��� ���       � ��     ���   �  �    ������         @ �*VeeXywg {euVXs�Wffizt!|fxWio���p���� "-8G�#.9H�$/:I�%0;JYh�&1<KZ������'2=L[j�(3>M\k�)4?N]l�*5@O^m�+6AP_n����������,7BQ`��CRa��
DSb��	ETc�vFUd�                           � � � � p p p p \ � \ � � �          � ��[>[>���          � � � � p p p p � � � � � � � ���������09090909LL�L��?��pUp�p�p�\�ܪܪܪת�����������j�j�Z�ګګ֫���U�������������    ������������  @@�����?�?�?�? � � � ������G�A�A�@�_�          ? � �������s�����������U�����������U���{�o��_�ߪߪ_U����������      � �� ��������������P�P���o�___�G�W�}���������A|��  �� � �      ��U��߫ګ֪�������������j�j�j�j�Z������������������������         P ��������������������A_@P���������                �|?W�������_�ߪߪߪת�������j�j�Z�ڭګ�U�������������        ���������?�?�?�?A@���� � � � 0 0 0 0                   ��_U������������������������������U����_�ߪ_U������������   � \ � ���� ���������p�p�p�p�\�ܪܪܪת����WU�������� � �               ���   ��U��ߪڪ֪�������������j�j�j�j�Z������������������������  ��UU��������������  �?<?<?<?<?<�ڪV�v��������W�������>�;�/          �?��       ���U����������_�ߪߪߪת���������j�j�Z�ګ�U�������������  � U5�֪Z�j�j�������j�j�Z��j�Z�����Z�j�j�����U�������������           0�      ��UU�����������  <??�?�<<<<�j�UU������������������          �p=p�\���������������~�{��_�ުܪ��WU������������        �?������   5 � Zjj�=��������j�j�Z������~�{�~��_�߯\� � �         ��|UW������������U�U�U�UU�U�U�U�V��߶��������W���������;�/        �?<????�??��pUp�p�p�\�ܪܪܪת�����������������j�ګ�����U�������������  ��UU�����������j�j�j�j�Z�ڪڪڪ֪�������������U�������������        �?<?<?<�? ? �?U��_����������  �??????????��j��U������������+� � � � �   ? � �����_�������������������������������\����? > ; /         ?<?<?<?<?<?<� ���5�����Zjj?j?j�j�Z����������_�޾����׿�+W � � � �      ��_U���������j�V����j�j�j�j�j�j�j��U��������UU������������        �?<? � ??���UU��j�j�j��������ܪܪp�p��� ���U����������ZU�������������  ��UU��Z�ڪ�U������������� � . ; �U=��j�j�j�U�������������        ??????????<��\?�������������֭Z�j������������j�Z��j�V��������������+�   �\?��������������������p�p�p�p�\�ܪܪߪת��WU���������        �?0? ? ? ?0��?U������媽����j�j�j�j�Z���ֿ���������������.��� /        ��UU���������V�����U������jUj�����ZU��������UU������������      V�V�Z�:�  � �      ? � � � � � ? > ; . +                            ��U��ߪ֪���U�������U��Z�ڿ����������߾���/����������������       ����� >�.�??+ ���/. = =?.�>�� ��� �   =./���+     ���������������  �????????????  �?<?<?<�??<  ?<?<?<�??<?<?<??�? ? ????�  ���������?��  � � �� � � � ��� � � � ���������?���������?�  ��������/���  ��������?�?�?������������?�?�?�?�������  ������ � � � �  �������������� � � � � �����������������������  ?@?�?�?�?�?�?�  ������   �??�?�?�?�?�?�?�?��?�?   ������  �/�?����������  ���������������������������     � 
� PRU����쐬���������U WUkU����   � �               ��
*  @ UTUU�����k�k�k�k�������U� �U�������  ����         � ���� P�U�U���������������������������� � ����      ��*� T [U�����������_��k��FR@PT�k����_�����������               � ��?�?<�����UUUU�U����������������������������������������o���   �� U������?�� � � ��?�����V�j���UW  BUKUUU/U/U/T/T�T�T�P�R�RϪ�  ����  ��  UU������<��� ��� �����UUU���UU      UUUU�� RRERRDQ ��UUUU����  ����  �
 �  U�V�������o?k�[�Z��V�V���UU      UUUUZ�p�q�p�q�q�q�p�_�UUUU����  ����    ��      ���A�U���������UU����UU    TU�j�~�~�~�~��_�_�_�_�V������   ����      �
 �    *�/�o�[�[�V�V�V�UU����UU  UUUUUUU�U�U�U�U�U�U�U�U�U����� �    ����        * �
 � � � �ooU[UZ�U*�U��U��?��������>��������������������������             ( � h �  ��
TU�����?�������_��k�[�VF@P�+����_�����������T���
*`@�Vՙ���uU��� �W����������������������������������� o���W��+ UZf����k�?[���Z�  0?<�����  ?<�<�????<?<?<�
  �U�U�j������/���3���3���/  �??????????�?�/���� � ? �?  ? ? ? ? ? ? �?  �?? ? �? ? �?   B@<V�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L��Lh�L��L�� �0��)�	�0�0� ��`����� ���@�3��JJJJ)�1� �2���2 �L�� �0����
�� �� k��0�0� ��` ���-� � �������-���.� �  ��` ���-� � �������-���.� �  ��` ���0�@��-��.�
���������` @�� @�� @�� @�� @�� @�� 	@	�	�	 
@
�
�
 ���3
���!��"��#�1)����#�1� � © �&�*�$� �!�(�1)� G� p¤*� �2�.�($�+ �¡%+($����ȥ&�+�$ �¡%+$�L����+ �¥($%+����ȡ�+ �¥&�$%+�� �&� e#� �*�-�LC��.�.����1������ e-e-� �
� 8�-8�-�  ��L;�`�@��0� JJe���� e�� ���`�.�-� � �1����	� e-� ����	� � 8�-� `�()�JJ�)JJJJ))�)�()

)�)�(





)�(`�0� )��(&&(&&���`��,�+%,��+,�+,,��`�i0���`���`	�Ɔ�I������>�bÆê������:�^���^Ŗ�T<��j�������U�U�Uk������T�T<������j���U�U�U����j��T�TA��o��o��o��WU�WU�����o��o��oTATA��~��~��~��?WU�WU���?��~��~��~TA�Uj�}�}�}U�U��U}U�}j�}�}�iUAU�U�}�}j�}U�U��U}U�}�}�}j�iUAUUEU�V��f��v�U�U����U�U�v��f��V�UEUUEU�W��g��w�U�U����U�U�w��g��W�UEU       <  7 ��pU�� 7            <�w���U�\U5]UuWU�WU�]Uu\U5�U�{��<�UUUUUUUUUUUUUUU����oU����_W_}}�W�WU_�U��u�_�}��WU_�_��u�W�}�W�WU_�U��u�UU}�W�WU��U��u�������WU����_���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�W}���W�__���}��}��}_�}_}�}_}��}��}_�U_��}_���}��}_�U_}u}�}��}��}_�}_}��}]����W�_��w}_UUUUUUUUUUUUUUU ��?�  �?< ��U� �?� � C� �7 C�5 �? _ �_  � UUUUUUUUUUUUUUUU���]��_U������}�_�}��UU�����_�}�_����_U�����_�}�_����UU�����_UU�_�}��UU�����_�}�_�}��_U���_�}UUUUUUUUUUUUUUUU                �?W�W�W�W����?�0<87�3��[��?W�W�W�W�W�W�W�W���UUUUUUUU�������?W�W�W�W�W�W�W�W�W�W�W�W����?��WUWUWUWU�������?U�U�U�U����?WUWUWUWUWU��������WUWUWUWUW�W�WiU�U�U�U�U����?�?U�U�U�U�U�U�U� l&�l&� ?    �?\5\5�? ?    �?�?�?�? ?   ��}=mz^���W���WUWUWUWUWUWUWUWUU�U�U�U�U�U�U�U���UUUUUUUUUUUUUUUUUUUUUUUU��������WUWUWUWUWUWUWU��t=mz\���W���������������������U�W�W�W�W�U���������W�W�������������������������UUUUUUUUUUUU����            ����Uu]u]u]U_u_u}����������������������������������� ��� �?��?��������?�������� ����� ��� ��������������� �������� ���?�?��������������������������������������c� ?��� ������Z� ����������_�_��������u�u�u�u�u�u�W��]_]_]]]U]W]___��W�����������W����0��Â��Â��>833333>8������������������ ��������� �������������� ��������������������������������� ����� ����� ��C}mz^:��W����L5\6\�\��:�:]:�:_:l:l:\:\:w����Gqmz\:��W�����������y99999999�:���������^�� �� ^U^U����   ��  UUUU����   ��� �U�U����� ��?�S�S�S�S�����  �� UU��999 9U9U9�:�    �@:999999� \U\U����  �*V�F�V���V��* � ��������?�/�/����/�?���� �� � � � � � � � ���������������������������������������?�?����������/�/�?�?����������?�����������������/�/�?�?����������  ?�?��������������?����   �?�?�?    �����?   � � � � � � �����������?��� � � � � � � �  ��?����������� ��?������������ � � � � � � ������� � ?    ��������������������������������������� � � ��������������?�?�?���� � � � ����������������������� ��?�������������������������?�� ���?����     ���������������޽޷�����}޷�����}ܷ�� �     ��������Z��������������}�������}�������}����� �o�o�n�~L���������������������������������������U�  V�V��������������>����>���;����;��������U�fPZ�����������������0 �� � �@�0 ����������������������������������������￿���������  
 � �
�/�/�k�k�����n�n�����n�n�����n�.��    llllllll�ll�lo��l~�nk ��_DYDVUDVYDUUEUEUUUUUUUUEUUEUUEUYUVWUWV_�\�\��� D�UDUQUDUQTUQTUQUTUQUTUQUTUUUTUUUTTUTUUTUETUETQETQ_TpQ�T�U W | �    U�UUU�UU5U�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUD_��  _�U5U�  ? ��U?E51U41D41U4U� 5�E1U41E41E4�D4�?            5 �         0 � ���l�lkn�~[�[�olol[lWl\lllo�_�\~�nll�nl~��l�lolll��U�U�U�UU�U�U�U���
 ���UbUb�b�b�  �?<?<?<?<? ? ? ? ? ?<?<?<?<�  �?0?0?0?0?0?0?0?0?0?0?0?0?0�  ?0?0?0�0�0?3?3?<?<?0?0?0?0?0?0  �?��������������  ���������������  ?0?0?0?0�0�0?3?3?<?<?0?0?0?0?0  ?0?0?0?0?0?0?0?0?0?0?0?0?0?0�  �?? ? ? ? ? ? �?? ? ? ? ? ? �?�<<<< <  ����  ���bUbUbUbUbUbUbUbUbU�U��
 ��      ��  ��UUUUU��������������������UUUU��  ��      ��  ��UUUU�_�W�U��  ��UUUUUUUU�W�_�W�U�U�U�U�UU�_���_U_U_U�WUUUU��  ��      UUUU��  ��      ��  ��UUUUUUUU���* ���U�U�U�U�W��_�_�����U�U��U�U�U�U�W�W�U�U�UUUU��  ��      U�U��� ��*          ��
 ���UbUbUbUbUbUbUbUbUbUbUbUbUbU�U��
 ��      ��  ��UUUU�����������������UUUU��  ��      ��  ��UUUU����������������������UUUU��  ��      ��  ��UUUUUUUUU��_�_�_�_�_�_�_U�UUUU��  ��      ��  ��UUUUUUUUU�U�W�W�W�W�W�UUUUUU��  ��      �* ���U�U�U�U�U�U�U�U�U�U�U�U�U�U�U��� ��*     �� ?<�   �? � �U��?� � C�C��_�_ �  � 7 5 ?      �"$(P�B�X$� ��000?�����?< ��0�Чڧ�S��? ��Ϝ?[��5G4��  �<��=�W���\%�� ��z����z�  ��?<<<�?���� �����0�������� ��� ���0�0���� ������� ����� �������0�0���� ��� ��� � ���� ��� � �������� ���0��� ���������� � �������?�?�?�?�?�?�?�����������������������0�0����������������� ���� � �0�0�0�0�0��� � �������������� ������� ����� ���0�0�������� �������������� ���0�0�������� ��� ��� � ��� � ������������������ �����������������0�0�0�0�0� ���������������������������  �*������  ******�*******  �������  *(*(�(�*�****(  �
***** ****�
  �** * �
* * �*  �
*(*(*(*(*(�
  
(**�*�*******  �
******�
* *   �*(*(*
*
*�*
*  ****�*�
���  ��? �? ���0 CCCCC000�� C  0 �     � p p \ \ \ � W ����U��WUW@W����� \ \ \ p p p p p � � �    �(�(�(� � � � � ��������~�~����������W�������ZUjUjU�U�V�V�Z�j          ��                     @ @ @ @ P   DQD�����W5���[�oU�����U�����U��U�PU�����>���;�������������U�U�ժ�������� � � � �     U U U UU U U U                             ? �0�T���eAe@iPPTƕ1e� <���+� ���Z�       � 0?�1�0?�?Ϗ���0��������������������������:�:��� :      �
�(� � � � � � � � � � � � �(�
         � ����<������������������������������ � ��>p�?p�>p�      ��|Z�j��������ꪺ�������������ޫ������ۮ�������������������������� � � � � � � � � � � � � � � � � � �      �������>���������������? �� ��_C����� \ p� ��� ��p_p���U�UVUVUVUVUV�U��������������������������{�_�UU_UVUVUVUZUZUZUZUZUZUjUjUjUjUjU�U�U�U�U�V�V�V�ZVZVYVU       ? ���?������������������ ��5�U�<< �   � � � ���p�_�E0�O?@@UUUUUUUUUUU����������������ի����w�]�W�U�UUS��555M�M�������������������_�W�t�s����n�z��Z�UUUUUU�U�U�U�U�����������������������������������������������������              ? � / � � � �������� � �<?��� ? 5 7 � � 4 � �?Ꙁ�
������������������������������P�A� ��������������������� �S�Z�EX������U��Õ
�
�
�
�
�
�
�
�*�*�*�*�*�*�*�*�*�*�*�*�
��
��*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�
� � � � � � �  ��  ����                � ��:
j������������3j�j��}��&�����������������Ϫ��?�?�?�?����뺫���������k���g�گ=j� ? : � � � � � � � 8 8 8 8 8 8 8 8 8 8 8 � � : � � � � � 8 8 8 8 8 8 8 8 � � � � � � � � � � � � � � � �*� � � � � �"�"�"    �j�      � � �
���� �                      8 0 � � � ��
****:�8�8�8�**��z_� 6  ���  ��
�
�        ��                                    �
�*�*�*�*�
�
�
� � � � � � � �
�*� � � � � � �*}�V�������������� � � � � � � � � � � � � � � �*�
� � � � � � � � � � � � � � �
�
�(�(�(�(�(� � � � �(�(�(�(�(�
D @ @A  D DA�A�BA�0��0�0�� "                                                                                 � � � � �       � � � � � � � � � � � @ � � � �  ��?<<<�?�  �������  ��?�?�? �?�?  ��? ?� ?�?�  �?�?�<?<�?�? <  �?�? � ?�?�  �?�? �<�?�  �?�? ?��� <   ��?<�?<�?�  ��?<�?�?<�  ��?<<<�?�  ��?<<�?<<  ��?<�<�?�  �?�?   �?�?  ��?<<<�?�  �?�? �? �?�?  �?�? �?�?    �?�? �?<�?�  <<<�?�?<<  �������   < < < < <�?�  <<?��?<       �?�?  ��?�<�<�<�<�<  ��?<<<<<  ��?<<<�?�  ��?<�?�    �?�?<<??<?   ��??�?�?<  �?�? �? <�?�  �?�?�����  <<<<<�?�  <<??<���  �<�<�<�<�<�?�  <??���??<  <<??����  �?�?��� �?�?  ����  ��� ��� ����� �� �    < ?��� ?    ���������?��  � � �� � � � ��� � � � ���������?���������?�  ��������/���  ��������?�?�?������������?�?�?�?�������  ������ � � � �  �������������� � � � � �����������������������  ?@?�?�?�?�?�?�  ������   �??�?�?�?�?�?�?�?��?�?   ������  �/�?����������  ����������������������������/���3���3���/ ���	����� ���`�
��T�	�U�
`�`������`���� �� �	�ȱ	����U���ȱ���������� � � ������ȥ�����L1�����ȱ���L1���ȱ�L1�HJJJ���hL1�ȱ� � �� h)� � �� ��� � ���� �� � �� �L�n�0!

�����8� �9� �:� �;� ���	��� � �0

�����P�( �Q�) ��R�* ��	��� �* `��d |!_� _= |� m�' r�t�z�x�|�d�0�(�������(�H�Z�x�x�@ @ !@ �  ! ����� � �@�@ @ @ !@ �  ! ����� � �@�@  �!@! �@�@� � � � �@�@ 1}@1}@ !A@1�}!h!@!!@!}  1}@1}@ !A@0�� � � � �@�!!@!!@@�@ !T!�!T!�A@  � �! � �!! �!!!@!!!@!T!!�!}!T!@!�!}!T!@!�!}!T!A@@   z�z�� !�!�!}@ !@!}  @ !@! ��  �!@  �  �1@!}!!@}�!��}!@@} � �   � !�!�!}@ !@!}  @ !@! ��  �!@  �  �1@!}!!@}�!��}!@@} � �   h !h!@!@ !@!}  � !�!}!h!}!@!�  h !h!@!@ !@!}  � 	� 	� !}!T1@h!}!�  ���	� 	� �}	@ 	@ !@	 	 �!@  	h 	h h	} 	} !}	� 	� 	� 	� !@ @	� 	� �}	@ 	@ !@	 	 �!@  	h 	h h	} 	} 	} 	} 	� 	� �}!�  	�	}	�	}	@ @�!@	h		h		} }	� �!@	�	}	�	}	@ @�!@	T	}	�	}T�@h}�  ~�~�A�1}hA@  @ 	@ ! � �!A@@ A�1}hA@  	@ 	@ !!@!h!}A�@ A�1}hA@  	@ 	@ ! � �!A@   �0�� � � �!!@!!}  !�  !�@ !@!}!@  !@!}!@  	@ 	@ ! � �!A@   �0�� � � �!!@!!}  !�  !�@ !@!}!@  !@!}!@  	@ 	@ ! � �!A@   �0�� � � �!!@!!}  !�  A�@   ���� �@@@} h !@  � �@@@} h !�  h h}�h�h!}	@ @ �!@T T@�����	@ @����@@} h !@  ����@@h  !�  @h}h�h�����!@�����@���� �`   j�j�T�T�!T �.}.}!�  ��!}!.T�T�!�  T�T� � �����!.  ����!.� ��!.!T  T�T�!T �.}.}!�  ��!}!.T�T�!�  �T�T �������!.  ����!. ��. �    6�6��  �@@@}�}@ �}��  �@@@}�}@ �  �@@@}�}� ����  �@@}�}  !@  �  �@@@}h}@ @@�  �@@@}h �   � ���.�� }T}T �T���@@T}T}�  .�.��	}1.T!}�	}A�\ 	�	}.1T	� �  A.  �	}1.T!}�	}A�} } 1���	T�@�  ��0�T .	0�}. .1ThT.�@�  ��0�T .	0�}. .1ThT.�@�    ����� 	@ 	@  @   � �   � � @ @ � � @ @ � � @ @ �p � � �  � � �  � � �  @p �  �@ @ �  �@ @ �  �������p �  ��� � �  ��� � �  ���@�p   ����1��!}!�!}!T!}!T!.!!}!�1�}!T!}!�"<1�}��A�  1��!�!�!�"<1��!�!}!!}1T. !!.!@�  !.!T!}0���  � � � � � �AT� 0�� � � � ������!}!!.1T. !!.! �! �0� !T0�� �1T.���.T1} "�  ����. .}. .}T � �0 T T�T T�} . }0 . .}. .} � �0 � �.}	 T�} . }0 � � � �� . �0  T!T!. } .0 T �T!�!T} . �0  � �!���..T  ����� �� � �� ���� � � � �	 ��@ �� �� � �� �@��� � ���� ��� !@    .�.�  	T	�T!}  �  N�N�����0� `�`���� � � �������-���.� �  ��`�9�� ���#��$��%��&�� ��i�9�)��i������`� ����
��`�%��&��+��i�������-��.`xآ�����& �� �� �� �������� �� ������@� �� ����� �
��������� �  �� � �� �� ��6 G��6��� �  �� � �� �� ��L����6����Z���&  ?�4��������� �  !�L����  !�4��  ��4�� �4�6�0� ��4�-��& � �5�6L�� ��4��  �L���	  � �L���  � � ��6��� �6L���ɉ���������
	�� �9� � �* ���s��������@� �`�����P�M�N�0����� �� ��`�9�3� �#�9� �(�-��.���������i�# ��#��`�  I����I�%��`�E����`�� ���K`�4
�����-����.l-  �π�� �� � �����0���� ���0�0� ��`��6`H�H�H�6� �� ��� �� ��槥s� �h�h�h@���& ������ � � �* ���  !����[��� ����������& ��Ť���� �� K����쥣���楧i<ŧ��`���Ơ`栥��>�]�:��8� 8�i0���i ����������������i0�����i ����㥢���  ���a�.�]�*�D 8����ȑ���� ��i0��i ������� ���_��a�Ș s��a�����`�`���ơ`���K�]�G��8� 8�i��i ��i0���i ����������������i0�����i ����㥣��� ���a�0�]�,�D 8��ȱ����'��� ��i0��i ���ߩ�����a�����`�`



}�󅥽��i ���J��� 8��e��i �������`� � ��@�� ��������`H)��S�hJJJJ�
ei@}c�` 0`��� P���@p��      

�� ��� � �����`� �/ ���� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������!���