�<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���* 0 � � 0 0 0   0����  У���#  �#���#���#
��#���#��# ��#���#���#  �����WUU��������< �< �< �< �< ����   ��������� �< � ����   ������ �� �� ������   ������0����0������   �         ? ���� � � � � �? � � �       ?��    �?�   ��< �         < ���   <      �     ��    ��    ��   ����  �    ��   ���   s��   s��   ��   w��   � �   �  �   � ��   p����pT��r���<��  ��  ��[���[������������  ��  ��  ��  ��  ���������    ���������?������ ��  �<  �  �����    �����?������ �� �� �����?������    ����<�?��������?��������<�?�����    �����ꬪꬪꬪꬪ����   ����������  ������������������������������������    �kU�kU�k}�k}�kU�kU髪ꫪ���� �� � 3��0��   �� �� ����� �?��?� 0�� ?< �� ��  �� � 3��0��   � �  ����� �?��?� 0�� 0< << �? �?  ��  ?�3� 3�00��00��3�00�?����������?����       UUUU            ��  ��? ����� ��#�0� ��� ���( ���� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                    ������? ��� ���� ����               <0 <��   �                  �PUU�0U�S��TUU�SUULUU<           0TUU�3U�S��TUUSUU?LUUU�            @�3U�S��T@?SU  ?LUT�          �*��3����Ϩ*�*?����?����          �*���3����Ϩ*�*?����?����          �*���3����Ϩ*�*?�� �?����          ����3����Ϩ��*?���2 �����          �*� 0����Ϩ��*?�������*�          0 �0��������?�������          �?�?�0���������?���������            ������������?�������?           ��?���������?��?�� <��?�             ��������?���������3��          ������������?������������          ���?�����?�? ����������             �? ���  �    � ��          ������������?  ����������          ����� ���� ��?  ����������          ����? ��� ��?  ���������                                                                                                                                                                          ��� ��   ��?  ���  ����           �   �  <    �  <  �  ?�          �TUU�SU�  �PU U0�T�          �TUU�SU�  0TU<�PUU��TC�          �T@�SU�  0UUU��TUU��TS�          ��*�����  � ��0�*��Ϩ*��          ��*�����  ��<��3�*�Ϩ���          ��*�����  ��<��3�*��Ϩ���          ��������  �� ��3�*��Ϩ�*�          ��������  �����3�*��Ϩ�*�           ��������������3�?� ���?�           ��?���< <�����3�?�����?�           ��?�?�� �������3�?������          ��?�??���������3�?����?��          ��?�??�����0�����������?�?          ����?�����0��?��������???          �����?���������������??<?          �   �?   �� �� ?  ��  � ?          �����?����� ���� �������?�?           ��������� ���? ���� ��?�?           ��������� ��� ��� ��?�?                                                                                                                   ?  �     �?   ?�  ��  0<  �  �   �    ��   <  0  �   �     �       �?  �?    ?     ��   �  ��   �    <      �  ��   ��  0<     0�  ����  ��  �     �?  �?  ��
�
�
�                                                    <<<<<<<<<<<<<<<<<<<<<<<<                          0                �0    3   *>2  p��  �"k  �'H  �P�  �� 0oe�?  ��+  ���  ���?  0��<  ��  �     �          �    � 0�   @V� C̠�  �̨ �4��gP7�KT �RUU � ��������< P��:@�?�kP�;o:1@<<��  �?���P	0 �    �  0����  � ��00�����  �  �����         �                          �300 0���� �?��� �?����������000� ���0030 ����  � ���� 0�<03��0030 ����  � 0��� 003�3���?� �?��  <�?0���<�?003��� 0  ����  �� � ���� 000�0�00�  ����  � 0 ��� 000  �����? �?���  ��0�?��ppp p pxxxxx��� � ���� � ���� � �� f f 
f f fp	p	
p	p pzz
zz z
�
�

�
� �	��
�� �*
***44
4>>H� f f 
f f fpp
pp p	zz
zz z
��
�� ���
�� �*
***44
4>>H� f f 
f f fpp
pp p
z
z

zz z��
�� �
��

�� �*
***44
4>>H� f f 
f f fpp
pp pzz
zz z��
�� �	�
�
�� �*
***44
4>>H� f f 
f f fp	p

pp p	z
z
zz z	�
�
�� �	�
�
�� �*
***44
4>>H� f f 
f f f
p
p	
p	p pzz

z
z z
��
�� ��	�

�� �*
***z44>f� f f 
f f fp	p	
p
p p
zz
z
z z
�
�

�	� ���
�
� �*
***44
4>>H� f f 
f f f	p	p
pp p
z	z	
z
z z
�
�
�� ��
�	
�	� �*
***44
4>>H� f f 
f f f
p
p	
pp pz
z
z
z z
��	
�� �	��

�� �*
***44
4>>H� f f 
f f fpp

pp pz	z	
zz z
��
�� ��	�

�� �*
***44
4>H� f f 
f f fpp
p
p pzz
z	z z�
�	
�	� �
��
�� �*
***44>>H�� f f 
f f f	p	p

p	p p	z
z
z	z z	�
�
�	� �
��	
�
� �*
***44
4>H� f f 
f f fpp
pp p
z
z
z
z z
��
�	� �
�
�

�
� �*
***44>>H�� f f 
f f fpp

p	p p
zz

zz z
��	
�� �	��
�
� �*
***44
4>>H� f f 
f f f
p	p

p	p p	z	z	
z	z z
��
�� ��	�
�� �*
***44
4>H� f f 
f f f	pp
p
p pzz

zz z�	�
�� �
�
�	
�	� �*
***44
4>>H� f f 
f f fp
p

pp pzz	
z
z z
��	
�� �	�
�
�
� �*
***44
4>>H� f f 
f f fp
p
pp p
z
z

z
z z	��
�	� �	��
�	� �*
***44
4>>H� f f 
f f fpp
pp pz
z
zz z�
�	
�	� ��
�

�� �*
***44
4>>H� f f 
f f fpp
p	p p	zz
zz z
�
�
�
� �	��

�� �*
***44
4>>H� f f 
f f f
pp	
pp p	zz
zz z�
�	
�
� �	��

�� �*
***44
4>H� f f 
f f fp	p	
pp pzz
zz z
�	�
�
� ��
�

�	� �*
***44
4>>H� f f 
f f fpp	
p
p p	zz
z	z z
��	
�� �
�	�
�	� �*
***44
4>>H� f f 
f f fp
p
pp pzz

z	z z��
�	� �	�	�

�
� �*
***44
4>>H� f f 
f f fpp
p	p p	z	z
z	z z
�	�
�
� �	�	�
�	� �*
***44
4>>H�ff
fffpp
p
ppzz	
z
zz
��

���
��
���*
***44
4>H�ff
fffp
p	
pppzz
zzz��
�����
���*
***44
4>>H�
ff	
f	f	f
pp
ppp
zz
zzz
��
���
�	�
���*
***44
4>H�
f
f

f
f
f
p
p

pp
p
zz

z
z	z
��
�
�
�	�
�

�
�
�*
***44>>H��ff

fffpp
p
pp
zz
zz
z	�	�	
��	�
�	�
���*
***44
4>>H�
ff
f	ff
p	p
pp	p
zz
zzz
�	�	
���
�
�
��	�*
***44
4>>H�f
f

ff	fp	p
pp	pz
z
zzz�
�

�
�
�	�
�	
���*
***44
4>>H�ff
f
ffpp
pp	p
z
z
z
z	z	��
��
�
�	�	
��
�*
***44
4>H�f
f	
f
ff	pp

p	p
p
z
z
zz
z��
��
��	�
���*
***44
4>>H�f
f

f
ffp
p
p
p
p	z
z	
zz
z
��
��
�	�
�
��
�*
***44
4>H�ff

f	f
f
p
p

p
p
p	zz
z
z	z	�	�	
�	�	�
�	�
��
�*
***44
4>>H�f	f
f
ffpp

pp
p	z	z

z
zz
��	
�	��
�
�
��
�*
***44
4>>H�ff	
ff
f	p
p
p	pp	zz

zzz��
���	�	�	
�
�
�*
***44
4>>H�	f	f

fff	p	p

p	p	pzz

z	zz��

�	��	��

�	��*
***44
4>H�
ff

ff	f	pp
pp	pzz

z
zz	�	�	
�
���
�
�
��*
***44>>H��  .  2  N  R  V . 2 N R V  .  2  N  R  V 0. 02 0N 0R 0V @. @2 @N @R @V P. P2 PN PR PV `. `2 `N `R `V p. p2 pN pR pV �. �2 �N �R �V �. �2 �N �R �V�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ���ة��8���  ��� � �?� � �@� �ߍ& ��" � t ���d%��&�� � �%����&��� ��X��>�#  I� o� �� ^� ~� ��	���P�� �� A� �� )� �� �� U� �� ���<� �� �� O� iĩ�<�:� ��d:�;�� �� �� �� Ué�;L�����F�	� F���F�	���i +�آ  7�����`�x���<�������y0, N����i��إ�i���(� )�� ���� ��LX� ^�Ls� �� a�`���A�	� F���P�	� F�  7���<��` �ȥK������	����
�� � �� �ȩ��D����E������ � �ȩ�� Q�E8��E�	 �� K�E�d�� �ȩ�� Q�Ei�E�	 �� K�EɈ�� 7� 7� 7� 7� �ȩ�� Q�E8��E�	 �� K�E�d�� �ȩ�� Q�Ei�E�	 �� K�EɈ�� 7� 7� 7� 7� 7� �ȩ�� Q�E8��E�	 �� K�E�d�� �ȩ�� Q�Ei�E�	 �� K�EɈ��` ک ������P�� �Ѭ   ;ۘ	�����	����� � ^�Ls� ^� ��LX��	�����	�����	�����	�����	�ɿд��i����� �� �ѥ�i���x��P�� ��Ls� �ȥK������	����
�� � �� �ȩ�� Q���"����	������ � �ک��A�	� F�
��P�	� F�  7���(��`L ĥK��� �x`��1�f�2� �x�1�9���2�2� �K��� ��2i
�2ɘ�� �إ1i�1 ĥ1���f�2� ����л��1���2� ���2�5�x�1�.� �K�2� ��18��1�0� �إ28�
�2 Nĥ2�\�	� ����п���x�� �x`ڥ1�
���x��	���>����#��1i�1����x�
�	���4����#��1i�1�`ڢ���2�	�28�
�2���#���`` �ȥEi�f��F���G�Ei�P(�� � ��Ei�0���0��x�F0i�F��#�ڢ � � ��x�F����G0�8�
�G���ߥF��G�	������
�� � ��`��� � � ��x����	�
� _�����`� �%�y� � �	�y�8��y����� �{� � � ��{i�{����z8�{�0� �.�{�z���1�08��� �
�1e1�1ʀ� �ť}e1�}�~i �~�`�0�0�
��P�	�1 +���P�	�  +�2�:`�����
��P�	 _�`����	�y +����	�~ +����	�} +�"���	�| +�`��� � ƀ�� �� � ��`� �1� �[���<�S�x�5�K��� � � �ǥS��J� �؅K� ���1 � �ǥS��/� ����иL�ƽ � � �ǥS��� ���1�� ��L��L�Ƣ �x��(�[���!Ɏ�"�K� �	 � ��L�ƽ � �� ��L�����̥K��� � � ��L|ƅK� � ȩ�1 ��L|ƽ � �	 � ��L|ƥ1�� �� ��`� �1�[Ɏ�d� �S�x�9�[���2�K��� � � �Ǣ �օK� ���� Q��1 �ǩ � � ����лL�ǽ � � �Ǣ ���1��> ��L�Ǣ ��Ɏ�*�S�x�#�K� �� � L�ǽ � ���1��
 �ǀ���� ��`��� Q����K�0� �K�0� ��S�Ei�[ ��`��� Q� �� �ĩ����S�Ei�[`�  �ȥS8��S � 7�����`�  �ȥ[i�[ � K���
��`��� Q�x�
���� � �\��� �x�
����	��i
������`���D��E�	������� ��`���F�	� F�`�
������F�	 _�`�H���
��S��[�	 _�h�`�H���
��x����	 _�h�`�����D��E�	 _�`���
��F��G�	 _�`�  ��� ;�LX��	����/���� ���[i
�[Ɏ����[�Ei
�EɈL�ɩ��EL�ɘ	����/���� ��8�[�
�[�*0��*�[8�E�
�E�$0L�ɩ$�EL�ɘ	�����S��� ��L�ɘ	�� ��`H {� m�x� �  T� ;� 7�  ��� ;� {�Xh`�K� �f� �Ȧ��0�eS�S� 6ʥS�� �ȩ���[Ɏ����3�e[�[�	8�d�*0���� �ȩ����S�Ei�[ �ȩ���
�� � ��`����
��S��[�	� � ��`�    ��[����S8��x�������#��`��
����ȹ��� � ����� ȱ�xȱ���Ȁ�dz� � � ��zi�z����`����
�� �� � � ���x����	 ����#��` ���d	������� �������$0��� �	 �������$0�����	 �������$0�dd	����� ���	i�	ɠ��&�d	 ���	i�	ɠ�� ��(�	 ���	i�	ɘ�����	 �ک���	 �ک���	 �ک���	 �ک���	 �ک���	 �ک��
�	� F����	������ +���
�	� F����	�y +����	� F�`���E�"�D���[��S��F�R�Gd<d;d:d���������K� �Uâ � �x����#��`� �� #�`��� #�`��� #�`�   ;ۘ	�����	���� �d�d�d|d}d~Ls���L��L<Ԙ	����#�i��� � �ѥ�iɌ��P�� ��LA̘	���О�8������ �ѥ�8��<��x�� ��LA�` �� 9� 3ک ������P�� �� �� �� �� �� ե;��$�$�� W�d$������; �� >� (Υ<�  � �� �� }�  � � �ة�<�9к <� (Ω�9��`�=���������� )� ��d= �� ک ������P�� �Ѭ   ;ۘ	�����	��"��� � ^ڥ��L����LW� ^� ��LX��	�����	�����	�����	�����	�ɿЧ��i����� �� �ѥ�i���x��P�� ��Li� �ѩ��B��C�	������ � �� F� M������� �� F� M����� ��`� �K � �c� � � �U�x�S �M��� 0Fi�[ �>� �J�x�0���1ڢ � � ��J� �0�x�1i��� �K  �΀��x���L����xП��Б`�Z�J��d �0� �1� � �J�	���2� ���x�� � �J����20��1��2��1��x��1�0���� Q� 3�Z���� ��0 z�zz�`���B��C�	������� ��`���F��G�	������ � ��`������ �� �K� �%�� w�8�[��[� �� �K����S��[�	 ������`dG� � � ���� 0�x�F����G0��i�G��x���G`�  ��� ;�LX��!�!�0&d!�	�����Bi�Bi�F�`��Bi�FLS�� � �0&d �	����8�B��Bi�F��`��Bi�FLS����0*d�	����!� �K� ��c�K�Bi�S���[�����LSЊ	�� �� W�`����  m�mm"e}e<e;e9)�0 ���  m�mm"e}e<e;e9)�0�
�����ȹ����� ����.�d� ���)��������dȱ�Hȱ�*�+ȱ�, �����`�Z�H
����'ȹ��(� �'��� 
ѥ+�*�,i�,Ȁ�z�`�Z� � �1�1
�1�!� � ��)� �*�x�,���	��x�� �����	�*i�*��z�`��d	����� _�`�����x����	� 0 _�`�����S ��[ �	 _�`�����B��C�	 _�`�����F��G�	 _�`����������	 _�`������ ���������	 ��`�:�G���J� � �J� ]���x�� � �J�����ɀ�	 3ҩ��=� T���x�����å�����:`ڢ � �J� ]ѩ � ��x��J�� �d �`ک����� ����x����	� 0 ���`�Z��}e0�}�~i �~ة$���	�| +�"���	�} +����	�~ +����*�� ��z�`� �������� �� ��5�����5��ȹ5��	ȹ5�� ��Ȁ�
�������	 _�
������@�	 _����	� F�$���	�  +�"���	�  +����	�  +����*�� �ة��D�	� F�@���Z�� �ة!��P�	��i +�`��F� �G���C��B  ϩ�c� �G� tK����� � �x����x���$� �=��8�<�;�:�9�}�~`�   ;ۘ	�����	��L�̘	����#��i��� �� �ѥ�i� ���� ��L�Ә	���и��8������� �ѥ�8������ ��L��` �� 1� 3ک ������P�� �� �� �� m� �� �ԥ;� ֥�����; r� >� pե<�  � � n� M� &�  � � �� �ة�<�9о �� pթ�9�����Z�0�~�00P����:�0�~� 0@����*�0�~�00�����0�~�0 ����
�~�0����!��P�	��i +�`���Z�0�~�00P����:�0�~� 0@����*�0�~�00�����0�~�0 ����
�~�0����!��P�	��i +�`� �K � �� � � �q�x�S �i�[ 8����^� �K �%��� Q�Z������0 z�z� � �K  B� X�L�թ�� Q� �ڢ � � ��I� �0�x�1i�����P���L����PЃ���Lr�`� �K � �I�x�0���1`�  eCeBeee;e:)�0�i�I�  eBeCeeee;e:)�0�����0� � � ��I� �0�x� ��Lq���P��`�:��� � � � B�����ɀ�� � ���=� ����P�٥�����:`������ �� ��x����	 ��`���F��G�	������ � ��`������ �� �K� �#�K��S��[�	 ��8�[��[� �	� �K�� X�����`dG� � � ��x�F����G0��i�G��P��`�  ��� ;�LX��!�!�0&d!�	�����Bi�Bi�F�`��Bi�FL�� � �0&d �	����8�B��Bi�F�0`��Bi�FL����0d�	�����	�����c�c��Cdc�cL����0*d�	����!� �K� ��c�K�Bi�S���[�����L؊	�� �� W�`�c��Bi��Ci�	������� ��`�����x����	 _�`�����S ��[ �	 _�`�����F��G�	 _�`�������� ������	 ��`�x���� i�`� �������� �� ��5�����5��ȹ5��	ȹ5�� ��Ȁ�
�������	 _�
������@�	 _����	� F�$���	�  +�"���	�  +����	�  +����*�� �ة��D�	� F�@���Z�� �ة!��P�	��i +�`��F� �G���C��B  ϩ�c ة �G� tK����� �=��8�<�;�:�9�}�~`�   ;ۘ	�����	��LWԘ	����#��i��� �� �ѥ�i� ���� ��L�٘	���и��8������� �ѥ�8������ ��L��` ����P�	�
 F���d�	� F�`���<�	� F�������� ��
��P�	 ��`� � � ��x��� � �d����� � �K����dHdIdJdcdy� �x`H�Z�
��h���h���� ��e��i ����e��i �� ��@��	� ��i0��i ����e��i �� � ڱ�� ���1�
���Q����������i0��i ��e��i ���z�h`H�  ����h`Hd8�  ����8�(0�h`H�  �������h`H�Z��ŉ���ŋ���������L�ۥ�������L�ۥ�ŉ���������L�ۥ�������接�Ŏ�LE�)� ����L�������L�����0��L�ۢ���������D���JJ�����L��接�Ŏ�LEܥ�)� ����L)������L)����0��L)ܢ���������D���JJ�����L��z�h`� ������ !� %�� � � � � � � � �* d�d�� ����d�`�������� !ॵ� ���  {�漥�ŷ� �ݥ������� %� �Í  ���ɥ���� �ݥ����J�������� !ख़� ���  �ޥ������� %१� ���  (�栥�ś� '�殥�ũ� Dޥ���� )� ��`������ȱ���ȱ���ȱ���ȱ���)
��W셞�W셟��)0��ȱ������Ȅ�d�d���� �L�ݤ� ��� �
��� �d���Ȅ�d���������ȱ���ȱ���ȱ���ȱ���)
��W셺�W셻��)0��ȱ������Ȅ�d�d���� �� ��� ��)��	����d� ��`������ȱ���ȱ���ȱ���ȱ���)
��W���W�ȥ�)0��ȱ������Ȅ�d�dʥ�� к� ��� ��)��@Ы����d� �݀�������ȱ���ȱ���ȱ���ȱ���)
��W셬�W셭��)0��ȱ������Ȅ�d�d���� й�� ��� �
��� �d���Ȅ�d�����
��������ݱ܅�ȱ܅�`��
������ݱ܅�ȱ܅�`H�Z��)?	@�̤�;��%̤̅������)@��J��̥̅��8������)0��Ȅ������ơ��d��̍ z�h`H�Z��)?	@�̤�;��%̤̅������)@��J��̥̅��8������)0��Ȅ������Ư��d��̍ z�h`H�Z��)?	@�̤�;��%̤̅������)@��J��̥̅��8������)0��Ȅ������ƽ��d��̍ z�h`H�Z��)?	@�̤�;��%̤̅ʱǪ��)@��J��̥̅��8��ˀ��)0��Ȅʱ�����ʥ�dʥ̍ z�h`� `� `H�Z������ک��م��)?
��i���i��d� \�z�h`d��* d�`����ȱ��ȱ��ȱ��)
��W���W�ҥ�)0��Ȅ�d�dӥ�� T�d�`H�Z�����L�΅ץ�;��)��פӱѪ��)@��J��ׅץ��8��ր��)0��Ȅӱ�����ӥ�dӥ�)�̥�)����
�@����̥̅׍( ������* ���Х���� \�z�h`H�Z�  �ޠ  ��d�d������ '� D� �� (� )����z�h`H�Z��� ���� �dߥ�)?�ߐD�� �>��
��3셳�E���3셴�E��d�d�� ������)������ �ݥ����� �� )�z�h` �� � �
� � �
� � �
� � �
� � 
� � �
� � �� � �� � �� � 
� � 8
� � ?
� � 8
� � ?
� � K
� � _
� � T
� � K
� � G
� � ?� � K� � ?
� � � �     � �� � �
� � �
� � �
� � �
� � 
� � �
� � �� � �� ��� � 
� � 2
� � _
� � T
� � K
� � G
� � ?
� � 8
� � 2
� � /
� � *� � ?� � ?
� � � �     � q
� � d
� � _
� � T
� � K� � � � T� � � � �(� � �
� � 
� � q
� � d
� � _
� � T
� � K
� � G
� � ?� � T
� � K
� � _� � � � ?
� � G
� � K
� � T
� � _(� �     �.� \� �.�  \� �     � �� � �� � �
� � �
� � �� � �� � �� � �
� � �� � �� � �� � q� � � � �� � _<� � _� � T� � j
� � j� � T� � _� � q
� � q� � q� � j� � �
� � �� � �� � _<� � _� � T� � j
� �     � j� � T� � _� � q
� � q� � q� � j� � �
� � �� � �� � �P� � Gx� � Kx� � T� � j
� � j� � j� � j(� � K� � T� � _� �     � q
� � q� � q� � q(� � _� � T� � _� � j
� � j� � j� � j(� � _� � T� � _� � q
� � q� � q� � qP� � Gx� � Kx� � T� � j
� �     � j� � j� � j(� � K� � T� � _� � q
� � q� � q� � q(� � _� � T� � _(� � j(� � q(� � (� � �(� � _� � q� � �<� �     ��� �:�  :
� �:
� �:� ��� �:� :
� �:� ��� �:�  �� ��� �:� �}<� }� �T�  �
� ��� �T� �}� �
� ��� ��� ��� \
� �\� �\� �}<�  }� �T�  �
� �     ��� �T� �}� �
� ��� ��� ���  \
� �\� �\� �:P� x� .x� T�  �
� ��� ��� ��(� .� �T� �}�       ��
� ��� ��� ��(� }� �T� �}� �
� ��� ��� ��(�  }� �T� �}�  �
� ��� ��� ��P� x� .x� T� �
� �     ��� ��� ��(�  .� �T� �}�  �
� ��� ��� ��(� }� �T� �}(� �(� ��(�  �(� �:(�  }� ��� �:<�      � ��� ?��}�� _��}�� ��� (�� ��� ?�� ��� ?
�� q
�� ?�� ��� _(�� ��� K�� �� 8�� �� G�� (�� ��� ?�� ��� _
��}
�� _�� ?�� �(�� ����� ��� ��� �(��     � �� �� ��� /�� ��� K�� ?(�� �� �� G�� 
�� 8
�� �� K�� /(�� _�� %�� ?�� �� ?�� #�� ?(�� �� �� K�� /
�� �
�� /�� �� (�� ?�� ��� _�� K�� _(��     ��(�\(���(��(��\(��(��     �}(�.(��}(� �(��.(�}(��     � �
�� /d��     � ���     � ���     � ���� ��� _��� K��� ?��� /���     � _��� _��� ���     � ��� _��� K��� ?��� /��� %���     � ?��� C��� G��� K��� T��� _���     � ?��� /��� %��� ��� ��� ���     � ���� G��� *��� ��� ?��� ���     � ���� ���� ���� ���� ����     �
	��
�
�
	�
	�
	 �

		�
	���'���-��H���  ��  ��j���x�  ���@���  H� �  ��"�  j�j�j�j�j�j�j�j�L�^�v������6�`�L������������s����?� $  o  $ � �� � ��      D   D   D   D      D   D   D   D   D   D   D   D   D   D   D   D      O   O      �    �:    ک2�;�`�Z�;� �� ���z�`�Z�:� �� ���z�` �� 7��� ��`����	���%���2�� � �ک��P�	� F���d�	� F���x�	�	 F�����	���!����� � ��`H�Z���7� ������� �
�����	�
� ���r� ����d�������	�
�� ���� ������	������� ���D� �L� � ��	���
�� �� �
i�
� ������ �8��� ���T� �La� �� (ߩ��� Q�z�h`xH�Z��
��3�%�3�	�)��&��0��1�	���-�D�.�JJ��%%7�-�%i�%�&i �&�1�1� �Ȁ��0�0� ���1�L��z�hX`H� �7 ����7h`H�Z�/���� ���� ��z�h`����Z�P���� ���� ��z�`�Z�%���� ���� ��z�`H�Z�	���e��D�i �� � ���0�����z�h`H�Zd%�@�&� � � �%����&���z�h`
	
	
	


	


	
������
		xndF2(
		
Ò-����k�Ք<����z��K�������W���+�����f�Л:����u�ߝF�������U���&�����d�ˢ����؂���r�Z���N�
�2�Z�����N�҄��΅�����W�ϐG�0�7�o������������������*�7�H�U�f�{�	�	�	������������	��	��	���������� ��	��������	���	����	
��������
������������������������������������@@@@�� ������@�����	xH�Z�/�a��$��b��%��c��&��d��'��J�%�r�&��0�	���-�D�.��%�-�%Ȳ%�-�%��0�0����z�hX`H�Z�)�JJJJ�/ ��)�/ ��z�h`H�Z
��$�5�$�6� �5�$��a�8�7�/ ��Ȁ�z�h` GAME  OVER $PAUSE$LEVEL  :$HEIGHT :$CLEAR$BLOCK$SCORE$aaPLAYaBLOCK$aaFILLaBLOCK$aaaHITaBLOCK$CONTINUE$END$AaBaCaDaEaF$STAGE$SORRY$aaaYOUaFAIL$SELECTaDIFFICULTY$HERRO$aaaYOUaPASS$q�~���������������������� ���  0@P`p��������  0@P`p��������  0@P`p���������������������������������������� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____H�Z�8�<��<�;��;�:��:�9��9(z�h@H�Z����� �� �ܭ' )��8�>�# �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �� ��