UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUU���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUZUUUUUUUZUUUUUUUjUUUUUUUjUUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�VUUUUUU�VUUUUUU�ZUUUUUU�ZUUUUUU�jUUUUUU�jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUU  PUUUU   UUUU   UUUU    UUU ��?UUU ���UU ����UU �*��UU �> �UU ��� UU  Z� UU   �TU      �      ���     �����   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU UUUUUUU  @UUUUU   @UUUU    TUUU�?  VUUU�� �VUUU� �VUUU� �VUUU� ��VUUU ��VUUU ��VUUU ���VUUU ���VUUU ���VUUU���VUUUUUUUU���UUUUU���UUUUU���UUUUU�j�UUUU��j�UUUU��Z�UUUU��V�UUUU��U�UUUU��U�UUUU��U�UUUU��V�UUUU��V�UUUU��Z�UUUU��Z�UUUU��Z�UUUU��j�UUUU��j�UUUU����UUUU����UUUU����UUUU����UUUU����UUUU����UUUU����UUUU����UUUU����UUUU����UUUU�����jUUUUUU��UUUUUU��UUUUUU��VUUUUU��VUUUUU��VUUUUU��ZUUUUU��ZUUUUU��ZUUUUU��jUUUUU��jUUUUU���UUUUU���UUUUU���VUUUU���VUUUU���ZUUUU���ZUUUU?��ZUUUU?��jUUUU?��jUUUU?���UUUU?�UUUU?�VUUU?���VUUU?���VUUU?@��ZUUU?@��ZUUU?@��jUUU������ ��������U�������U�������U�������U�������U�� ����U�� UU��U�� UU��U��UU��U��TU��U��TU��UU�PU��UU�?PU��UU�?@U��UU�?@U��UU��@U��UU�� U��UU��U��UU��T��UU��T��UUU�P��UUU�P��UUU�?P��UUU�?@��UUU��@��UUU�� ��UUU��������VUUU����VUUU�Z��VUUU�V��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUUjU��VUUU*U��VUUU*U��VUUU*U��VUUU*U��VUUU*T��VUUU*T��VUUU*T��VUUU*P��VUUU*P��VUUU*P��VUUU*@��VUUU�@��VUUU�@��VUUUUUUU����UUUU����UUUU����UUUU����UUUU�O��UUUU�O��UUUU���UUUU���UUUU���UUUU���UUUU���UUUU���UUUU���UUUU���UUUU�P�UUUU�P�UUUU�P�UUUU�P�UUUU�P�UUUU�P�UUUU�P�UUUU�P�UUUU�P�UUUU��UUUU� �UUUU� �UUUU� �UUUU� �?@��jUUU>@��jUUU>@���UUU:@���UUU:@տ�VUU*@���VUU*@U��ZUU*@U��ZUU�@U��ZUU�@U��jUU�BU��jUU�BU���UU�JU���UU�JUտ�UU�JU���VU�jUU��VU�jUU��ZU��UU��ZU��UU��jU��UU��jU�� �jU�� ���U��
 ���U��
 ���V����? �V����? �Z������Z������VUUU����UUU����UUU���UUUU��UUUU�?�UUUU�?�UUUU���UUUU���UUUU���UUUU���UUUU����UUUU����UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��� ��VUUU���VUUU���VUUU���VUUU���VUUU���VUUU���VUUU�?��VUUU�?��VUUU�?��VUUU����VUUUj���VUUUj���VUUUj���VUUUj���VUUUj���VUUUj���VUUUj���VUUUj���VUUUj���VUUUj���VUUUjU��VUUUjU��VUUUjU��VUUUj�VUUUj �VUUUj ��VUUU* ��VUUUUUUU� �UUUU� �UUUU���UUUU��jUUUU�  UUUU�  UUUU�  UUUU�  UUUU����UUUU����UUUU����UUUU����UUUU����UUUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���U ��U��� �jU�����ZU���
��VU���
��UU@��*�jUU ����ZUU ����VUU�����UUU����jUUU����ZUUU����VUUU����UUUU���oUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUտUUUUUUտUUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU* �jUUUU*��ZUUUU*��VUUUU*��UUUUU��ZUUUUU��VUUUUU�jUUUUUU�ZUUUUUU�VUUUUUUjUUUUUUUZUUUUUUUVUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUZUUUUUU�ZUUUUU��ZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU UUUUUU  UUUUU   UUUU  �UUU   �UU   ��UU  ���UU?  ���UU�  Z�UU�?  @�UU��  �UU���   UU���  UU���� UU� ��? UU� ���UU� U���UU� U���UU� UU��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUU@UUUUUU  TUUUUU  @UUUUU   TUUUU�  UUUU��  PUUU��  UUU��� PUU
���  UU��  TUT=  �UU  ��UU   �jUU   ��jUU  ���jUU ����ZUU ����ZUU�����ZUU��j��VUU��U��VUU�VU��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUU��ZUUUU���ZUUU����ZUU�����ZU������ZU�����ZU����իZU���VիZի�ZU��ZիjUU��ZիZUU��Z��ZUU��Z��ZUU��Z��ZUU��Z��ZUU��Z��ZUU��Z��ZU���Z��ZU���Z��ZU���Z��ZU���Z��ZU���Z��ZU���Z��ZU���Z��ZU���Z��ZU���Z��ZU?��Z��Z�?��Z��Z�?��ZUU� UU��UU� UU��UU� UU��UU� UU��UU� UU��UU� UU��UU� U���UU� U���UU� U���UU� U���UU� U���UU� U���UU� U���UU� U���UU� U���UU� U���UU� ����UU� ����UU� ����UU� ����UU� ��j�UU� ��j�UU� ��j�UU� ��Z�UU� ��Z�UU� ��V�UU����V�UU����V��TU��UUU�TU��UUU
TU�jUUU
TտjUUU
TկjUUUTկZUUUT��ZUUUT��VUUUT��VUUUT��VUUUT��UUUUT��UUUUT��UUUUT�jUUUUԯjUUUUԯZUUUUԯZUUUU��ZUUUU��VUUUU��VUUUU��UUUUU��UUUUU��UUUUU�jUUUUU�jUUUUU�jUUUUUïZUUUUUïZUUUUUUUUUUUU�UUUUUUU�UUUUUUU�UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU�?UUUUUU�?UUUUUU�UUUUUU�UUUUUU�UUUUUU�UUUUU��UUUUU��UUUUU�� UUUUU�� UUUUU�?@UUUUU�?@UUUUU�?@UUUUU�UUUUU� UUUUU� UUUUU� UUUU�� UUUU�� �UUUU�� ���Z���Z��Z���Z��Z���Z��Z���Z��Z���Z��Z� ��Z��Z� ��Z��Z?@��Z���?@��Z���?P��Z���P��Z���P��Z���T��Z���T��Z���T��Z���U��Z��� U��Z���@U��Z��:@U��Z��: U��Z��
 T��Z��� P��Z���@��Z��� ��Z���? ��Z���� ��Z������Z��Z���ZUU��U�UU��U�UU��jU�UU���jU�UU���jU�UU���ZU�UU���ZU�UU���VU�UU���VU�UU���VU�UU���UU�UU���UU�UU��jUU�UU��jUU�UU��jUU�UU��ZU�UU��Z �UU��V��UU�����UU�����UU�����VUU����jUUU����UUUU���ZUUUU��jUUUUU��UUUUUU�VUUUUUUZUUUUU�VUUUUU�VUUUUU�VUUUUU��UUUUUU��UUUUUU�jUUUUUU�jUUUUUU�jUUUUUU�ZUUUUUU�ZUUUUUU�VUUUUUU�VUUUUUU�VUUUUUU�UUUUUUU�UUUUUUU�UUUUUUUjUUUUUUUjUUUUUUUZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�? �UUUU�? �UUUU�� hUUUU��@UUUUU� UUUUU�? UUUUU�� UUUUU��UUUUUU�UUUUUU�?UUUUUU��UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��Z�?��Z��Z����Z��Z����Z��ZU?�Z��ZU��Z��Z  �Z��Z   �Z��
  ��Z��
  ��Z��
 ���Z��
����U��
���ZU�����jUU�����UUU����ZUUU����UUUU���VUUUUիjUUUUUU�VUUUUUU]UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�������_�������[�������[�������[�������[�������[�WUUU��[��UUU��[��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��ZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   UUUUU   UUUU   UUUU   UUUU   UUUU ���UUUU ���UUU ���UUU ���UUU �ZUUUU ��ZUUU ��ZUUU ��VUUU     UU     UU      U      U�������U�������U�������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU    XUUU    XUUU    ZUUU    ZUUU   �ZUUU���ZUUU�� �VUUU�? �VUUU���VUUUU��VUUUU��VUUUU ��VUUU ��UUUU ���UUUU ���UUUU ��UUUU ���UUUU����UUUU���jUUUU���jUUUUUUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUUU�UUUUUU��UUUUUU��UUUUUU��UUUUUUտUUUUUUտUUUUUUտUUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU����UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UUU��Z��UU���Z��UU���Z�UU���Z�UU���Z�UU���Z�UU���Z�UUտ�Z�UU���Z��UU���Z��UU���Z��UU���Z��UU���ZU�������U�������U��Z��U�U��Z��U�U��Z��U�U��Z��U�U��Z�jU�U��Z�jU�U��Z�jU�U��Z�jU�U��Z�jU�U��ڿjU�U��ڿjU�U��ڿZU�U��ڿZU�U��گZU�U��گZU�U��گZU�U��گZU�U��گZU�U����VU�U����VU�U����VU�U����VU�U����VU�U����VU�U����UU�U����UU����jUUUU��jUUUU��jUUUU��jUUUU��ZUUUU��ZUUUU��ZUUUU��ZUUUU��ZUUUU��ZUUUU��VUUUU��VUUUU��VUUUU��VUUUU��VUUUU��VUUUU��UUUUU��UUUUU��UUUUU��UUUUU��UUUUU��UUUUU��jUUUUU��jUUUUU��jUUUUU��jUUUUU��jUUUUU��jUUUUUUUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUU���UUUUU���UUUUU���UUUUU���UUUUUտ�UUUUUտ�UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUU���UUUUU��
UUUUU��
UUUUU����UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��UU���Z��U���Z��U���Z��Uտ�Z��Uտ�Z��Uտ�Z��UտگZ��UտگZ��U��گZ��U��گZ�
 ��گZ� ��֯Z�  ���Z �����Z������Z������ZU����UU�U����UU�U����UU�U����UU�U����UU�U���jUU�U���jUU�U���jUU�U���jUU�U���jUU�U���jUU�U���jUU�U���ZUU�U���ZUU�U���ZUU�U���ZUU�U���ZUU�U���ZUU�U���ZUU�U���VUU�U���VUU�U���VUU�U���VUU�U���VUU�U���UUU�U���UUU�U���UUU�U���UUU���ZUUUUU��ZUUUUU��ZUUUUU��ZUUUUU��ZUUUUU��ZUUUUU��VUUUUU��VUUUUU��VUUUUU��VUUUUU��VUUUUU��VUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU��UUUUUU�jUUUUUU�jUUUUUU�jUUUUUU�jUUUUUU�jUUUUUU�jUUUUUU�ZUUUUUU�ZUUUUUU�ZUUUUUU�ZUUUUUUUUUUU��UUUUU��UUUUU���UUUUU���UUUUU�+�UUUUU���UUUUU�
 UUUUU� UUUU��  UUUU��  UUUU����UUUU����UUUU����UUUU����UUUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����� �V�������U�UU���jUjUU���ZUZUU���VUVUU���UU  @��jUU  @��ZUU  @��VUU  ���UUU����jUUU����ZUUU����VUUU����UUUU���oUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��jUUU�U��
   �U��   �U��    �U�?    �U�������U�������U�������U�������U�������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�ZUUUUUU�ZUUUUUU�VUUUUUU�VUUUUUU�VUUUUUU�VUUUUUU�VUUUUUU�VUUUUUU�UUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?    0<<?�?�<<0  ���?    �?��    �������?���?<  <<  <�  �����?� ��  �?  �  �      �  �  �  �  �  � ���������������� �  �  �  �  �  �   0 < ����< 0         ����      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                UUUU���  p  p��p��p��p��p��p��p��p��p  p  p���UUUU��������WUUUUUUէ�UUUU�ڧ�uUUu�ڧU�UU]UڧUUWUWUڧU�]�]UڧUUwuWUڧUU��UUڧUUuuUUڧUU��UUڧUUuuUUڧ�U�_U�ڧ�UUUU��WUUUUUU�����������������WUUUUUUէ�UUUU�ڧ�U�WU�ڧUU]]UUڧUU�wUUڧUU]]UUڧUU�wUUڧU�]�UUڧUuWuWUڧU�U�UUڧUuUUWUڧ�]UU]�ڧ�UUUU��WUUUUUU�������������WUUէ��ڧ��ڧUUڧUU�WUU��UU�WWU�W�U�Wuw�W���WUw�WUw�WUw�W���Wuw�W�U�WwU��UU�WUU�WUUէUUڧUUڧ��ڧ���WUU���������WUUէ��ڧ��ڧUUڧUU�WUU�WUU�WUU�WU��WUw�W�]�WwW���U���U���U�WwW�W�]�WUw�WU��WUU�WUUէUUڧUUڧ��ڧ���WUU�������������  �  �  �  �  �  �  �  �  �  �  �  �������������������������                                                                     <    <          <    <                                          <    <          <    <                                                                     ������������������������UUUUUUUUUUUUUUUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUUUUUUUUUUUUUUUU��������                                                                                                                                                                                                                                ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       @U    TU       |Y   @U       Y   PU      �U   T       ��U%   U       ��U  @U        ��Z  P        ��^  T        ��SU  U       ���CU PU        ���@UU        ���@TU        ���PUUU        ���TUUU         ��?TUU         ��TUU          ��TUU	         ��T�Z)         ��P��%         �  P��%            @��&             ��
             ��
             ��
             ��
             ��
             ��
     @      ��
     T      ��
    @U     ���
    TUU    ���
    UUU�  ����
    UUU�i ����       ��) ����       ��� ����      ���������      ���������       ���������       ���������       ��������*       ��������*        �������*        �������*        �������
        ���ꪪ�
        �������
        �������         ������         ������         �����            ����            ���*            ���*            讪
            ���
            ���
            ���            ���             ��              �              �;              �*              T
              T	              T              T              T              T              U              U              U             @U              PU              T              T              PU              @U               U               T              P              @                                                              �               �             ��             ��?             ��?             ��            ���            ���    U      ���   @U     ����   T       ���   U      ����  P       ���� @U       ����_UUU        ���WUUU         ��UUU         @UUUUU         U�UU          @UUUU           PU�UU           TUUVU           UUUVU          @UQUU          PU@UV          U UU         PU UU�       UUUU TU�      PUUU  XU%      TUUU  hU*            ���            ��j            ���
            ���)            ����           @����           ����j          ���j�          @����	          `����
          ����j*          `����*          `����*          ������          ������          ������         h�����         ���ꪪ
        �������
        @��ꮪ�*        �������*        �������*        ����ꪪ�        ��������        ��������        �����       ��ꪪ����      ������n��      ���������
      ������kZ�	      ����SU      �������CU      ��ꦪ��`U       ������
U       �ꪪ� T        �Z�� P        �W   PU         P   @U         P   @U         P    U        P    T        @    T        @    T        @    P        @    P        @    @        @    @        @    �e        @    @U        @    @U       @            P     �       P     	       TU     UU                U    @U       PU   Te=       @U   Te�        P   TU�       @U   XU�        U  TU�        T  ���        P  T��?        @U  U���         U U���        TU@U��        PUD��?        @UUU���         UUU��         PUU��          UU���         `UU��?         h�V��         X�j��         X�j           ��j            ���             ���             ��*             ��*             ��
             ��
             ��
      @     ���      @     ���
     PU    ����    @UU    ����  �jUUU    ����
 �ijUUU    ����* h��       ����� ���       ���������
       ��������
       ��������
       ��������
       ��������
       ��������
       ��������        �������
        �������        �������        �������        �������        �������         ������*          �����*          ���*            ���*            ���*            ���+            ���*            ���
            �j�            ���             �              �+              �              �              �              `              P              P              @              @              @U              @U              @U               U              U              T              T              U              U              U              @              @              P              T                                                ?              ��              p�             |Y_     T     _U_U     @U    �_U_U     U   �_ZTU    P   ��@UU    @   ��? TU     U   ��? PU     T  �� T     PU  �� U     @U �_U@U      UU TU TU       TUPVUVU       @UUUVUVU        TU�ZUZU        @U�ZUZ          T�j�j          @����           ����           ����           ����           ����            ����            ����            ���;             ��*             ��*             ���            ����            ����           ����
           ����
           `���&           ����*           ����j           �����         ������         @����j
         ������         ������	         ��j���)         h�����&         ��j���%         ������*         �������         �������        ���i����        ���ꪪ��        ��������       ��������       ��������       �������j       ��������
       �������j
       ��������)       ��������*       ��ꩮ����       U��������       U����
�     @U  ��� �     @U  T�
      @U   T ��      PU   T         P   T         P   T         T   T         T   T         U   P         U    P        @U    P        @U    P        PU   P        PU   P        TU    P        U    P        U     T       @     T       P     T             U                                                          �      �?      |?      �?    �
�?    ��V5    ���    ���    ���*    ����    ����   ����  �����
  ���*�  �����  �����    �*�    ��*    ���
   ����   �*
�    ����    ����    �)��    h���    ����   ��
�   ����   ����   ����
   �*��
  ��*��
  ��
 �
  �� �   �  �  �
 ��   �
 ��   �
 ��   � �*   � �
  ��  �  �*  �  �  �   �  <   �  ?  �   �  ?   �  ?  �?  ?   �   ?  �?   ?  �     �                                               �      p-      �?      Կ      ��      x      �      P      �     ��     ��    ���
    ���
   ����
   ����
   �
��
   ���
   ���*   � ��*   � ��*   %����  ��*� @����   ����
   ��*     ��*     ��
     ���     ���     ���    ���    ���
    ���
    ���*    ���*    �*�*   ��
�*   ���*  ��* ���� �* ��� �
 �?   �
 �   �
 �   �
 �   � �    � �    �     �     �? <    ���     ���     000    ���                             7      ��      ��     ��     �W     �U      `V      @U      �     ��*     �**    ��**    ��
�    �*��    ����   �����   �
���   ����  �* ��� �
 ���
 � ���
 T ���
 T ����*  ��*�*   ��* �   ��* �   ��� �   ��� �    ��      ��    ���    ���
    ���
    �
�
    �*�
   ��
�*   ���*  � �* ���* �* ���
 �* �?   �
 �   �
 �   � �   � �    �  �    �      �       �      �      ��0     ��0         ���                 �      �      @3      ��      0�      �_�*    U��    PU��   Zժ�  �jժ�  �����  ����  ����  �����  ���.�   ���>�   ��.�   �n *   �x��*   ����   ��*
   ����*   ����*   �����   �����   �����  ��ꯪ
  ��ꯪ
  �����
  �����*  (����*  ��
�*  ��
�*  ��
�>    �
��    � �   � �   � �   �
 �*   �
 �*   �* �*   �* ��   �*  �   �*  �   ��  �   �  �   �  �   �  �?   � ��   P 0�   � ��  0��  �  ��  �  ��                     �       �      x      �?      �      �>      T-      T      P      P*      ��
     ���     ��*
    ��*�    ��*�   ����   ����
   ����
   ����
   ��� *   ��� *  P���X  ����P  �/��
@ ���
     ��
     ��
     ��     ��     ��
    ���
    ���
    ���*    �*�*    ���*    ���*    �*�*    �
��   ����   �
���  �
 ���� �* ���� �*   �� �*   �� �*   �� �
   �� �    � �    � �    � �?    ���?    <��?          ���                     0       �       �     �_     ��     ��      U
      �	      U      �      ��     ��*     ���    ���
    �
�*    ����    ��*�   ��*�*   ��*��  ���* � ���* � ���* � ���� @ ���  ���  � ��
   * ��
   * ��
    ��     ��    ���    ��*
    ���*    ���*    ����    ����    �*��   �
���   �
 ��  �
 ���� �
 ���� �*   �� �*   �� �*   �� �*   ��  *    �  ?    �  ?    � �?      ��     ��     ��     000     ���                                                                                                                                    �   �  �? ��  ��  __ __ �� �� __ __ ��  �5  � �    �� ���  _?  _/ ��� ��� �_� �_� ���  �� 0_? 0\� 0�� 0�  �  � 0� 0�� 0\�  _? ��� ��� �_� �_� ��� ���  _  _? ��� ��     �  �  �5 �� __  __ �� �� __ __ ��  ��  �?� �                             ����<������ }= w}= ��? ��  �                                ��� ��3��� }= w}= ��? �0  �                             �  <���� ��7 |}� |}� ��� ��� �                                 ���� ��7 |}� |}� ��? �0  �            � � @P �P  <  \  ]  u  � �u��u�  �7 ���                � � �� �C� _} \] ]] uW �U  u]  t  s�  �0 � 0          
�  ((     �  0  0  �?  �  	�  �  _�  �?  ?�                0�0 �3 ��  �  1  0    �,  >2  0     �               0  �� ��� ? �?� �"� ��  �                         �   � ����G� =��3 0�?�>�< 0  �   <                             ? ���0�� �� ���?���0' ��  0                             ���0��?�< ����� <�� �  �  <                                   T: @�� ijZ����6WW�?�W� �  �              UU      UU      UU      UU      UU      UU      UU      UU      UU      UU UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU     UU      UU      UU      UU      UU      UU      UU      UU      UU   UU      UU      UU      UU      UU      UU      UU      UU      UU      UU    UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UU      UU      UU      UU      UU      UU      UU      UU      UU                                                                                    UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU      UU      UU      UU      UU      UU      UU      UU      UU      UU   UU      UU      UU      UU      UU      UU      UU      UU      UU      UU    UUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUU     UU      UU      UU      UU      UU      UU      UU      UU      UU      UU      UU UUUU UU UUUU UU UUUU UU UUUU UU UUUU UU UUUU UU UUUU UU UUUU UU UUUU UUU  UU UUU  UU UUU  UU UUU  UU UUU  UU UUU  UU UUU  UU UUU  UU UUU  UU      UU      UU      UU      UU      UU      UU      UU      UU         UU      UU      UU      UU      UU      UU      UU      UU      UU      UU UUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUUUUUU UUU  UU      UU      UU      UU      UU      UU      UU      UU      UU    �|=_��������?��<<O�S�_���?�                                                                                                �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?    0<<?�?�<<0  ���?    �?��    �������?���?<  <<  <�  �����?� ��  �?  �  �      �  �  �  �  �  � ���������������� �  �  �  �  �  �   0 < ����< 0         ����      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                UUUU���  p  p��p��p��p��p��p��p��p��p  p  p���UUUU��������WUUUUUUէ�UUUU�ڧ�uUUu�ڧU�UU]UڧUUWUWUڧU�]�]UڧUUwuWUڧUU��UUڧUUuuUUڧUU��UUڧUUuuUUڧ�U�_U�ڧ�UUUU��WUUUUUU�����������������WUUUUUUէ�UUUU�ڧ�U�WU�ڧUU]]UUڧUU�wUUڧUU]]UUڧUU�wUUڧU�]�UUڧUuWuWUڧU�U�UUڧUuUUWUڧ�]UU]�ڧ�UUUU��WUUUUUU�������������WUUէ��ڧ��ڧUUڧUU�WUU��UU�WWU�W�U�Wuw�W���WUw�WUw�WUw�W���Wuw�W�U�WwU��UU�WUU�WUUէUUڧUUڧ��ڧ���WUU���������WUUէ��ڧ��ڧUUڧUU�WUU�WUU�WUU�WU��WUw�W�]�WwW���U���U���U�WwW�W�]�WUw�WU��WUU�WUUէUUڧUUڧ��ڧ���WUU�������������  �  �  �  �  �  �  �  �  �  �  �  �������������������������                                                                     <    <          <    <                                          <    <          <    <                                                                     ������������������������UUUUUUUUUUUUUUUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUUUUUUUUUUUUUUUU��������                                                                                                                                                                                                                                ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������          �     �? 
  @���
 @֟��  �V��Z* �u����  V����  Xe�V* T�Z��  @UUU*   TUeT  UiU  TEYUU   @IYU   �V�Z)   �� ��   �*  �                          �     �? "   J����   j֟`�   �V���  �u�j�  �V�j*  TXe�
  P�Z�    UUU*    PUUd     UUd�   TUd�
   @d�B   �YUU   �	U     	P    T      P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �G�����? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ����������������������������������������                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                     �               �                    @�               �                    @�               �                    �?                �                    �                �                   P�                 �                   �>                 �                   �                 �                   �                 �                   �                  �                   >                  �              ��? �  ��              �             �U�� � �_��            �            �GD��� U<?            �            |U �>� �UE �0            �           �WU ��� <Q�3            �           �QUE���<�CT�?�            �           _UQ��?0D@�?�           �          �SE �>?D�:
�          �          0U  ��  � �?          �          EP@   ���  �**�0          �          Q   ��   ��*(3          �         �@AT         ���*0          �         0D  �   <    ��*�         �         p@ �?  �?    � ?         �          E   �  �    ���(0         �             � ?    ��*��         �             ?�     ��
�        �              < �      ���*        �            �� �    ����+        �        �     �U��    ���         �        �     |U=|U    �����        �        �     \U5_U=    ��(�3        �        �    �WU�WU5     ���0        �        0    �UU�UU�     �����        �        0    pUU�UU�    ������        �        0    pU��UU�   �����        �        0    |U��UUU      �?�        �        0    \U��}UU   ? � �  �    �        0    _U���UU   �8�<� ��    �        �    WUU��UU    �< ? ��    �        �   WUU�UU � <���� ��    �         �   _U�UU   �3�?  ��    �         �?  �W� WU�   ��?� ���     �          �   �? \U� �����?  ��?     �          ��     |� 0  ���   ��     �           �?    �?  0�� �   ��     �            �       < *��   ���      �             ��      < ��    ��?      �              ���������?     ��      �                             ��      �                            ���   U  �     T          �������    ���UU�  �TUUUU�       ��      �    � ���WU�������      �     �   �?  P5@�����?�������     �     �    �� T@�����?�������     ?      �      �0 UP�����?�������    �       �       @� P? �O���   �   �      �?       P5 �? ����        <       ��     � T �?@����       �      ��.     0 U �@����       �      ��     @� �@����       <      0 �     P5 �@����             ?��0    � T0 �@����      �      ���3    0 U� �?@� ���      �      ����0    @� � ��@� ���      �      ��� �    P5 � ��W� ���_      0     0����   � T � P���U����     0      �:��   0 U � @��������  @ 0<     0��> �   @�  �  ����� �T� @U= 0�    ���. <   P5  ? UU���� �P�@U�? 0      �3�  � T �? �_��� �PPU��? � �    ���?   0 U �? ��_U  �PQU���� � ��    ��    @�  � ����W �P_����� �  �   ��     P5 �? �����? �P����?� � �?   ��    � T �  ����? �P���? T    �? ��:    0 U��>   ���? �P��?  �     ��:    @�����   @��? �P�  @�      ���    P���?�    U�?  �P?   U�      ��   � T�����   T��   �P=  T��      ������? U����  @��   �   P���      ��   @Տ��0 @U��    �  @U���  0     ��  P5����0 P��    �  U���?  0     ���� T���� 8 ��?     � U����?  0     ��� 0 U��?� ��     � �����  �    �< @� ��3� ���    � ����  �  �  � P5 �� ���U   � ��@�    �� ���6� U<��?  ���_U � �? P�      ����50@���� <@ ����  � P P?     ��UêN5T= �?��@� ����  � P P? U  ��Uë�5S� ���#� @� ���  �    �T� < �����>�U? ������ P�_ ��  �    �C�� 0 ��� �>��  ��0;�3 T��W P?  �    �W�� � �?  �:   ����0(< ���@=  �   @���� �     ��    ��??
  ���_    �   P��?      ��   �
���   ���E  �   ����T�     ���   ����@����_  �   �����  <   ���   ��2� P�? ���  �   ��?P��  �  ����   ��2���? ���  �   ��T�� �����  ���������?  ��  �  @�?@���   0�<?   �?� ���?<  ��  �  P�T���  <������ ��
� ���   @�   �  P?@����?  �0� ���#�*��    @�   �   @U��@�   ���
�*?�*��̰�`�    @9   �   UW�� �   �?;����0�?��H?         �   ���� �   ����"��������R?         �   ���� �    �����������P?   P     �   ����? �?          ������P�   �    �   ��?@�@�              �P�   T?    �   P�@�@�W               P�  P?    �   P� ���             PP�  P?    �   @� �T�?             �@�  �?    �    � �P��            @�?@��  �?    �    �?   T��OUU      U���C�� �    �    ��  ���O��UU   T������?U�    �    P� @���O����  T��?��?�����     �    @�7 T��O���� T�����?��T����     �    @�� ��O�O��� ���S�����O���     �     ��C��C�C�P�?@��@���P�?���     �     ��S��P�C� �? �? @�W� ��P��      �     P�T��S�S� �? �? @�_� ��P      �     P���_�S� �? �?  �_���        �     @U�����S�  �? �?  �_�C��?        �      ��� ��S�  �? �? @�_�W��        �      P�? ��S�  �? �� U�_��T�       �      @� ��P�  � �� U�C�� @�?       �       � ����UU� ��U��C�  �       �       T ������� ����@�  �       �       T  ������� ���? @�           �          �������  ���  �           �          �?�?��   ��@� �?           �          �?�?T�   P� � �?           �          �?�?@�  P� �? �?           �         @�?�? �  P� P� ��          �         @�?�? �?  P� @���          �           ?�? P�  P� ��?           �           @�� @� P� ���           �           @��  � P� P�             �                � �� �             �                   �?                 �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �����������������������������������������                    �� �� �� � � �8� �� �� �� � �� ��.0� �� �� �� �� ��. � �� �� �� �� �� �� �� � � �� � q � �� �    q� 0� �� �� � � �� �� �� �0�.� �� �� �� � q� � � � ��.� �� �� �� �� �0�   .�.�}�T�.���}���.�.�}�T�.�}���}� ��}� �� ��.���.� ��.�}�.�}�}�����}�   T�. �}�T�.�}0������ ���.� ��.0�}�.�.�}� �� �� ��. � ��}�.�.� �� ��}��0�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?    0<<?�?�<<0  ���?    �?��    �������?���?<  <<  <�  �����?� ��  �?  �  �      �  �  �  �  �  � ���������������� �  �  �  �  �  �   0 < ����< 0         ����      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                UUUU���  p  p��p��p��p��p��p��p��p��p  p  p���UUUU��������WUUUUUUէ�UUUU�ڧ�uUUu�ڧU�UU]UڧUUWUWUڧU�]�]UڧUUwuWUڧUU��UUڧUUuuUUڧUU��UUڧUUuuUUڧ�U�_U�ڧ�UUUU��WUUUUUU�����������������WUUUUUUէ�UUUU�ڧ�U�WU�ڧUU]]UUڧUU�wUUڧUU]]UUڧUU�wUUڧU�]�UUڧUuWuWUڧU�U�UUڧUuUUWUڧ�]UU]�ڧ�UUUU��WUUUUUU�������������WUUէ��ڧ��ڧUUڧUU�WUU��UU�WWU�W�U�Wuw�W���WUw�WUw�WUw�W���Wuw�W�U�WwU��UU�WUU�WUUէUUڧUUڧ��ڧ���WUU���������WUUէ��ڧ��ڧUUڧUU�WUU�WUU�WUU�WU��WUw�W�]�WwW���U���U���U�WwW�W�]�WUw�WU��WUU�WUUէUUڧUUڧ��ڧ���WUU�������������  �  �  �  �  �  �  �  �  �  �  �  �������������������������                                                                     <    <          <    <                                          <    <          <    <                                                                     ������������������������UUUUUUUUUUUUUUUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUU  TUUUUUUUUUUUUUUUUUU��������                                                                                                                                                                                                                                ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������H�Z���8 � �� ��� ��� ��� ���� �� �  �� �  ���� �r� /�ά ��h�� ���� ά �� �  �� � � �� ��� ���  ��έ έ �� �  �� � ��� ��� ���  ���� �D� /�L� /� /��� �  ��� �� � � �� ���  ��� i�� �  ���� � ��� ���  ��� 8��� �  ���� �\� /�LL� �� �� �z�h`xH�Z�� 
�� �� � �� �� �2 �� �3 �  ���� ���� � JJ��-8 �� i� � i � �3 �3 � �Ȁ��2 �2 � �
�� �3 �L϶z�hX`H� �8  �����8 h`H�Z�/���� ���� ��z�h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ���ة��  ��� � �? � � �@ � �ߍ& ��" � t ���� �� �� � ����� ��� � �� � �� ��XL��H�Z�9 �= � ��<�=  D��= �: � ��<�: �' �� �р v� � ���:  ��z�(h@@                ���(�� �ـ��+ �y  �� �� �� p� �� �� %® ��� �  � Hí� ��
 � ����� � �� �� <ҩ��- � ��� �  �� bʮ, ��� ������y �G ��y  �� ƭ4 ���L���. �/ �0 �G �y  ��' �����& L�����& L�����8 �<�= �- � �� �� �� ����$�� �� �� �F�� �R�� �A�� �N�� �K�� ��� �. �/ �0 �� ��� �* �; �< �1 � �, �� �� `H�Z��' ��� �@�(  �� ڢ �
 �٭  ������ �Q� �� g����߀� ��z�h`H ܩ� ���  � #ܩ
�  �� � #ܩ� ��  � #ܩ� �2�  � #ܩF�  �� � #ܩ� �Z�  �  #ܩ� �n�  �! #ܩ
�  �$� �)�  zܩ�'  ��ɿ�> u߭' ���$� �
�  �)�  zܩ�' �֩$� �  i�  �)�  z��' ���з�' �����& ����& h`Hڢ �H����� ����� � �� �� ѩ��- �  ���� �ٜ- ��h�� ���h`H � �� �Щ
� ���  � #ܩ-�  �
� � #�� � ��  zܩ
� �A�  � #�� � ��  zܩ
� �U�  � #�� � ��  zܩ-�  �� �)�  zܩ��  ��ɿ�> u߭� ���� �-�  �)�  zܩ�� �֩� �  i�  �)�  z�� ���зh`H�Z ܩ*� ��  �� �� z������ �  i�  ���+� ��  �� �� z�� � �  i�  ����  � i� ��� �� �Щ� ���  � #ܩ� ��  ��  zܩ �  �����8 u߭ ��8�
� ��  z�� L��i� ��  z�� � � L�����8 u߭ � �i� ��  z�� L��8�� ��  z�� � � L�����J u߭  �"� 8��  � � ��  zܭ 8�� L��iT�  �� � �  zܭ i� L�����M u߭  �j�#i�  � � ��  z�� � � � L��8�T�  � � ��  zܭ 8�� L����L�ĭ �  �ک	�(  �z�h`ڢ �2 �� ��� ���2 �	������� �`H�Z���- ��� �Э  ���� �ٜ-  Fƭ� �� �� �� ������ n�z�h`H�Z�� �. �:� ���  Z� yǭ. �� �/ �� �0 �� L	ǭ� �/ ���ԭ� �0 ���ȭ� �. �6����  Zǭ. �� �/ �� �0 �� �X�� �/ ���ح� �0 ���̭� �. �3���� �. �� �/ �� �0 �� ��� �/ ���ۭ� �0 ���ϩ�� �ߍ& � �  �ک�(  ����
� �و����� �D�  �� i������ #� ������ ��z�h`Hڢ �� �� ����� �� �� �����h`Hڢ �� �� ����� �� �� �����h`H�Z ܩ� ��  ��  zܩ� � #ܩ� ��  [�� � ��  [�� � ��  [ܩ� �-�  ��  zܩ� � #ܩ� ��  [�� � ��  [�� � ��  [ܩ� �<�  ��  zܩ� � #ܩ� ��  [�� � ��  [�� � ��  [ܩ� �x�  � #�z�h`H� � �� �Щ2�  �� � #ܩ� �Z�  � #ܩ2�  �� �)�  zܩ �4  ��ɿ�< u߭4 ����� �2�  �)�  zܩ �4 �֩Z�  �� �)�  zܩ��4 ���й�4 ���L�� � �� �ЩF�  �� � #ܢ ����� ܩ� ��  � #ܩ� �$�  � #ܩ� �B�  � #ܩ� �V�  � #ܩ� �t�  � #ܩ� ���  � #� ����� �� ���h`H�Z �� ���)��&  �� � � �� �Щ� ��  � #ܩ� �2�  �  #ܩ� �<�  � #ܩ� �P�  �
 #ܩ� �d�  �" #ܩ� �n�  � #ܮ  �� �٩��, L^����! �٭' ��������& �- H �h�- L������ �٭' ��������&  �� �� �, z�h`H�Z �� �����R� � ���� L4��"��� L4��(��'� L4���	8�� L4�������������i� L4����R� � ���� L4����� L4��'��(� L4���	i� L4�������������8�� L4����M� � ���� L4����� L4���	i� L4�������	i$� L4�����8�� L4����M� � ���� L4����"� L4���	8�� L4�� ����'�	8�$� L4��(���i� L4����L�ͭ� ��L<���L�̮ ��� ɠ�LI�ɀ�L�̮ ���� �  (� 6�LIν�� ��m� Ɉ�	� Ɉ�4�]� Ɉ�V8逪�q� � 8逪�q�  � (� �� ���� LI�8逪�q� � 8逪�q�  �� (� �� ���� LI� (� �ϩ�� LIή ���� �  (� 6�LIν�� ɀ��� �� (� �� ���� LIή ��� � �.�p8� ��7��d��2 �� �2 �U��!�2 �2 �2 �2 �� 8� ����5� ��x� �2 � � �2 � � ��2 � �� ��2 � �X ��LIή ��� ɀ�LI�Ʉ�	 �� ��LI�Ɉ�	 � ��LI�Ɍ�	 E� ��LI�ɐ� v� ��LI����L+έ �'��- i)�- LI��(��- i)�- LIΪ��� ɀ� �- )�	 M� ��LIέ- )�y ^� ��LI�Ɉ�'8逪�q� �- )� o� ��- )�N �� ��LI�8逪�q� �- )� �� ��- )�' �� ��LI��� �ɀ� ��� � ���  ��z�h`Hڮ �i)_��h`Hڮ �i@)_��h`Hڢ� �  M���i���h`Hڢ� �  ^���i���h`Hڢ� �  M���i���h`Hڢ� �  ^���i���h`Hڮ ��2 � �� ��2 � ��h`H�Z� �Έ�� � ��z�h`H�Z� �Έ�� i� � i� ��z�h`H�- i )��- h`H�Z�- ) �P� ���  +�(�7�� �c�� �� �C�C������$� i� � i � �C i0�C �D i �D ��(z�h`Hڮ ��� �� �� ڀ�' �� �� �� � �� g��h`H�Z� 8逪�q直��2 �i���3 �� �3 ��i��i���2 �z�h`H�Z� 8逪�q�i����2 �8����3 �� �3 ��8���8����2 �z�h`H�Z� 8逪�q直��2 ��3 �� �3 ��Ȁ�2 �z�h`H�Z� 8逪�q�i����2 ʩ�3 �� �3 �ʈ��2 �z�h`Hڢ �  �� ���$���h`Hڢ��  �� �������h`Hڢ��  �ک�(  �������h`xH�Z �� �� �� �� �� �� �� �� �� ��z�hX`�Z����  �� ������ ���  �.  [ܩ
� ���  �/  [ܩ� ���  �0  [ܭ� � �� ���   zܩ%�  z�z�`xH�Z�- )��'�* i��� �*  � �� �� � �� �� �� 6�(z�hX`xH�Z�- )��\ >�' �� �� �Ҁ%�� @� �Հ�� �Հ�� *ր��� d� �� �  ������ �� �� � �� �� �� 6�(z�hX`H�Z� �  �� � �� g�����(z�h`H�Z�+ �+ ���+ �+ � �� �������� �
���0��@� �������z�h`Hک`�( � ���  ���  x������h`Hڮ1 ��� �K�  �  �" ��4�G� �! ��1 )��W�( �D�V�( �=�1 )��U�( �/�T�( �(�1 )��S�( ��R�( ��1 )��Q�( ��P�(  x� �! �  �" �1 ��� ���  �  �$ ��4�G� �# ��1 )��W�( �D�V�( �=�1 )��U�( �/�T�( �(�1 )��S�( ��R�( ��1 )��Q�( ��P�(  x� �# �  �$ �1 �;� ���  �  �& ��4�G� �% ��1 )��_�( �D�^�( �=�1 )��]�( �/�\�( �(�1 )��[�( ��Z�( ��1 )��Y�( ��X�(  x��1 �P���1 � �% �  �& �h`H�Z�� �� �a�( � �Q�C �Q�D  ���Q�C �Q�D  ���Q�C �Q�D  ���Q�C �Q�D  ���Q�C �Q�D  ��b�( ��Q�C �Q�D  ���Q�C �Q�D  ��
�Q�C �Q�D  ���Q�C �Q�D  ���Q�C �Q�D  ���Q�C �Q�D  ��c�( ��Q�C �Q�D  ��d�( ��Q�C �Q�D  ���Q�C �Q�D  ��e�( ��Q�C �Q�D  ��f�( ��Q�C �Q�D  ��z�h`Hکg�( �1 ��� �K�   x�h�( �1 ��� �+�   x�1 �o��1 ��1 �h`Hڭ1 )��i�( ��j�( �1 ��� ���   x��1 �( �( �k��( �( �1 �M� ���   x�1 �W��1 �h`Hک� �8� �1 �1 ���1 �1 
��qm1 �( ��C ��D  ���h`Hک� �T� �1 �1 )�1 
��mm1 �( ���C ���D  ���h`H�Z�b� �� ���   z�(z�h`xH�Z�- )�$�< � ��a� �� ���   z��< � ���< (z�hX`H�Z�c� �� ���   z�(z�h`xH�Z�- )�$�; � ��a� �� ���   z��; � ���; (z�hX`xH�Z�2 � � � �2 �\i����8����� � ��	�@2 ����	����	����	����	����	 ����	����	���	@�2 (z�hX`xH�Z� �

�Laح' ��"� �)
��Q�C �Q�D �� �� � �ڢ � �C�2  ;׭2 �C�����3 � �C�2 Z�m3 ��Cz�CZ�m3 ��2 �Cz����3 �3 ���� �%�' ���C i(�C �	�C i0�C �D i �D ��(z�hX`xH�Z� �



�L>٭' ��"� �)
��Q�C �Q�D �� �� � �ڭ' ���C i8� �D i� ��C i� �D i� � � �C�2 ��C�2 ��� �����O�' ��$�C i(�C �D i �D � 8�(� � � � ���C i0�C �D i �D 8� �0� � � � ��(z�hX`xH�Z�- )�g���8 �0 �0  �ٍ0 �`�B�0 �/ �/  �ٍ/ �`��/ �. �.  �ٍ. �� ���  �.  [ܩ
� ���  �/  [ܩ� ���  �0  [�(z�hX`�2 )�
0�m2 )��2 �2 `�Z�P���� ���� ��z�`�  ���� �� �� �� ��`H�  ����h`H�9 �  ����9 ���h`xH�Z�� ��� � ��	�( �( 
��c�E �c�F  �ڢ � �E�C�� ���� �%�C i0�C �D i �D �E m �E �F i �F �ɭ( �@��ߍ& (z�hX`xH�Z� � �5����C ���D �� �� � �)�( �* 



m( i�( L��ɀ�"8� ����C ���D �� �� � �( L��Ʉ�"8逪���C ���D �� �� ��( L��Ɉ�"8鄪���C ���D �� �� ��( L��Ɍ�"8鈪���C ���D �� �� ��( L��ɠ�"8錪���C ���D �� �� ��( L����R8頪���C ���D � ɠ��� �� ��( �>ɤ��ɡ��� �� ��( �%�� �� ��( �� �C �@�D �(� ��� (z�hX`H�Z� �@� � � � ����� ���z�h`H�Z
����6 轝�7 � �6�$��a��b��c�8�7�  z�Ȁ�(z�h`H�Z�)�JJJJ�  z܊)�  z�(z�h`xH�Z� �a��$��b��%��c��&��d��'��7�� �c�� ��2 �  ���� ���� � �-8 �� Ȳ-8 �� ��2 ��� � (z�hX`H�Z ܩ�  �� �	� ��� � �  z܈��  i �  �� ��ީ� �g�  �)�  z�� � ��  zܩ�  zܩ�  zܩ��  �� � #ܩ*� ���  ��  z� z� z� z� zܩ*� ��  ��  zܮ� � ��i���4 ���B ��A �
�� �  �����LOޭ� �$�B�A ��L���A �A � ڬ  Z�A � �B �  �$�  z�� � � �A z�  �� ���%�Li߭A �"���� � �4 i7�� �4 � ڬ  Z�A � �B �   zܭ �A z�  �� L�����8 u߭ �
�i� �*�  zܭ� i�� L��8�� �*�  z�΁ L�����8 u߭ ��8�� �*�  zܭ� 8��� L��� � �*�  z�� L�����J u߭  �� i`�  � � �*�  zܭ� i�� L��8� �  � � �*�  zܭ� 8��� L�����I u߭  �n���  � � �*�  zܭ� 8��� L��i �  � � �*�  zܭ� i�� L�����L�ݩ$�4 �� z�h`� � �$�  z�`xH�Z� ��� �4 � � �4 � � �� �� �ɢ� �ր!ɣ� �ր�' �� �� �� � �� gح � �'�7�� �c��  +�� �C�C������$� i� � i � �C i0�C �D i �D ��(z�hX`H �ڭ ɀ��C i"�C �D i�D �,Ɉ��C i�C �D i �D �ɠ��C i �C �D i�D h`xH�Z�' ���� �� ����� �� �
�� ��   �( 
��c�E �c�F � � �EC�C�� ���� �%�C i(�C �D i �D �E m �E �F i �F ��(z�hX`H�� �C ��D �  � ��C i(�C �D i �D ���C m �C �D i �D (�h`xH�Z���C �
�D � � � �C�� ����p��C i(�C �D i �D ��z�hX`xH���C �
�D � � �p�  ��hX`xHڢ �  �� g������hX`xH�Z�( 
��c�E �c�F � � �E�C�� ���� �%�C i(�C �D i �D �E m �E �F i �F ��(z�hX`xH�Z�� ��� � ��	
��c�E �c�F �� �)
��Q�E �Q�F � ���C ���D �� �� � � �E�C�� ���� �>�C i0�C �D i �D �� ��� � ��E i�E �	�E i(�E �F i �F ��(z�hX`H � �� �Щ� ���  � #ܩ(�  �� � #�� � ��  zܩ� �<�  � #�� � ��  zܩ� �P�  � #�� � ��  zܩ(�  �� �)�  zܩ�y  ��ɿ�> u߭y ���� �(�  �)�  zܩ�y �֩� �  i�  �)�  z��y ���зh`�* `� �J �K  �� �� � � � � � � � �~ � `H�Z�J ���Q�K ���.�V � ��O �P � �  ��c � ��\ �] � �  ���V �V �Q � F��c �c �^ � �K ���.�p � �� ��i �j � � � �  5��p �p �k � ��(z�h`�L �M�O ȱM�P ȱM�Q ȱM�R ȱM�S )
�����T ����U ȌL �V �W �Q � �L��X �z�M ȱz�N � ��M � ��X ��ȌX �L LF�`�f �g�i ȱg�j ȱg�k ȱg�l ȱg�m )
�����n ����o Ȍf �p �q �k � �#� �K  �� ��O �P � � �\ �] � � `�Y �Z�\ ȱZ�] ȱZ�^ ȱZ�_ ȱZ�` )
�����a ����b ȌY �c �d �^ � �(�e �|�Z ȱ|�[ � ��Z � ��e ��Ȍe �Y L�`H�Z�R )?	@�s �R 4��-s �s �W �T��S )@��J��s �s ȌW �T����W �S �W �s �~ ��~ � z�h`H�Z�_ )?	@�s �_ 4��-s �s �d �a��` )@��J��s �s Ȍd �a����d �` �d �s � �� � z�h`H�Z�l )?	@�s �l 4��-s �s �q �n��m )@��J��s �s Ȍq �n����q �m �q �s � � �~ � z�h`� �~ `� � `H�Z�y 
��K��z �U��| �K��{ �U��} � �z�M �|�Z ����L �Y ��X �e  F� � �� ����J z�h`H�Z����g ����h �f ��r  �� 5���K z�h`H�Z����g ����h �f ��r  �� 5���K z�h`AaaSEEaCOMPLETE$PICTURE$YOURaNAME$WONDERFUL$aaGOOD$aCORRECT$CHOOSEaACT$CHOOSEaMELODY$CHOOSEaSCENE$SCENE$SELECTaaRESTART$PAUSE$MELODY$CHOOSEaBLANKaBLOCK$ACT$CONGRATULATIONS$CONTINUE$END$BYE$PROGRAMMEDaBY$MUSICaBY$GRAPHICSaBY$FRANKaGU$LIVYaSHOU$JOHNaBAN$MAGICaCUBE$RACINGaINaWOODS$ROLLINGaBALLS$HAPPYaANGELS$BRAVEaSKATER$CHARMINGaDANCER$ANYaOTHERaKEYaTO$=�M�U�_�i�p�y������������� � � �����������&�0�9�D�T�b�o�|��##55GGYYll !"#$$#"! 
	  $(,048<@DHHHHHHHHHHddddddddddddddddddddddddddddddddd`\XTPLHD@<840,($ 	
$#"! 
	,,,,,,,,,,,,,,,,,,048<@DHLPTX\`dhlptx| $(,044444444444 	"!!!!!!!!!!



!$~tj`VRRRRRRRRRR",6@JT^hr|��vlbXND:0&&&&&&&&$.8BLV`jttttttttt																				

	%$#"!!!!!!"# $(,048<@DINSSSSSSSSSSSSSSSSSSSSSSW[_cgkosw{JJJJNRVZ^bfjnrvz~ $(,047777777777777777777766666<BHNRRR	
#"!!!!!!!!!!!!!!! 
	 !"					  nnnnnnnnnnnnnjfb^ZVRNJFB>:62.*&"
RRRNJFB>:640+&"~zvrnnnnnnnnnn
  	

		

     %+17=CIOU[agmsy%+17=CIOU[agmsy%+17=CIOU[agmsy%+17=CIOU[agmsy     
		
 
		 ",6@JT^hr| *4>HR\fpz#-7AKU_is)3=GQ[eoy *4>HR\fp!+5?IS]gq{	'1;EOYcmw ����
��
�
�UKL
YF VN 	KQMK
	 
M CX	
  �@���@��� �`�`����             ���������`�@� � ���������`�@� � ���������`�@� � ���������`�@� � ���������`�@� � ��������`�@� �� �����                         �@����� �@����� �@����� �@����� �@� � ������������@�     �@����� �����@� ����
�
�
�
����DLT\����     ����!� ����	
���"����#������DLT\��������CCCCHHHHMMMMRRRR $ $@@XX@@@@XXXX @��CHMR$d��CHMR $[[[[[.� �� �� �(��@� �� �(� ���.� �� ��    �(� �
� �
� �� �� �� �<�� �� �� �(� ��� �� �(�    �� ��� �� �� �(� �
� �
� �� �� �� �<� �� �� �� �(� �� �� �� �(�    �� �� �� �� �� �(�� �� �� �(�    ���.� �� ��@� �� ��� �� ��� �� ��� �� ��   � �� �� �� �� �� �� �� �� �<� �<� �<� �<�    <� �� � _� (� �� �� � _(� � �� �� � _�    K(� T
� _
� d� q� T� <� �� q� T� q(� � �� q� T(�    q� � �� q� T� G(� K
� T
� q� d� _� T<� K� _� d� q(� w� K� Y� j(�    q� � T� d� q� ?(� �� T� j� q(�    � �� �� � _� �� � _� �� w� _� �� q� _� �� j� Y�    �� j� Y� � _� O� � _� K� G<� d<� _<�    K� Y� q� w� d� q� �� � �� �� �� w� w�    q� � �� �� �� w� w� q� � Y� d� �� �� q� w�    �� � �� �� �� �� �� �� w� �$� K� K� Y� Y� j� j� � �� d� ��    Y� �� T� � T� T� d� d� w� w�    � �� q� �� d� �� Y� � Y� Y� q� w� d� q� �� � ��    �� �� w� w� q� � �� �� �� w� w� q� �    q� d� q� d� K� q� � q� d� j� d� j� d� K� q�    � �� �� �� � �� �� �� �� ��    �� � �� �� �� �� �� �� � �� ���.� � �� �$� ��   .$� <��.�T����� <�.�T�h���   �� � �� �� �� � �� �� �� �� �� �� � �� �� �� ��    �� �� �h�T�.�� �h�T$�.���    �� �� � �� � q�  � �� �� �� �p� � d�    d� q� �� �� � q�  � �� �� �� �p� �� �� �� ��    �� �� �� � �� q� � q� q� q� q� q� _� � q� �� �� �� T� T� T�    T� q� q� d� q� � �� � q� q� _p�    _� K� ?� K� ?� 8� ? � K� T� �� �0� �� �� � q� d� _� T� K�    ?� 2� 2� 8� G� G� ?� 8� ? � K� _� T� 0� ?� G� K� T� _� d� q� �    _� _� _� _� _� T� K� ?� K� 8� ?� 8� 8� 8� 8� 8� /� ?� 8� G� K� T�    *� *� *� *� 8� 8� 2� 8� ?� K� ?� 8� 8� _0� ?� K� ?� 8� 8� _�    �� �� �� �� �� �� �� �� ��� �0� Y� K� C� K� Y0�    �� �� �� �� �� �� �� �� ��� �0� �� �� �� �� �0�   h�h�.� �� �� �� ���.���   h�h�.� �� �� �� ���.���    �� �� �� �� �� �� �� �� ��� �� �� �� �� �� �� w� w$� �� ��    �� �� w� �� �� �� �� �� ��.� �� ��.��.��.�h$�   .�h�h�.�h�h�.��.��h�h� H�   ��������h�h���   h�h�.�.� ��.�h�h�����.��� �h�h�h�h�.���h�   .�.�h�h�.������������$�    ��  /2�    �� �� �� � �� �      �





		�	
	 �
�_�������k�e�������y� ���  ���  ��=������k�  ������2���  ��A�����+��  ���^�����R�  ����#�����[�  ����6�u���  �P���
�  D������  �����  ��2�@� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0�@P`��� ��������������������������������������������                                                                                                           [� ���