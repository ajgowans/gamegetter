                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �                                                                            �                                    "�                                     "                                     "�                                    , ��                                    ,��                                    ,���     �������������������  ���?      ���     0                      0     ,���     0                      0     ,���     0                      0     ,���    0                      0     ����    0                      0     ����     0                      0     ����     0                      0     ����     0                      0     ,  �     0                      0     ���     0                      0     �  �     0                      0     ����     0                      0     ����     0                      0     ����     0                      0     �
 �     0                      0     ����     0                      0     �
 �     0                      0     ����     0                      0     ����     0                      0     �"��     0                      0     �"��     0                      0     �"��  �  0                      0     �"��     0                      0     �"��     0                      0     �"��    �0                      0     �"��  �  0                      0     �"��  � �0                    ���?     �"��  ��0                            �"��  ��0                            �"�� ���0                           �"��  ��0                  (         �"�� ���0                  (�
        ���� ���0                  *�        ���� ���0                  "�
   �  ����� ���2                   �
�
 �  ����� ����2                   �
� �  �� � ����2                  , �
�* �������������2                  ,  �*�� �* ���������2                  , �� 
 *�������"2                  ����  
�* �������" 2                  ������*���
�"���  8                  �������*� �"����*��8                  ���"���
��(��"��  ��8                  � ��������(��"�� �*�:                  ����*�����* �"��  " 0                  �(��
�
���*
�"��
��"0                  ����� ���*
�"��
��"0                  ����������* �"��
��"�2                  ����
 ����*��"�� ��"�2                  ����*��������"�� ��"�:                  �������������"��*��:                  �������������"�� ���:                  �������
  ���"�� ���:                  ������    ���"�� ���:                  ���      ���"������:                   �����������"�����"�:                  ��
  
  
 ���"��*��"�:                  �     
 ���"��*��"�:                           ���������"�:                           ���������"�:                           
��������"�:                  ��        ��
�����"�:                           ���������"�:                          ��������"�:                        *  ���������"�:                       �� * �������"�:                      ��*   
" �����"�:                      ��  
  *�����"�:                           
�**�����**0                           �  �����*8                           ���������*�:                           ���������*�:                           ���������*�:                           ���������*�:                           �����������:                           �����������:                           �����������:                  *        �����������:                  �        �����������:                  ��
       �����������2                  ��        ����������
0                  �
        ���������* 0                           ���������  0                           �������� �?                           ��� 3����0                           �� <       0                                  ����?                           �������   0                           ��         0                  ��               ���?                  ����            �   0                  ������?   ��   �   0                   �����������  �   0                     �������
 < ��   0                       ����� � ��   0                           
   ���
   0                  <           ����   0                  �    ����   ����
   0                  �   �      � ��    0                    ��       � ��*   0                   ����       � �
    0                   ���        ��
   0                   ���        ���    0                   ��*       �  �
   0                   ���         �
    0                   ���      �   �
  0                   ��          ��    0                   ���      �* ��   0                   �
�
        �    0                   ���      ����
 ��  0                   ���+         �*    0                  �*   �              0                    �
        ��  (  0                   �
��              ��������������������
   (        ��            �*          ��*             �*      ���   ��*        ���                     ���*              ��                       �*
          (�                            "                                  �          ����                      ������           ��                          ��        �                                                                                *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��                               0   ��?�                              ��    ?��?                              ��   ���                              �?   ���                              < �   ��?  ?                            �  �� ��                                 �� ��                              <  �� ���                              �  ��  ��?                              � �������                               �������                              < �������?                              � �����?                                ������                                �����3                                  ����                                  <���?                                   ����                                   ���                                    ���                                 �����                                 ��?���                                �������+                               ���������                               �� �����?                             ��   �������                            �   𿪪
��                           �    ����
 ��                          �    ̬��
 ��                         �    ���
  ��                         �    ����   �                        ?    ���*    �                       �    � ���    ��                       �   �? ���     �                      �    � ���      ?                      0    �����                                �? � �                                 � � �                                 � �  �                               ��  �  �                               �?  0  �                               �  0   ?                               �      ?                               �       <                               �       �                               �       �                                     �                                     �                             �                                     �         ?                             �         �                                       �                                       �                                      �                                                                              ?                                       �                                       �                                      �                                       ?                                       �                                       �                                      �                                       ?                                       �                                       �                                      �?                                       �                                       �                                      �?                                      ��                                       �                                      �?                                      ��                                       �                                      �                                      �?                                       �                                       �                                      �                                      �?                                       �                                       �                                      �                                      ��                                       �                                      �                                      �?                                      ��                                       �                                      �                                      �?                                      ��                                       �                                      �                                      �?                                      ��                                       �                                      �                                      �?                                      ��                                       �                                      �                                      �?                                      ��                                       �                                      �                                      �?                                      ��                                      ��                                      �                                      �                                      �?                                      ��                                      ��                                     ��                                      �?                                      �?                                      ��                                      ��                                     ��                                      �                                      �?                                      �?                                      ��                                      ��                                     ��                                     ��                                      �                                      �?                                      ��                                      ��                                      ��                                     ��                                     ��?                               �?    ��?                              �?    ��                             �?��   ��                            �   �  ��                           �?      � ��                          �?����?  � ��                        ��     ��?���                       ������   ����                      �?  �?�   �3 ��                   ��?   ?�?���<  ����                 ��    � 0�� ?0 �              ��� 0�<���� ��  �<�            �?     �<  0�   � ��<�       ��<� �0�        �3 00<��< �  @   ���� ��0�����000�  3 �<   @ U�?    ��   � ��� �? �03  ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?      ���                      ����������������                  <<�������?�  ��:�:�:�:�3 �w=��\=�5  0  <<��W�W�\5��<?��������<����.�;��;��PT�W�_�_�WTP<0���?��?��?�0��?���������?����W�����W����??���?��?���0000��������?�?�����0������0��?�������?0<<?�    ?�<<0H�Z� �� ��� ��� ��� ���� �� � �� �  ���� �r� 
��� 8��� �ܩh�� ���� �� 8��� � �� � � �� ��� ���  ���� 8��� � �� � ��� ��� ���  ���� �D� 
�Lʃ 
� 
��� � ��� �� � � �� ���  ���� i�� �  ���� � ��� ���  ���� 8��� �  ���� �\� 
�L0�z�h`xH�Z�� 
��{� �{� �� � �� � � �F�� ���� � JJ��- �� i� � i � � � � �Ȁ�� � � �
�� � �L��z�hX`H� �  ����� h`H�Z�/���� ���� ��z�h`����? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                           C� �Ʃ  �� �ĭ2 ��  �ɩ��  \ŭ � ��Z�  V� V� V�  ��L&��k ���L�� #ív ���L؇� � �����	 �� �Lx���	 �� M�Lx��� �� {� B� {� B� {�Ll���	 �� ]�Lx���7���  N� ��Ll�� ��  N� p� �� ��} � �Li� �� :� �� �߀�`H�Z  �7 �C 0N��6 �B 0D��5 �A 0:�7 �@ 0P��6 �? 0F��5 �> 0<�7 �= 0J��6 �< 0@��5 �; 06��L Ո �� ��[� �D ������/ �- ;��[� �P ������/ � Ո (��[� �J ������/  N�z�h`�> �A �? �B �@ �C � �J �P ����`�; �> �< �? �= �@ � �D �J ����`�5 �; �6 �< �7 �= `�5 �> �6 �? �7 �@ `�5 �A �6 �B �7 �C `H�Z�/ � �Ld��(� �� � �� h� ������ � �$�  V� V��  �
�a �a � ��  ���@ B��a �� H�a� ��  �h� ��a �a � ��  ��� B��a ��  ������� �$� ,�L~��
� L~����� �$� I�L~��#� L~��� 늀I��� 늽�  �� �� �L~�� �L~����L~� 늽�  ����  �L~�� �L~�z�h`�� �P� � ��� �d� � ��� �x� � ��`�
� �P� �=  ��<  ��;  ��
� �d� �@  ��?  ��>  ��
� �x� �C  ��B  ��A  ��`Z�
���� ȹ��  ��� i7� �z`Z�/ ��
���� ȹ��  ���8�7� z`H�Z8�7� � � �� ��$� h`H�A8�7� � � �� ��$� h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ���ة��  ��� � � � � � � �ߍ& ��" � t ���� �� �� � ����� ���  �XL �H�Z�  	ǭ0 ����
� � �� � � �� �- ��
� � �� (z�h@H�' )�	� � �# �$ �% hX@                                                                                         @� �Ơ��  �����  Nʜ �  ��� B�� � �2�� @Ʃ��  ��  � � �  �� V�� � �2�� M�L-� �� d� C� �Ʃ  �� �ĭ2 ��  �ɭ- �� �í0 ���� S� \� �­k ���LU� #ív ���L(­w ���
�x ���LO� ��Э  ���� ���L-��� 7�L��ɿ�L�����	 �� �L�����	 �� M�L�����3�0 ��'��# �� {ܭk ���: .�  ����L�� �� {�L�� �܀���	 �� ]�L��������  N� ��L��� ��  N� p� �� ��} � � ŭl ���I �L�� ��0 ��	�� :� :� �� �߭- ���8 �d0� '� ��Ld��m ����8 ��Х����  �� �� '� +�5 �6 �7 �~ � �4 ��L-�Ld����  N�`�H� � ��(� � � �	�[ ��� � � ��� h�`Hک �v �w �x ��� � ��x � � ��v � � ��w �h`H�Z� � �� �\ �0�0 ��0 � �\ 
����� 车�� � �	 �� �����	 ��� ��	 �	 �� ��z�h`H�Z� � �� �\ �0�0 ��0 � �\ 
����� ���� � �	 �� �����	 ��� ��	 �	 �� ��z�h`���� ��  �� 1�`� �� ��  �� ��`� � �� ���  Nʭ5 �iP�5 �6 i �6 �7 i �7 ة�� �� �7  ��� �6  ��� �5  �� V�� � �0����� `���  ���\ �[ �[ �0�0�0�0��[ ������0 ��Z i�Z ة �� ��� �U� �Z  ��  V�� � �
��`�
� �� � �𩇍 �� � ��� � �� @�`HZ� � �� � �� �	��	0�� ����l zh`�. ���
�
������3 `� �3 �� ����o ����p ����q � ȹ���r ����s ����t ��u �	�i ��j  �o �r �p �s �q �t ��i ��j  �� � �k `Hڪ�j�




� ��) �& �h`H�Z ��
��d�# �d�$ � �! �@�" � � �#�!��(���! i0�! �" i �" �# i(�# �$ i �$ ���Ωߍ& z�h`��- �. �0 �1 �Z � � � �2 �[ �\ � �~ � �5 �6 �7 �; �< �= �> �? �@ �A �B �C � �[�D �J �P ����$�D �J �P   �`�u �} �8 � �k �m �l � �� � � ���������  �` Ĝ � � � � � � � �� �� �ߍ& `H�Z�� ���Q�� ���.�� � �ɭ� �� � �  �ȭ� � �ɭ� �� � �  1�� �� ͘ � ��� �� ͥ � oȭ� ���.�� � �� �ɭ� �� � � � �  ��� �� Ͳ � 	�(z�h`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��ڍ� �ڍ� Ȍ� �� �� �� � �'�� ���� ȱ��� � ��� � ��� ��Ȍ� �� ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��ڍ� �ڍ� Ȍ� �� �� �� � �#� ��  �� �ɭ� �� � � �� �� � � `�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��ڍ� �ڍ� Ȍ� �� �� �� � �'�� ���� ȱ��� � ��� � ��� ��Ȍ� �� ��`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����Ξ �� �� �� ͼ �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����Ϋ �� �� �� ͽ �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����θ �� �� �� � �� � �� z�h`� �� `� �� `H�Z�� 

��_ٍ� ȹ_ٍ� ȹ_ٍ� ȹ_ٍ� � ���� ���� ȱ��� ���� �� �� ��� ��  �� o� �� 1ɩ��� z�h`H�Z�� 
���ٍ� ��ٍ� �� ���  	� �ɩ��� z�h`.
� �
� �
� �
� �� �
� �
� ��.
� �
� �
� �
�    �� �
� �
� �� �� �
� �
� �
� �
� �<� ��    �� q� �
�    �
� �� �
� �
� ��.� �
� �
� �
� �
� �
� �
� �<�   \�����\�\���������.�}�.� �� �� �� �� �� ��.�   }�\���\���������\�����    �� �� �� �� �� �� � �� �� � �� ��    �� �� �� �� _� d� q� � �� �� ��    �� �� �0�    � �� �� � �� �� � q� � �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��    �� �� �� � � q� � �� �� �� �� �� �� �� �� �� ��    �� �� � � q� � �� �� �� �� �� �� �� �� �� �`�   \���\���\�����\���:�\�������\�:�������   }���}0�\���\����0��0���\�������\��0���\��0�   ��\��0��0��0��`�    /�  ,�  *�     G� C� q� K� O� �� Y� G� 5�    2� /� .� ,� *� .� %� .� *� &�    ��    �� �� �� ��� ��� �� �� �� � d�    �� /2�    �� T@� �� T� T� �� T� T� O� T� Y� T�    G@� O� T� _� T� _� d� _� T� _� T� _� d� _�    T� _ � j� �� � �� T@� �� T� T� �� T� T� O� T� Y� T�    G@� O� T� _� T� _� d� _� T� _� T� _� d� _�    T� j� @� j� O � O� O� G� O� T� O� G� O � T� T � ��    _ � _� _� T� _� d� _� T� _0� j� � j� O � O�    O� G�  � T� O� G� O0� T � G� q � q� q� j� q� w� q� j� q@� _�    0�� �@�� �� ��� �� �� �� �� �� ��    �@� �� �� �� �� �� �� �� �� �� �� �� �� ��    �� � � ��� �� �@�� �� ��� �� �� �� �� �� ��    �@� �� �� �� �� �� �� �� �� �� �� �� �� ��    �� �� @� �� � � �� �� �� �� �� �� �� � � �� � ��    � � �� �� �� �� �� �� �� �0� �� � �� � � ��    �� ��  � �� �� �� �0� � � �� � � �� �� �� �� �� �� �� �� ��    � � ��� �� �� �� �� �� �� ��� ��.�   �@�h@�   `� � � �� �� �� w� �� �� � � �� �� ��    �� �� � �� �� �� �� �� �� �`� � � �� �� �� �� �� �� � � ���    �� �� �.�� ��� �� �� �    �`� �� �� �� w� �� � �� �� �� w� � � �� �� �� �� ��    � �� �� �� �� �� � �� �� �� �� �� ��    �`� �� �� �� �� �� � �� �� �� �� �� � � � ��� �� �� �`�   ��\�h ����. �� �@���   � ��h���\�\�   � � ������� � ���@�� ������   h���� �� ���@� �� �h�h�h�� �� �.���� �\���� �   \ �� �@����� �@ ���������.�   � ���.�� �� ������� �� ����� �� ������� �    ����� �� ������� � �� ���@�@�� �� �� �    �	� �	� �	� �	� �	� �	� �	� �	� 	� �	� �	� �	� �	� �	� �	� �	� �H�   }	�.	��	�.	��	��	�}	�.	��	�}	�T	�@	�.	�	�	� �	�}H�    �� �� �� �� w� �� �� �� ��� ��@�.$�    C� O� Y� d� ;� G� O� Y� d� C� q� O� ��   	

	�	�	�		�		��
 �

		�
	�wىٓ٣ٳ�����������������$���$�^�p���C�  �͖���Z�  Fυ���&�o����  mѱ���Rқ���7�  ���ә���.ԕ���"�f�  �������b����`�  ��  �  c�  ��  zʹ����  I˫�  {΍ν�����9�  ��������!�.�T�H� �  ���� �0�h`H�  ����h`�Z �� �ɩ�)��&  -� V�
� �� �
 ��  ��� -ک� � �� V� V� �� 1ɩߍ& z�`H�` 


m_ m` �h h`�j �` � � �� �i �_ � 0+ �ڬh �� ��u ������_ � 0 �ڬh �� �	� � ?ۀ���y `�j �` � � �� �i �_ �	/ �ڬh �� �#�u �� ����_ �	 �ڬh �� ����� � ?ۍz `�h 8�	��� ��h i	��� ����� `�i �_ �j �` � � ��  �ڬh �� ��u � ����`  �ڬh �� ����� � ܍{ `�i �_ � � �� �j �`  �ڬh �� �%�u � �"���`  �ڬh �� ��` ����� �
�` �� ܍| `�h ��� ��h ȱ� ����� `�i H�i �i �  �ڭy ���h�i �h�i  <� �i  �`�i H�i �i �  �ڭz ���h�i �h�i  <� �i  �`xH�Z�j H�j �j �  �ۭ| ���h�j ���h�j  <� �j  � �k z�hX`�j �a �j �j �  �ۭ| � � �­a �j  <� �a �j  � .�Эa �j `�
 H� H�` �a �` �` �  Qݭ| � �$�a �` � �  ���� � �a �`  �� .�ɩ ��  Nʭa �` h� h�
 ` �ڬh �� ��` ����� � �| `� � �� �u ��L��� �L ޭi �_ �d �j �` �e  �ڬh �s ��
 �j �c �g �i �b �f �`  �ڬh ��+�` �c �r ��	 �` �`  �ڭ` �g �h �t �� L/߭t �� �` �g �` �`  �ڬh �` �c �r ��	 L/߭i �d �_ �j �` �s �]  �ܭ` �e  �ڬh �s ��
 �i ʎb �_ �j �` �r �]  �ܭ` �c  �ڬh �r ��	 �i �f �_ �j �` �t �]  �ܭ` �g  �ڬh �t �� L/߭i �d �_ �j �` �s �]  �ܭ` �e  �ڬh �s ��
 �i �b �_ �j �` �r �]  �ܭ` �c  �ڬh �r ��	 �i ʎf �_ �j �` �t �]  �ܭ` �g  �ڬh �t ��  3�`� �@��! �B��# �D��+ �@��" �B��$ �D��, ��} � �b �!�c �#�	 �+ȭd �!�e �#�
 �+ȭf �!�g �#� �+`H�Z�� �� �� �� �� �� �� �� �� ��� �� � � ���@��� �+Z� ��� �z�!z ୀ ����!� �#�  v� Y� <� ����} ��z�h`�Z� ��.�� � � �
��(��% ȹ(��& � �%� �
� �Ȁ��ҩ��� �� z�`� �� �� ����� �
��0��' �8��) �(��% ȹ0��( �8��* �(��& `Z ?� � �_ �'� �` �)� � �%�_ �_ � 0D�` �` � 0:� �8�
� �� � �� �!�� �� �� �� ��_ �'�` �)� �%� ��� �_ � �` � � �_ �_ �	D�` �` �:� �i
� �� � �� �!�� �� �� �� �� �%� �_ �'�` �)���� �� �� �� �� �� z`Z ?� � �_ �'� �` �)� � �%�_ �_ �	D�` �` � 0:� �8�� �� � �� �!�� �� �� �� ��_ �'�` �)� �%� ��� �_ � �` � � �_ �_ � 0D�` �` �:� �i� �� � �� �!�� �� �� �� �� �%� �_ �'�` �)���� �� �� �� �� �� z`Z ?� � �_ �'� �` �)� � �%�_ �_ � 04� �� � �� �� ��� �� �� �� ��_ �'� �)� �%�­ �_ � � �_ �_ �	4� �� � Ȍ �� ��� �� �� �� �� �%�_ �'� �)�¬� �� �� �� �� �� z`Z ?� � �_ �'� �` �)� � �%�` �` � 0:� �8�	� �� � �� �!�� �� �� �� �� �'�` �)� �%� ��� �` � � �` �` �:� �i	� �� � �� �!�� �� �� �� �� �%� �_ �'�` �)���� �� �� �� �� �� z`xH��_ ��` �n �]  ��n ��� ���n hX`H�Z�} � �� ��B� ��� � �  ��� � � V� V���  �� V� V�ة��  N� ����  @�z�h`�� �
� �Z  �𩑍 �� �  ��� �~  ��� �7  ��� �6  ��� �5  ��`� � �� � �� � �0�L��] �� � �
��0��' �8��) ȹ0��( �8��* � �'�_ �)�`  ��� � � �L��`� � � �� � �� � �0�L��] �� � � � �� �� � m} �} m8 �8 � �m m m5 �5 �6 i �6 �7 i �7 � m~ �~ � i � ؘ
��0��' �8��) ȹ0��( �8��* � � �'�_ �)�` � �_ �!�` �# �ک � �� �h �+�� �� � � � �L��`�} � � �� �
 � �
 0U�
 ���#� ȱ#� � ;� �#�� �#�!� �+� ȱ!� �+� � �!� �+�� �!� �+�
 � �
 ��� � � � Ў`�} � ���g � �	 �!�_ �+� �x����m �#�` �g �g �_�_ �b �` �c �_ �_ � 0 �ڬh �� ���_ �b �_ 0C�c �`  �ڭh � �` �` � 0� �ڬh �� �� �h �� ���	 �	 � �L9�LJ�b �_ �c �` �_ �_ �	 �ڬh �� ���_ �_ �b �­c �`  �ڭh � �` �` � 0� �ڬh �� �� �h �� ��`� �+�x���} 0����m �c �_ �c �c �G�` �_ �	� �ڬh � �� ��_ �c �` ���` �` � 0� �ڬh �� �� �h �� ��`� �_ � �`  �ڬh ��]  ���` �` �0��_ �_ �	0�`xH�Z�u � �u �u H��3� �/����' �ۭ| � �R `ۭ{ � �H� �u  <�h�u  ��LX��0� �u  �ڭy � �" �ڭz � �� �u  <�h�0� �u  w�� �u hz�hX`Hڮr �s �r �t �s �t  ��h`�j �` �i �_ �u � ��_ ��_ �t �]  ��i �_ �s �]  ��i �_ �u � ��_ ��_ �r �]  ��`�i �_ �j �` �u ���` ��` �t �]  ��j �` �u ���` ��` �r �]  ��j �` �s �]  ��`xH�u � � w��� ����� w�hX`xH� H� �  �h� hX`H� H� �  �h� h`  �� �� � ��� �(� � ��� �;� � ��� ��  ��� ��� � �� �� �� ��`�� �� � � � ���� � �� � �� B� �<�թ|� �� � � � ���� � �� � �� B� �<� V��)��&  �� ��`  �� �� � ��� �;� � ��� �N� �	 ���4 �4� �;�  �� j� B����
�����/�� �  ���� �4 �4 �0��4 �;� ��N�  �퀿 �� 1ɩߍ& `�4� �o�  �� -� j� B���������������"�� �  ���� ��1 �1 �0� ���`�(� ���  �� �2 ��� �� �&�  ��2 ��  �� j� -� B������������ ���2 �2 � ���4��2 �1�� ���2 �2 ����� �2 ��  ��2 ��  �ɀ����#�� ����� �	�� �� � �F�� ���� � �Q�� ȲQ�� �� ��`�� ��  -� j� B�������Cɿ�r��n�� �  ���� �. ��	��. �;���	��. ����. �'�  �퀯� �  ���� �. ��	��. �'����	��. �;�Ω�. ��ũ �  ���� �
�^ ��  �`�1 ��] �H� �n�  @��] �] �	� i� ��`  ��- �0� �X�  -� j� B����
�����/�� �  ���� �- �- �0��- �X� ��d�  �퀿` w� � ��� �_� �  ��`H�_� �� � � �  ���� � �� �  �� B� �|0թ� � ��� �X� � ��� �d� � ��0� �X�  ��h`� � i� � � i�
 ��^  ��`�
�^ �@� �A�  � V� B� Q�d�  � V� B� Q驌�  � V� B� Q�d�  � V� B� Q��^ �� �l� �<� �n�
  ��`� � i� � � i�
  ��`�Z� ���� ���� ��z�`�Z�P���� ���� ��z�`�Z������ ���� ��z�`ڭ  ���� ��`H�Z�0� iL� � �
  ���
  �� B� �� �  ���� � �
 � �0ל^ � �  ��� ���  �� B� i�
 �/0�z�h`H�Z� �m� �m� �8� �j �j � �� i� � i � �j ��z�h`�� �� �9� i�
 � �  T��� � �  T� B� i� 0�`��^ � 

� i8�  ���^ � 

� i<�  ��`��^ �4� i<� ��� ���
 � �  ���� � � i	�
  �� B� �y�`xH�Z�^ �m� �m�  ��z�hX`� JJ� � �F�� ���� � JJ��- �� i� � i � �� ����
 ��`H�Z� �@� � � � ����� ���z�h`xH�Z� H� H� H� H� i� � i�
 �1 ��� ����	�
�����m] ����� ����  ��h� h� h� h� z�hX`xHڮ_ ��� �` ���  @��hX`H�Z
��<� �<� � ��$��a��[��d�8�7�  �Ȁ�z�h`H�Z�)�JJJJ�  �)�  �z�h`xH�Z� H� H� H� H� �[��$��a��%��d��&����� �	�� �� � �F�� ���� � �- �� Ȳ- �� �� ��� � h� h� h� h� z�hX`PRESSaSTARTaBUTTON$NORMAL$FLASH$BEGINNER$AVERAGE$EXPERT$MUSICaAaBaC$GAMEaOVER$CONTINUE$END$PAUSE$LEVEL$TIME$SCORE$BLOCKS$aaaPLEASEaSELECTaa$ENTERaSIGNATURE$�������������������������,�D J P  � � ������'������ �c� PdxD J P F<2(
F<2(
F<2(
F<2(


  �
 ���  ��
�* �
  �
����  ����* �
  �
���� �����* �
 ������ �����
�� ��������*�
�� � �*��*� ���  � �*����+  ���  ����
��*�+�*��*  ����
��*��������*  ����¯�*��������
  �
���+�*  ��* �
 ����
�*  �
�� �������* �
�� � �*����� ���  � ��������  �* ��� ������ �*  �* ��+ ������� �*  �
���
��*����* �
     ��
��   ��
  ���*�   ���  ���*�  ���� ��
�
�*  ���� ���*�*  �*�� � �
�
 ��
�� �+ �
�
 ��� ���¯ �� �� ������ �* �� �����  �
 � �
��  �
 �+����* �� �*����* ��
 �
� �*�
 �� �
� �*�
 ��
�� ���ʯ����*�� ��������*���
 ��������
���     �* �� �
 �*   ���
���*���
 ����
���
���
��
�*��ʯʿ
 �� �
�*���� �
�* �
���
�
   ��
   ��� �   �  ��* �   �   ���
 ���  �*   ��� ���
 �*   ��
   �
 �
 �����
   �
 �* ���*�
� �
 �
 �*�
�
�
�� �*��
�
�+�*�� ����¯�
����  ���*���+���*  ���
� �+���  ���<  0�� � �? <  �� �             0 ���� � ?���  ���3�    ���3� �  � ��3�   � � ��  � 0 0 �� �� ?�             ��?���������?�                                                                       �                  0                                                              �    �            0    0                                          � 0 <             0 0 � �             0� 0             00            �  0 0      �����?  0 �      �       �        �              ��               �?   �                                  �                  �   0 � �������     �   � � ������� �0 0    � � ��� � < 0   � � �*���*� 0    0 � �+���+� �0     ��� �,� ��<0     ���������0   �  �/������/��                  �    �              �                      0   3              0   �          0      �    ��    �      � � � �     �   0 0� �  �    0  0 ��0 0   �? 0   �0  ��0    ���     � 0      � � �   0 0        0  0    �        �  0               �              ��                  0                  �                   ��������������^a�JW�UAE�BCD5�68:<>�UBD=-(�$.8B:2���9�p����K�uvwxyz{|}�lmnopqrstuvwxyz{|}�cdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}��08@HPX`hp�$,4<DLT\dlt|����  0@P`p��� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____P  0@P`pP��������P�  0@P`P  0@P`p������������������������������������  0@P`p��������  0@P`p��������  0@P`���������������������������������������                                                                                                                                                                                                          O� ���