     			      

 !"!"!"#$%&'()*+,    -.-.-./0123456  7878			9:;<3456  =  >?@     
AB!"CDEF   GH     IJKL-.MNMNOPQRSTUV  WXYZ		  [\]^_`ab  cde   fghijklm  nopqrDrD  stuvwxyz      MNMN  {|}~  �            ��������            ����� �             ��������   �        ����       �������� ����       �������� ������ ����         ������ ������������                 �j�Z�V�W�W�W���������������������?�?�?�?�?�?�?���������������着�?�?�?�?�?�?�?��WUWUWUWUWUWUWU�?U5U5U5U5U5U5U5       @ P T U@U       
 * � ���������������  �?�?�?�?�?�?�?  ���?����������  �?�?�?�?�?�?�?  WUWUWUWU��������U5U5U5U5�/�/�/�/PUTUUUUUUUUUUUUժ
�*������������PUTUUUW�W�TUUUժ
�*j�ګڠ������           ��
(�  ��"�˺��?��  � �<
<*���.��             
 @�_p����ۼ_l� �   � ��� � � @         � + �0 � �30   � ����ઠ��  
 � �����
�/�/�/�/�/�/�/  �������?������  �/�/�/�/�/�/�/  U�U�U�������������������������������,�� ��
 �  ��+�� ?    ���?*<������ �" � ��
*<��? ��������|����� ��?�?�?����  ����権 � j ���
"
�
��� � � � � �    �   ? � � ?   ������ � � � �  ���?��� ?           ��bb��        j	�/
t T@����������� z��jE�j��i��i��i��i����������������""DD�""DD�""DD0""DD0��WUWUWUWW�W�W�?U5U5U5T5S5S5T5 7 � � 7  �    ���
�(4�     �������� �EEE�jE�? PUTUVUVUVUVUVUV�  @����@         � � k�[�       � � ��������?������  �/�/�/�/�/�/�/  V�V�V��������o�O����������������U�U�U���������ϯ�����������������[ k � �      ��� �         @ T@��e W�V���VU��UViU�UvV��iY   V e*e��X�              �?���� � � � �  ���?��� ?        @���� 
��      ���( �     @�Ӱ���
 �      � ��� +          �� 0��        0<���       �� 0����      <0�0�Ό�T]tU4���P�V �  WUU�3�?1�Z��
  !�e����efe�Z �   @ �)�b   ��|?� ( 0      �:�:#?
        ��~��\�0     �����     ��㌎0�����    ���?�?�?��     �㌎0������     �?�?�?���?     T�Z��d�vT��U�̕ji��S�UUu�ͩ�      Y J%�! @ � ��찬��@     ����]  @ � � ?����6      ?�:�:�        �0<0�β        �  ��2      0�<˳��2      �  ��2�2����������PU U  �Y�%�e?iL�U���  �e�%be&XY�j���      f !��Z  U�U�U��������o�O��� �����0�    � � 3 � �     ��0 ���0��    � %# �      �2���/���� �    �2�2�2����    ���/�������?    �2�2��� �       @?�됯�p� � �   ��O��W � < �@�𬓰�@� � � <���:OW �   �0@��W���  Pt��44���u � p      n]�  0 @     ���u � � 0     N]�   p          UP��UU    ��=D�U       @UP�� ��?     4��?�?      � �� ��* ��"��  

�
�/ �*�� ��b
�*h���b�� ����*�/��*�  Tt��  �0P�T@@�
 ���0� � � 0  �*� /3      X ���0� � � 0  & � /3     W|�P U        U ?�UU    @00W0�� �      U� �� �    ����[���[����   � ��0��� ���   ? ���0�� �   �0����� � �0�   ?0���� �0  5@�@�@�@�U�U�0� ( ���00 � 0 �0� �30 0 � �� ( � ��0 � <  �� � 3< �   j�@�@�U�U�j�@���       ��(         * � 
 ( (       �( ����      + �;(8( P@� � P �(A���% � g � & ��V   P U@�P�P�T��   U Vj��� �  # l�T p2   C!0� �P   ( �� �       ( *�
�*       (8�� �      �( *�
�*       ����P`@� T  =P�S'SZU   ��T�P�P�@� U P  ���jVU    � T c�� ��  �P� �� 8  �  UU �U�U�U�����UU QUQUQU����������������������           � �                                                                                                �������?��� ? ������������ � �                                                                                                               � �                �         � �            �����������   ����0   � � ���?����  �  ����������������?�� � ?    ������� � � � ��?��?������������� ������������� ??   ������� ��0�                                                                                    � ? � �� � � � � �������    �   ? ��� � � � � � ���         ? � � � � � � � ����� �   �� �������?�����?�? ��?�?�?�?���� ������� �0�����  ? � ���?��   � � � ���������������  �  ��������� � �����?    �� �� �� � �0�0� �   �   �   �   �            ��33�<����33�<����33������33����         � 0 0 �            ���<�<����������<�<������������� �?��0�0�0�0� �0� ���              ��?�����?����������� � ? ? �������� � � � �     0 �                                                                     0               ? ? � � ������� � � � ����������?�? ? �     �      0       ���� ��� ��  0����������������  ? � ���?��   � � � ������������?� �� ������<�� ��� ������??� ?�� �������� ������������� �� 3��������������0������� �� 3�3�����������003   �0�? ���   ��0��  ����  <        ������?���0������ � ������������0�������������� ������� � ��0�<�������3330� ?   ����3 �� � � �����330� ?   ������� � � �������? �   3 �       <0 ��������� �0��� ��?�?���?�������<�<��� ��?�?���� � �����������<�� ����������?���00�������� ��� ���������?���0 ������� ��� ��0�       3 � ��   �  � 3    ��0  � � 0    �������� ���3�  ��                ? ?��??�?���� � ���0�<�������? ���?��?���� �����0��������� �0�  � ����0�0�� � �  ����0�  ? �����0�� � � �� �������?�   � � ������ 0  � � ��� ? ?� � ��� � 0�0��� � ���?�?�� ��������� � �����? ? � ��������� � � �����?�����?? �0���������0� ���������������� 3�  ����� ���3� � �������?  �0 ��������� � �?��������?�?�?���  ������0� ���0�  �??<?� � ? ��<�0� �� 0� ������� �3�������?��� � ?�?��� ?�3��?����� ��������������� ?�3��?������ ���������������� �� � �������� ����  ����?���� �?�������� � ��� �����      ��      ���?���?0�?0������ ? �0� �0����?�??�0��3������ � �0� �0�����? ? ? ?    ���� ??���?���� �� ���������?�? ����<��?���� �� ����������  ? ?      ? ? �������?     �������� � � � ��������?     �������� � � � ��? ���?��<0 ��� � ��� � �� ���� ?     ���� � � � � � ���������������������������������    ? ������� � � � ���������    ? ������� � � � ���������00����? ���� ����� � ���    ? � ��� � � � � � ����������?������?��?�����?����������  �?              ��        xآ����IՅ ��I� �)d ��� �� ������ ��Ս����� �� �  � ��d g� ܜ ԩ���� 9�  �d���8�F��� mƩ�� m�ddddd�@�A�B�C�D�E�F�G �� ؙ���2��dL䘩��� mƩ��� mƩ�� �d�������u���v��o��p �۩�o�
�p Gԩ�o�
�p GԤȘ �� �Ԡd 5݈��L�**************           **  Stage ?? **           **************  � � .� �� N� ^� 9� �� ��� �0 ��Lؙ��� �� VӠ2 5݈��`��� mƩ�� mƠ� 5݈��������d	d
ddd`�բ� mƩբ� mƩ��d��y�u���v��o��p �۠� 5� 5݈��L��***************            ** Game Over  **            *************** �  )p�6��m��n� ڽ H�m�o�n�p G�h ���m�m�m����m�n�n���@��`8�0JJJJ�g�8�0)�Jeg�� `8`� �?� ���'�\��� ���q
����q�������7����6
�����u��v��7���u��u�eu�u��v���dv
&v
&v
&v
&v
&v
&vip�u��ev�vd�?Z�uH�vH�u�����
� ƛL���  ��h�vh�uz��`�g�'�\��`Z�g	��\� u������ E�)?i
�����$�L�tz`��%�H� /��� �� �u����u����u����u` (*,.0PRTV�hJJJ
idv

�g
&v
&veg�u��v�h)
ieu�u��v�uiq�w�vi
�x�ui�u�vi�v`�g)



iH�g)�
i�h`���s0���si���  )��  )��4��l�� 5ݭ  )��  )��� 5ݭ  )��  )��� 5ݭ  )��  )���`� �{���|� �}���~����������?�dd	d
ddd�� �@�X��ddd`��
�� B� ���� ���X��X��`�d���e����e��


e����


������_�����`�����a�����b�����c�����d��_���`�� �FH� 
���m�����m���� m���ک V��� /�� ��uȑu��uȑuh�����`���	`���	`   � �   �� �� �� ��  �������	��L[��  ) �  ) � ٞ��4��0�  )�  )�%�  )�  )�/�  )�  )�;�  )�  )�E`������������`�������ک���`��ͤ����ĩ���`�����������`��� �� ���
� ���� ���� ����� V�`��@��@�`�g�O��X�,��X�g�@� ɀ�ȥ



yW��H�



yY��P΢`   ٞ���������
��}��u�~��vlu `|�}���������         �ڽ@�8~jL*���@ɀ���}PH�}Hz ���	��@�2�}H�H�oɠ��:�}P�P�pɠ��@���jL*���@�� ɀ���B��u�C��v�J��K�H�H�z� ����0L��`    ����    z {   ���'��\ `����`)��H R� ��h�����`L��LϠL�L_� ��8�

�� )��i
�����u����v���o���p�i	��� ��L��� � � @� � � B ��8�


�� )��Ƚ����ȹ��u���v���o���p�i	��� ��L��� � � � � � ������L�L�����\`
��Y��u�Z��v���o���p�i	���L��hjl��0&��)�����u����v���o���p�i	���L�۞\�i	����L��oqH�� E�)i�� Eݝ� Eݝ$h`�dg���g
&g
&g
&g}L�L�g}��idg�$�g
&g
&g
&g}t�t�g}��j�i�i�i�j�j�j�	ei�k�	ej�l�i�j ��,�k�l ��#�i�l ���k�j ��8�i���8�j���`� ��`�



i�g�



i�h��i8�g����i8�h�����`���g���h��@k������yH8�g��W�yP8�h��K��\ɑ�ɐ��Н\Lܢ���\����Z� V�z��@���!� �@� m����m�����`���`�



i�o�



i �p� )��=�ep�p����eo�o���ep�p A�Lȣ  �����!��&��E��'`dg��&g�
�&g�g���`�
)��ƣ`�)��ƣ`dg�
�&g��&g��&g�g���`dg�
�&g��&g��&g�g���`   � ���	
 �
����u���v���g�+��h�pɠ�dp����h�eu�u��v� �g�hL��  
  Z \    ^ ` b � � � )�^��o��p���u���v �ۭ��=���>���? �ϥG �ԤF�E �ԥ )�'��o��p GԠ�{ �ܩ�o��p Gԩ: �ԥ ��`Score: ��5�e�� e��`�J8����)��JJ��ܤ�0[�`[��[��[��[` ?�����/[������u���vdo��pL��  Force: �������&�u���v��o��p �۩��`*************          ** Time out **          ************* ��{���| Yܩ�o��p�ʅu���v ��L��� �{���|�㥬� ���奬� ��`���y�T�z�$�HZ�u�v�� �� <�zh�y��z����`(c)1992Thin Chen Enter. � � � �                                                                              	
                                                                                             !"#$%&'()          *+,-./0123                                                                                                                                                                                        � � �          � ��W9W�WU    ��l\_  � ���p5p\0? ��p�     �    � � � W W W�         0              � � � ���pU\�W�  �    5 � W WsW×� ;    UU[����\UpU�U�� � �  UU9U:��?   � ��UpUpU�����0 4�5���� � � ?               �� � � � � � � ��   QU��5 : : ?    _\���  ������5�5�0���@��:p����U� p @               � � \ \ W  �������? �?�              �U�U�U��������  UUU�U��:��     W W l � �    �wUuUu������    5 5 : :    �������5�5�5�0����>��p�p�p5,0�?����U�U�U� �            �����\\W > � W\\��� ���W� � �  �>���7�� � ��? :�:�5\�WU� 0��� � :         �1�5�5�5������  ,�pUpUpU������  �A�U�U�UΪê��    ��Uժ:��  �WU\U\U���� �  @�U�UU� >    �UUWUWU��� �  5���U�U���>��  ��\�p�p�����      5 � ��  ��dd L� <� <� <ݭ  )����� <����ȐL���  )�����d ���  ) �3�  )�<�  )��C�  )���  )�Σ�  )� �  )� Lª�����1���L*��������L*�`��o��p���u���v �۩�o��p GԤȘ �� �ԩ�o���J�Ȅp Gԩ*L�� Stage:?? START ���d`� ���������  ��� �����-���� Ԡ Z���Iw� z����o��p� �u��v ��L�`�������������_^FNNEzz#W4W2Yw� �o��p Gԩ��u���v G��
�o��p Gԩ��u���v G��L��(H� � Z�u ��z�����eu�u��v����y���C����y����`ey�y��z�h:м`�g�g� ���Jjj(**HJ~�~�~�~�J~�~�~�~�hJ~�~�~�~�J~�~�~�~��з����`            x   �   ?�  ��   ��   �� ��� ��?� ��� aÁ� aÃ� aÃ� Ã� �Ç� ���� ���� ���  ��  ��� ��� ���  ?�  �   �        �   �  �               � ��������  0�                   p   | |  | >  ><>  <><  80  ?0  ? g�� ����� � |p 0w� 8�����~s�  s�  � 8��������g   w   �   �  ��` /�p x<x |x|~ <x|g <y�g�s�c��`��`� � �?  �   �   �    @            

      

                                                                                                                                                                                                                                                                                                                          					 		  		  			   					                     
                                                                                                                                                                                                                                                      	 	 	 	                
 				  			                                                      		                                                                                                                                                                  
              

                                         			  		  		  			                                              								                                                                                                                                     				   		   		    				                 	   	   		 		 		 	  		 	         	   		  	
   	
	  	
  	
		
  	
	                   


		 	


   


  		


								                                 				   	
	  		  	  		   				                                             

   

                                                                                                                  							                                              	   	        

    

               	  	  	   	   	   	     	                     		          	           	  	 		 	
			
		 	
		 	
		 	
		 	  	            � ��@���������`�����[������ds���s������ _� ������������si<�s��`

�� �W�� � �����`� �/ ������`������@�]�<��8�� dťi0��i �������������i0���i ��������  ɼ���a�1�]�-�D dŢ���ȑ�� ��� ��i0��i ���ߩ��� ���_��a�Ș B����a�����`��`�����`���M�]�I��8�� dťi��i ��i0��i �������������i0���i �������� ɼ���a�1�]�-�D dŢ�ȱ����'��� ��i0��i ���ߩ�����a�����`��`



}������i ��J��� dŹ��e��i ������` � � ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �ɍ& ���  ��� � � � � � �� � �( ���򩠅��� [ũ@�d�� �������`��������� 0ĥs)��������)�S����L������������� ��������� ������i ���L��@@@@@@8  0@P`8@@@@@@p�����Т ���	��8��������p����	��i��������������i����ɀ�LV�ds�sɴ��  ����  ����`

��h����i����j����k���������i����������i����� ��������`	
+,)*78'(56%&34#$12!"/0 -.                   P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������s)����`����������0'� �����������������Z ��z�����۠ �������������������Z ��z�����ة ��`��������������������� dŭ�JJe��i ����



e��i ��JJJJe���)�������������
.�.�
.�.����Q�ȭ�Q�ȭ�Q��i0��i ��i��i ����L��`es�s��`� �����`H)��ŅhJJJJ�
ei@}�Ņ` 0`��� P���@p��      Hژ��,
�h� h�`�;�<� �;H
���ōg��ōh� ����
`lg�����Ţ �;� �����`� �;� �����`� �;�( ��������;`� ��� ���)�� ���E� ����"�� � � �( ����`d 'Ƣ!�E�����(����` mƥ��`�(t���!����L'Ɯ��'�(� � �'���������,� �)�
����/�0�1�`��`�/��L�����0��0�`� �/�1m��0�,�
�)�	�)�� L�Ƚɪ��%� �&�/� �%0LX����L[����Lt����� �,����� ɱ%�1m��0 �L����� ɱ%��%8��%�&� �&L�����L{����������}ɨ���%���& �L�����- ɱ%H ɱ%H��}ɨ�%���&������h�&h�%L�����' ɤ/�ɠ �%�������%i�%� e&�&�/L����� ɱ%Hȱ%�&h�%L�����2�ɹ)��:�� �� ��%���ɦ/�)L�� � �L������/��)��)��� ɦ/L��ɀ�(逼�

���ə��ə��ə��ə ɦ/L�Ƥ/�
��ɨ�Rɝ ��ɝ �� ��  ɠ �%���ɦ/�) ɥ/
��%��&� �/��
��
��`�.��+��+�L�Ƞ �#���� �.L����� $ɱ#��#8��#�$� �$L��

� $ɱ#���Ʌ+ $ɽ�ɍ( ��ɍ) ���)�* 	�* L��   �%��&`�#��$`H���
�hJH��m�hnn���`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   ��C���  <				



				�0      �				



				

		��  4            
  
  
  

  
  
  
            0                  
  
  
  

  
  
  
            ���̽�����  ���  6���������  <���  &0 ���9�N�� �  <  
 	  ���  0 0���=�>� 8�=H� �>�h`H�=E=�=�I�i�hI�i ��$=� 8�EH� �F�h`H���E
�FhJH��eF�FhfFfE��E�F`�>EBH$>� 8�=�=� �>�>$B� 8�A�A� �B�B ��h� 8�E�E� �F�F� �G�G� �H�H`� �H�G�E���FF>f=��GeA�G�HeB�HfHfGfFfE��`�=�>E>�>I�i��=I�i B�(I�i`�=�>� �H=�*�>��>�h*��`�>EAH�AI�i�A$>� 8�=�=� �>�> ��h� 8�E�E� �F�F`��EJ�F�?=&>&?�?8�A��?&E&F��`�@EBH$B� 8�A�A� �B�B$@� 8�=�=� �>�>� �?�?� �@�@ �h� 8�E�E� �F�F� �G�G� �H�H`��EJ�F�G�H�C�D=&>&?&@&C&D�C8�A��D�B��C�D&E&F&G&H��`���Eϐ��EϘ` 	$1@Qdy����=�>��A��B�F�E�=&>&E&F=&>&E&F8�E�A��F�B��F�E��**EA*�A&B���FBjFBj`��8��
��i
�=�



=`�=�>��=��ϥ>��ϐ
�>�=��υ=8&E&F���E�F`    
  ( P d � � ���@�E�=�(Х>�)Х?�*А�?�=�(Ѕ=�>�)Ѕ>8&E&F&G����`        
    (  P  d  �  �   � � � @ '  N @� �8��@� 5�I \хA�I WхB�N�A `ͅg�h�MH�B `�8�g�g��hg*�M�N�B `ͅg�hh�A `�eg�g�ehg*�N`�J \хA�J WхB�L�A `ͅg�h�NH�B `�8�g�g��hg*�N�L�B `ͅg�hh�A `�eg�g�ehg*�L`�K \хA�K WхB�M�A `ͅg�h�LH�B `�8�g�g��hg*�L�M�B `ͅg�hh�A `�eg�g�ehg*�M`I�8i@�@�!���"

JJ(�I�i )?����(�I�i � `�� `����` 	"%(+.0369<?ADGILNQSUXZ\^`bdfhjlmoprsuvwxyz{||}~~8�S�O�W�T�P�X8�U�Q�Y�V�R�Z� �[�\�]�^�\�h�[FhjFhjFhjeO�S�\)�heP�T�^�h�]FhjFhjFhjeQ�U�^)�heR�VLpҥ\�h�[FhjFhjFhjFhjeO�S�\)�heP�T�^�h�]FhjFhjFhjFhjeQ�U�^)�heR�V�We[�[�Xe\�\�Ye]�]�Ze^�^`�)�A�JJJJ�B�i)


8�A�=�i)�J8�B�>�j)


�?�j)�J�@�ge=fE8�o�jEE.�=e?8�A�E�E� �he>fE8�p�jEE�>e@8�B�E�E�8``H�ZE����e����充��  E��� �� %��s��tz�h@��+� �� �����m���� � � � �`
�
m�� �qә������`�,
� � 8� � 
�@@ 
��<� ( �  �S����l��@�?�  �����  � � � � � � � � � � � �	�& ���d��<���x�����,�h����멀� �q
������p���L[Ʃ �u�@�v�����CԠ'�u���0eu�u� ev�v��� �������	�����` U���p


 ]ԥo
ey�y� ez�z`dz
&z
&z
&z
&z�y�z
&zey�y�ez�z�@ez�z`H� ��hHJJJJ ��h)	0�:���H�Z�uZ�vZ ��z�vz�uz�h`8� dv
&v
&v
&viZ�u��ev�v� Z�u�i �Ԡ�y �Ԡ �y�0ey�y� ez�zz����8�y�~�y�z��z`���Z؅g���Z؅hFi�	Fh*Fh*L �Fg*Fg*Fi�	Fh*Fh*L3�Fg*Fg*Fi�	Fh*Fh*LF�Fg*Fg*Fi�	Fh*Fh*LY�Fg*Fg*`        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l���  �U� h� �� :�`�; q���`�i`��)�J�udv
&v
&veu�u��v�yJJJeu�u��v�qeu�u�
ev�v�i�y)�Ȅg����)�Ȅh� �@u�u��g���eu�u��v�h��`dodp GԢ �_�q
��� �� ������q���	 �� �������`�ey�y� ez�z�_�_I��_�Xey�y�ez�z`�; C���`�i`����e}�i�-e~�j�i�k���l�� ]ԽyJJey�_� ez�`�_�y�`�z ���ei�i��j��e_�_�e`�`�l��`� Z�i i��ey�y��zz��k��`��)�J�JJ�o��udv
&v
&veu�u��v�yJJJ�peu�u��v�qeu�w�
ev�x�{eu�m�{ev�n�i�y)�Ȅg����)�Ȅh GԠ �@w�wZ�m ��z�y�y��z��g���g�gey�y��z�eu�u��v�em�m��n�hк`dv
&v
&v
&v
&v�ue�w��ev�x�}eu�u�~ev�v��eu�u�ev�v� �u�g�w� 1yg�y��u�g�w�1yg�y��u�g�w�01yg�y��u�g�w�11yg�y��u�g�w�`1yg�y��u�g�w�a1yg�y��u�g�w��1yg�y��u�g�w��1yg�y��u�g�w��1yg�y�	�u�g�w��1yg�y�
�u�g�w��1yg�y��u�g�w��1yg�y�z��u�g�w� 1yg�y��u�g�w�!1yg�y��u�g�w�P1yg�y��u�g�w�Q1yg�y�z`�i����o�y�p���u���v�-`�<���x�����,�h�����`L���p GԠ �u�����u��v������� ��L��`�g�h�ue{�w�ve|�x�yH�zH �h�zh�z`�zH�yH�g� Z�w ���ey�y��zz����hi��yhi�z�ew�w��x�h��`dodp� Z�{�� ��z���Z�|�{��	�| ��z�����`H G��o�oI��o�phdvi��v
&v
&v
&v
&ve{�u�|ev�v� �u� �y��u��y��u�0�y��u�1�y��u�`�y��u�a�y��u���y��u���y��u���y�	�u���y�
�u��y��u��y�z��u� �y��u�!�y��u�P�y��u�Q�y�z`�s�s��`�s���s��`�sEtM  e�*��E���e���&�E���`u�g�w� 1yg�y��u�g�w�!1yg�y��u�g�w�P1yg�y��u�g�w�Q1yg�y�z`�i����o�y�p���u���v�-`�<���x�����,�h�����`L���p GԠ �u�����u��v������� ��L��`�g�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                .                    �Kw�    ..                   �Kw      PCTOOLS EXE           ss9��� AT86    COM           �^�K�  AFC     EXE           c�`��  256     COM           P�f�  DS      EXE           @�ok$Y  SPEED   COM            `a�!A  XDEL    EXE            (���)  TREE    COM            (���%  HEXOBJ  EXE           [L���"  POPDROP COM           �Z��?"  POPPRO  COM           [Z��O  TY      EXE            hA�  SETUP   COM            !��  PRCOLOR EXE           ;W��Ґ���