@<  ��1 �� � � ��� �� � �   ��   � � � �� �   ��� �	� � � �   ��    �� ��	  �  � �  �  �   �� �   �  � ��	 � � � ��� �� �      �	 �� �
 ���   ��  �
 � � �� �
��   � �� �� �  � �� ��  �  �    ��  �   � �� ��  �  � �� ��  �� �
�
 �   �� �  �	�
 � �� �� ��	 �   �	�  � ��
 �  ��    �� �         �  � �
 �� �� �   �    �     � ��
 � �� � � �    � �	�
 � �� �
� �
 �  � � �  � �� � �	   �  �� � � ��    �� � � �  ��	 �   �� �� �  �� � � �   ��   � �� ���  ��    � �   ��  �� ��� �
� � � �
 � � ��� � � � �$ ��� �L �� �� �� �� �� �� �? � �� � �	 �� � �� �� �� � �� �� �� ��
 �� ��� �	 � �� �� � ��� �	 � � �� �   ��� �	 � �     � �� �� �	 � � �� �� �� �	  �� �� �� �� �� �� �� � � � ��� � �
�	 ��    ��	 � � ��� � �	� ��
 �� �  �	�� �
�    � � ��	 �	 � ��� � �� �� ��       �� �� �� �	 �� �	� �� �   �� � ��	    �      ��� �     � � � �	   � � �� �     �� �    �	   �    ��  �     ��
 � � �	   � � ��   �       ��	 � � �	   � ���       �    �� �    �	       ��� �    � � �� � � �	   �� �� �  � � �� � �� �	  �� ��� � �	 � � � � �	 ��  �� �	 � �� � �	 ��    ��� �	 � �� � � �� � ��� � �� � � � �� � ��� �	 �� �	 � �� � �	 ��� �
 � � �� � �	�� � � � ��� �! �� �� �!�!�!"!""#B"%b"'�")�"+                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                @<  ��2 � � � � � �� �� ��  � � � �� �   �   �
 �  � � � �� �   ��	 � �� �� �    ���  �
� �  �� �     �
 � �� �� �     �     �  �	 �� � ��� � � ��    �	 �
  �	 �   ��� �      ��
     � �
     � �   ��� �� ��
 � ��    �   � �   ��� � �  � �   ��	 �	   � �    ��   � �      �
 �    �   �   ��       ��      ��       ��    � ���      �   � ��     ��    � ��� � � �	     �	    �� � � ��  �   � ��  � �
� � ��       �
 � ��	 �  � �    ��       � �	   � �� � ���       �   ��  ��
 � �� � ��� �  �  � � �� �  �� � �� �   �  � � �  �  �    ��
 � �� �	 �� � � � � � �� � �� �
 �� � � �� �   �� � �� � � � �� �� � �� � � �� �� �� �� �� �� �� �~ �� �? ��9 � �� � � �� �� �� � � �� � ��� � � � �    ��  �
 � �� �  �	�� �� �� � �	  ��� �� �� � ��
 �	� �� � �	 � �
� � �    �� � �� � ��   � �	�� �
   � �
�   � �	�� �	� �   � �
   �� �	� �� ��
 � � �� �� �� �� �� �� �	 �� �� �   ��� �	� �� � � � �� ��� �   � �� �   � � �   �� � � ��  ��    �  ���    � � �� � � ��� �� �� �� � � �� �     � �� � �   ��� � � ��   �� ��� � �	 � � � � � ��     � �    �� �  �    ��    �� � � �� � � �	� �� �	� �� � �� � � � �� ��	 ��
 ��	 �� � � �
 �� �� �� �� �� � � �
 �� � �� �� �
�  �� �� ��� �� �� �	�    �� ��� �� � �� � ��� �: �� ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ��� � � ��� � � � �)��� ȩ)����� � ������i��i ���� ���e � ���������	 ȥ )��������)�S����L������������� ��������� ������i ���Lƀ@@@@@@8  0@P`8@@@@@@p�����Т �*�	�,8��,�����p��*�	�,i�,���������i����ɀ�L]�d � ɴ�
������`

��h��*�i��.�j��2�k��6���)�-i�1�5���,�4i�0�8� �+�/�3�7`	
+,)*78'(56%&34#$12!"/0 -.                     � �              �     D3�L0�L3@� 1DD33DD            � 1@L�03D1���1 D 1��0�1� 1  � 1�@  D 1� 1� 1�D13@���3 D3��03��13�L13D3�3D    D 1�13��13��13@D 3@L 3@L3�L33 �  �           �          �  @    ��L 3�1�1� ��0� 1� 1� �1���� 1� 0�L3@�   �0�3L  �D1� 1� 1� ������13�L13��13���    D3���13��1� 1� �L33�L33�L03�L          ��           �    @�03�03�� 3 ��L           @  � 3��L���� @�3�L0� 1�  L 3�0�  � 1� 1� 1������ @�03��13�L13���3�    D�1�L13��13�� @L 3@L3DL3�L     �   �        �          0 �      DD13DD3 � 3�0�3D 03�D1� 1� 1D 3���@1� 1�0�� 1 D  @�1�   1� 1� 1� 1D ���@13��13�L13��13DD3D    �3D13��1�@1� 1D 33�L33�L13�L3@D� ��@���������`�����[������d ��� ������ �� Y������������ i<� ��`

�� ���� � �����`� �/ ������`������@�]�<��8�� �ǥi0��i �������������i0���i ��������  	����a�1�]�-�D �Ǣ���ȑ�� ��� ��i0��i ���ߩ��� ���_��a�Ș �����a�����`��`�����`���M�]�I��8�� �ǥi��i ��i0��i �������������i0���i �������� 	����a�1�]�-�D �Ǣ�ȱ����'��� ��i0��i ���ߩ�����a�����`��`



}:���;�i ��J��� �ǹ>�e��i ������`@�@� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  @<  ��/ ��% � � ��� �� � �� � �� �� �� ��    �� � �� �   � ��    �� � ��      �� �� �   � �� �� �    ��	   �� �   � �� �� �  �� �� ��   � ��	 ��  �� ��	    �      � �� � ���  � �
 � �� �    ��	 �� �	�� �� �� �     �� �  ��� �  �� �      �     �� �  �   �	      �� �� �� �� �� �� �    �� � �  � �	 �� �� �    � � �   � �� �� �      � �      � �� �� �    ��    �	  ��
 �	� �� �       �   �     �    � �� �        �    � �    � �� �   ��   � ��
 �� �� � �� �    ��	 �� �� � �
 � �    ��	 �	 �� � �    � �� �� �+ �	 �� �� �7 �� �� �� �� �� �� �� �F �! � �� �� �	 � �� �� � �� �� � � �� � � ��� �� �    � � ��� �� ��    � �   � ���    � ��  �� �   � ��   � �� �
� �  ��   �	 � � �
� � ���   �	 �	� �   � � ���      �� ��    � � ���        � �� �	� ���        �  � ��   ��  �   �� � � �      ���           � � � � �	�� �         �  ��  ��� �  �� �� �    �� � �� �	� ��   �� �
 �� � �  � ��� �	 �� � ��      ��� �   � �� � � �� �       � ��    � �   �� � � � �� �	  � � � ��� � � � �   ��    � �   ���    � � �   � � � � �� � � �� � �� � �� �
  � � �� �    ��� �
 �� �
 �� ��� � �� � �� �� �� � �� � �� � � � � �� �? �� **+�z-***�+�.�%-�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	
           !"#$%&'(    )*+,-./0123456               78     9::::::::::::::;   <=>    ?@ AB        CDEFGHIJKLMNOPQRST  UVWXYZ[\]^_`abcdef       gh                                                                                                                                                                                            ������W���	�	��������UU��    ��������պz�`�`��	�	�	�	�	�	�	�	          P��             @ �         } �             @�             PP�           UU���                                           `�`�`�`�`�`�`�`�         @ � �       T�����������_��������@������� �     U�� � �     �������               ��   �����������U_��������U����?����          � ��������      _ �T������_�����?����������������   @ �P��� � � � @��������            �     ��������}����\U����������_������ ���  @�T����?? T�������� �@U����?�            � � �        ����?�� | �  �?������� ��    �   � ����    � � �            ����  ��  ��� ��W�����W���������������� ����     �    U���� � � � �T�����             �   � �   �  ( �"�(� �  ���W�����    ��UU��������    z�պ��������                 P �            @�                          TU��           e �           @ � �          U�e�j � � � � � � � �j���Zj����j     @��j�        U@������        E��j��       U@������F      A��j j �����Z����Z����e  Aj��Zj        P��� �@�@�@�@� � � P�jAiZ �A�F����    T ���E�Z�Z        jj�j�j      P��j��*�       U@�������     T �A�F�����            � � � � � � P  �_����@   �������T  ������������EA  ������T  �G�������W�����UT�_�UW������_����P  _GA�@� � � P  �����     @_@�@�@� A  ������U   �E�A�G�_�_�_@  U@@@     ���U�����P  �����W�_��@� U  _������@           �W����@U        �               	
                               !"#$%     &'()*()+,-./01234*3456789:;<=>?6?6?6?6?6?6?6?6?OPPPPPPPPPPPPPPPPPPQPRRRRRRRRRRRRRRRRRRPSTPUUUUUUUUUUUUUUUUUUPPPPPPPPPPPPPPPPPPPPP�j����������ZT�0��3�3���0���������� � 0��<?���� 0 ������<��� �            �?���< � 0��? � � �������0������� � � � �� ������������ ������ ����� ����� < <�� � � �ꪺ��������ZT              UU��30�0 33��UU?��   �?�UU�000�030�UU�?3 3 �0 0 �?UU              U�� �  �   ?33?����  �����������  �     ?? ?  �                          UU �            UU?��UU�?3�3��?3 3 0 UU�?����]�eYUU�P�j��VU��& & %�$��j��UU��    <�j��UU�� � � ���j��UU��     0�j��UU�� ��3����j��UU��?   � ��j��UU��  ��� �j��U��� � � X������������ZT�������������VU��f�f�f���TU  U���U�i�Y��U  ����������      &?�?��&�&�$?�?���<��0�000��� �<0���� ��� ?�    �  �� ?0��3�������� 0  0�?�0�? 0 < ��?��?�  0 �?�<���?ZU�j�e�i�U��PU  U���V���f��U  �����������[�j�[��������$$ ��TU        �  ��UU        0   ��UU        ��  ��UU        �  ��UU        ?   ��UU        ��  ��UU         �U        �j�[�j�[�j�[�j�[UU������������UUTU������������TUPU������������PU@U������������@U U � � � � � � U T � � � � � � T P � � � � � � P @ � � � � � � @U�*�?�?�?�?�*UU�
�����
UU������UU � � � � � � U  * ? ? ? ? *   
     
          �QU����  ������  QU����  �������jQU����  ������  QU����        ��* *�*<*�*<* ���V ��0�� � ��V          ����������������������������� � � � ������ � � � � ������?���� ������ � � � � �����������?������������??<<����� � � � � �����������?�  ��������������������?�     �������������������?�?�?���������0        �� � � � � � � � �    �     � � � � � ��� � ������������          �  � � � � � � � ����������?�               ���������������������?   ?���             ����������������� ? ? ? ?�?���� � � ����?��� � ? ? ?�� ��  � ������� ��? ? ? ?�������     ���������� � ����?�?����������������� � ����?�?�� ��?���?���?           ��� ������� � � ���?����?�?�?�������?        ?��� ��� � � � � ������������������?�� ? ? ? ?     ������������ � ��������������?����������� � � ���������������������� ? ? ?   �������������������?����������  0      �      � � �������<  ? �  � � � � � � � ��� � ������                  � � �  � 0��������������?���?�?��������������������������������������  �������?��?  �         ������ � � � � � � ��  ��������������? � ������� � � ����������������  ����          ���������� � �������������?�?�?�?����������  ��������������������������  ���?���<   � ��              ���������� <   ������������������?����          ������������������������ � � ? ���������� � � ���?���� � � ��������     �������0?�<    �������� �  ������������� ? ����������������������� � � �                ������ � � �������?       <              ���������������������?���                 � �������������3 � ���?�?����� � �           � � � � � � � ���������?�0  ? ?  ?         ���������� � � ���������            ����������� � ����������?�����                ����������������     ������ � � � � ��� � � �����������         ? �? ����������������? ?    ? � � � �       ?�   03<���?�?�            0 �� � � � � � � � ���?��?�?�?�?����� � � � � � ���� � � � � ? ?�����?������������   ���������������?�������?  ? ? ��������������������������?  �����������������?���� � ?0 � � � � � �    �?�?�?�� ? � �? � � � � � �   ��?��� ? 0? <    � � � � ����������������������?�� ?  ?�� �       � ���� ������������������?�?��� �� � < 0       3 ���������������������������?�?��? ? � � < 0     �����������������������?�������?����������  ����������������?�?�����?�   0 � ��<��������������?������?�?�?��� �� � �  � �<������������?�� � � �� �<���?�? �������������       ? ����?����������������?<    �� ���������������������������������  3 <     �������������� � ��?�?�  ������          ���������� � ����������������   ����������0� � ������    ��������0� � � ��������?  �������� � � � ����?����?� ���� � � ��� � ������������    ��� ���0    ����������������   ? ��� �  � � � � � � � �  ? ��� � ?  � � � � � � � � ? � ���� ?  � � � � � � � �    � ���?�� � � � � � � � �� ��?����������             ��������������������������?�����������������������������������������?���?����������  �  ����������������������  ����� ? ? ? � ��� �� � � � � ���? ? ? � ��� ����0� ��� �� ���?    ? � ��  �0�� ��� �� ����������? ���0� � � � � ��?�?�?�?��������          �������������������3�3��     ��              �������� �    ������3�3�    �  �            �������� � �  �          ������� ? ? ? ? ? � ? ��������������������������<� � �� ? ? ? ? ? � ? ������������������������������� ��� � � � � �����?�?�?�?�?��? � � � � � � � ����?�?�?�?�?���?? 3      ? ?  ������������ �0�3      ? ? ?   � � � ������� �0      � � � ? ������ � � � � ������ <     � � � � � � � �?0� � ��������? � � �          �?�?����?���?������������?�?��������������������������������������� ����  <�?�?�?������� � ��?�����  <?�?�?���0�������������? ? � � � ����������� ���������� ������������� �  0�?�� ?����?�?������������ � � �   �������?�?�����������������   ��� � �         ������������ �0���                     � � w U u W    ? � ��W�      � � �<T��T    ? � �u]V          ���         ��@\C\C    ���?U7�e5          �?����                   �?����Tu�]TV               � � �        ���uUe�W]�w � �� _U}Wu_� \p\�\U\��] wPꥪ� U}W� / �� � � �        q=vU�U�ׯz��� �g�U5�5]U �         � _pU\UTu�]TVp��UUU���       5 5      |�UpUp��  p��UUU���_UpU��    5 5     �@�@���:�/ �?���
�
�
�@�/ � �@�@�@: � P �����
�
� � P@����}�      �����T         ���*�*�:�@�/ �              ���*�*�:�@�/\��  @ � � @   �WU���������  �    k ��: >�   @ @ @       ������������  �  j ����� � >               � � ����]@U��_gUm  ? ?  5]W5             � p          � ��               �     � ����]@U��      ? ?  5 p p �          U��U���������� ����֪4� � /  ? �P\P\Sp�p]pU�� w�wYY�5U5�5] \ W � <   � ���Ugeg_�XU�V�����]W5U��5��5
          �   @ �        �P
��                       ��T)h     @ � �������ꩪ����:    U ������ ��>< 0         ���@� � �      j j k          � � � ��T�PT  
�:�ꫪ�����UU     
 ZV         \ @ @ @ @      %XPPP��      5               ��TT � � � �A�U�U  �����ꫪ���      jAWUU                 @  � ����������  
               � � � �@�       ? �  �   @ ���
��m       �?���t�U�     J�:��Ѻ�n    �����Ъ             ���                   p \ W W W T�����_�U�U�V�[�  = � � � 5 
  � ���p�\�\��\�����_�VUVUZUjU��*               � p \\���������_�W�UWU^�����     * �� � � \ � �    ��
�i}u��WW]|�� �_	W	U	U	U�
        @�I�vh�@���P�@�w���kߪ{  ? ? ? � � �  � � � � � � P W�������� p   * k �  %  � � � � �     p���������WW�[
        5 ��誥�T���     �*�.�;���PW�� � �          ��ﮩ��䮀� T��:            ����Ъ������pW	�*��{�j�����p��z�ʌ� � � � � p�mU��������Ū% � � �����V �   � � @ � @ �    ����U � �   ����U ���� P  	@� $ 	 :     ������p�P`-       P $ 	@      ���p��]@V                      ���p�              @ � � � � j��p�������-Uު� @ � � � ��y � ������
��ת> @ � � ���J\��A�b���.��U�
                   �ppV�\UPU�+��+����Z%� ' � =               � �   ��* � �����髫��^̫        
            � �  �]@V � �����髫�                 �       @      :�T)h%X�V              �� @ P P P P @ ��j��VYQA5
     ` @      � � @ P P V X ��Ua�u5A% 	  P P T T P � �  �
�uQ]B �:@U h            ���jZU`U�U  �:               �C��UdUTUd%U�(
 
            � )�)         ���WC�P��U�UT�  
 
 
   ��  @ @j����      UUUUUU����        ��
         � | t T8P�T�U   = 1  �U	Y$ � | t T8P�T�U�o = 1  �U	Y$V!   � | t T X�W�{   = 1 �U	Y$Y!   � � p P @ h�V  ? � } �  �U	          �*���U  �w=�1dX�feUY           	 $ �o�_�_�� t � � �V!U%Y
�� � ���_�_�� t � � m�YU%Y
�� � ������� � � t � ��mV%U%Y
�� � ���U��<Z P p � � `U$U!f�&U	���*<Z ` �          �Z�W���iPW��ꪵV! % 	     
          � � ` P        �
�%X%X          	             @   �          ꫨ*�V                    �PT)h%X f�e���� V X � �UU	U	VV� ��Y�Y�Y f � � �  E� U� �  �Y`V`V`V�Y � � �E� � U� � P X X X X `   @U*E�U��
�: � � � �        �U�U�UUVUVVQ����) 4 $ %  	     H H X8Y~eU<TT�V�V�V�V�Z���k$ ! ! % e,Y�U�< `  H H Yxe~U?T�VT�V�V�V�Z���j	  ! ! e Y-U���VUUUU����       �����@����� j��    
 
  6 :     
 
 � vz �����@����� j��    
 
 " * :              < �  ����*�*�
�   � � @�� `�� ���
�
�"j*�:   � � @ � �   ��ꌾ�������뀪�� * *  
 ; � �L�����������������  * ; � O����ꬾ � � �@�: : ; � � � � �  ' � �����ꨪ����+�*�*����*�O � � �       @�:�:�;�������� @ � � � 5@� $@           P @ �          \
h�                         ��9��亨���@@   
 j ���  ��讨����@@   � 
  * * � P  ��@� � � i X   / 
 * �        � �            �:���ʰ�* �@   � @            �/�
�*��iX   � @             � � ��7��Ꜩ  :�*�:�ꪪ�����     +7�5�  ������ ڰ� �)��� � 2� 豩����������Ѕ����������\��[������ &� .�� �� �� W� k��s�� ���Z � � B� ȯ �� 8� z� O� � �� � s� <� ��]��]L��``�@�e��] ���
�������dpdq� ���`���`���`���@�����dodcdd���f�<��g�=��h�[�:)
��>��i�?��j� �g�kȱg�l� �i�mȱi�n`@GFEDCBANMLKJIH�@��� ��dX���� ��X��� ��8��Y��� ���$X����Y���$X�	���� ���$X������L���e � �� ����P�����`�� ٰ ƥ )���P��`������Q�\�P�Q0�P�� ����Q�PLi����� Vå[ ��L��STAGE �� �)��� � 2í�����	������� �ĥ[ �ʪ)��JJJJ �ÊL��`���x�`����������x��`���?����B���������B���?������ Ví��'���&���%L��������`������`������`���������������� Ví��'���&���% �ʥ/ �å. �å-L��  �]
�����^����_��]����^`PRESS START BUTTON  Copyright 1993� Thin Chen Enter.���������� �� �ƩV�� �ϩ��������� �ĩ����ƅ��� �ĭ ��� �� Xӭ�� ��L2�dbd`da�@�������i����b���i����b���qk�Pȭ�iqk�Q���qm�Rȭ�iqm�S ���`�`�R8�Q��P8�S�f`�P�R��Q�R���`��a`�S�P����`��a`	
���������ȴ �������	
�����������
	�`�
������`�Z)���]�L���������� �Y�������� �X�������� �W����L������X�L������
�Բ���L���߲m���� m���� m����o�
`��o�LXƭ���`���Y�`����X�`����i���`��)���}�� ����c�o�`��o�LXƭ���`����W�`����
�����`� y��� � ��d��o�LXƭ �` �ϩ�� �Ϡ ��[� �)��� � 2â��Lۮ�e��e�o��o���` �ϩH�� �Ϡ$ ��\� �\� �)��� � 2â��LۮGAME OVER�� �)��� � 2é��	������� ���<e � ����P�� ƥ )��P����L���Y�$��g�Uȱg�V�	�i�Uȱi�V�Y�U��P�R�V��Q�S�i�R� eS�S� �$�� �T�$�����U����V�����U����V� �T �� ��<e � ���U��V��R��S�� �T �� ��e � ���U��V��P��Q�� �T �� ��e � ���U��V��R��S�� �T �� ��e � ���U��V��P��Q�� �T �� ��e � ��L�ϥo�`�e����� Fϭ������ �eLy�F�n�����¶޶���.�B�V�j�~�������η���
��2�F�R�^���r�����¸ָ����&�:�N�Z�f���z�����ʹ޹���.�B�V�b�n���������Һ�������"�6�B�N�v�b�������ƻڻ���*�>�J� �� �   � �� �   � �� �   � �� �   �   �)*+�123�   �    �+*)�321�   � � 	��#$%�      �	 ��%$#�      � ,-� 45�=>?�      �-, �54 �?>=�      �./0�678�@AB�       0/.�876�BA@�       � 
��&'(�       
 ��('&�       ��� !"�      ���"! �      � � � �      � � � �      �   �9:;�CDE�   � < �CDE�MNO�XYZ�ghi�      �MNO�XYZ�jkl�      �ONM�ZYX�ihg�      �ONM�ZYX�lkj�      �PQR�[\]�mn �      �RQP�]\[� nm�      � ST�^_`�opq�        TS �`_^�qpo�        UPQ�abc� rs�        QPU�cba�sr �         VW�def�tuv�       �WV �fed�vut�          �FGH�JKL�   � I �JKL�wx ��� ��� �      �wx ��� �����      � xw� ��� ���      � xw� �������      �wyz������� �       zyw����� ���       � {|������� �       |{ ����� ���       � }~���������       �~} ���������        ����������       �� ���������          ���������   � � ��ԥ� ��� ��� ���      � ��� ��� ���      ��� ��� ��� �      ��� ��� ��� �      � ��� ��� ���      
��� ��� ��� �      � ��� ��� ���      ��� ��� ��� �      �������������       �������������          ���������   ��������� ��� ��� ���      � ��� ��� ���      ��� ��� ��� �      ��� ��� ��� �      � ��� ��� ���      ��� ��� ��� �      � ��� ��� ���       �� ��� ��� �       � ��� ��� ���       �� ��� ��� �       � ��� ��� ���      ��� ��� ��� �      �   ���������   � � �����   ���������   � � ��ԥ� ��� ��� ���      � ��� ��� ���      ��� ��� ��� �      ��� ��� ��� �      � ��� ��� ���      
��� ��� ��� �      � ��� ��� ���      ��� ��� ��� �      �������������       �������������          ���������   ��������� ��� ��� ���      � ��� ��� ���      ��� ��� ��� �      ��� ��� ��� �      � ��� ��� ���      ��� ��� ��� �      � ��� ��� ���       �� ��� ��� �       � ��� ��� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l��� ���  � � � � � � � � � � � ��" ��d`� ��@����'� ����0e�� e����`�


 ní
e�� e�`d
&
&
&
&��
&e��e��@e�`H� ��hHJJJJ ��h)	0�:���H�Z�Z�Z ��z�z�z�h`8� d
&
&
&i ���e�� Z�� Ġ� Ġ ��0e�� e�z����8��~����`���č���čN�N*N*L9�N*N*N�N*N*LQ�N*N*N�N*N*Li�N*N*N�N*N*L��N*N*` �U�L��� Và ��������������� ��L��`

����� ���6����C����,0)�*��,��)��+����i�nL��ȩ �)�*�+�,L�ĭ��e�nL�Ĝ���������  I�� �
>��`�H�H�H�H� �� � � � � � � � � 	� 
� � � � � � � � � � � � � � � � � � � � � �Сh�h�h�h�`��e�E����&E�m `��L������ ����������� ���L�ŭ�`��� �	� �� ���`�	�+� �
� �����
m�
��� � � � �	`
�
m�� �sƙ
������	`  8� 8�P8X 6� 8��8 p8v�8 ���)����� �������i��i ��i��i ���ة)������ � #�����ɨ��`�Z��J�"�JJ����e"�#���i �$�H� �#hz��#�$�



e��i ��JJJJe�� �ǥm��� ��ȱ��i�� e��i0��i ���� �Ǭ$�#`�����0�� iɪ�骍�`H)���ǅhJJJJ�
ei@}�ǅ` 0`��� P���@p��      )AYq�����1Iay������@ � � �Z�	�)��
�*���+���,�L�)
��	�%�
�&��'��(Z ��z�)�	�*�
�+��,��+)*� ��z������Љ`�)�%�*�&�+�'�,�(�')i��')Ji� �0� d!�%�'m:H���!E � h �ǭ(JJe��i ��&�



e��i ��'J�jJJJe��()�#� � �,'p�����0�� �ڪ�������#�!........��߬ �Q����e ��e!��m ��i ���L�` @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��H��
���


�h �ƭ���`��8��
��i
�%�



%`�E�%� ˥&�˥'�ː�'�%� ˅%�&�˅&8&-&.&/����`        
    (  P  d  �  �   � � � @ '  N @� �8��@� 5N�h�r���  6$
    0��  #0�U��y�m����  9000000	0		00	00	00	000	00000000000000000000000000000000	00��  $								    �m���1�U���  <)� ( )�  0)���  $	0	0"00$ � $	0��\�(�����  
�o�����o���  00 0 0�  000�  00�  �  0 0 000�  �  0�  00000��  '
0
0
0
00	0	000
0
0000	0000
000	00	0000000	0	00	00
0
00
00	0�(��Hژ��?
�h�3h�2`�N�O� �NH
��ύ��ύ�� ���G`l��&�4Ϣ �N� �����`� �N� �����`� �N�( ��������N`� �1�Y� �1��)�� �+��� �+��"�� � � �( ����`d1 hϢ!���+���(�Y�1��` �ϥ1��`�t1���-�+��LhϜ+�:�;� � �:�2��������?� �<�G�,��B�C�D�1`�1�`�B��L�����C��C�`� �B�Dm+�C�?�
�<�	�<�� L�ѽVҪ�2�8�3�9�B� �80L�����L�����L������ �?����� ^ұ8�Dm+�C ^�L%���� ^ұ8�K�88�K�8�9� �9L%����L������,�,�,}ZҨ�/�8�0�9 ^�L%����- ^ұ8H ^ұ8H�,}ZҨ�8�/�9�0�,�,h�9h�8L%����' ^ҤB�RҠ �8�M������8i�8� e9�9�BL%���� ^ұ8Hȱ8�9h�8L%����2�RҹO)��O:�O� �P� ��8��ӦB�<L�� ^� ^�L%�����B�R�)��O)�O�O�O ^ҦBL%�ɀ�(逼R�

��әM�әN�әO�әP ^ҦBL%ФB�G��RҨ��ҝ ��ҝ �O� �P�  ^Ҡ �8��ӦB�< ^ҥB
��8�2�9�3�B��G��G��`�A��>��>�L�Ѡ �6���� �AL����� eұ6�W�68�W�6�7� �7L��

� eұ6��Ӆ> eҽ�ҍ( ��ҍ) ���)�* 	�* L��   �8��9`�6��7`H���K
�LhJH��mL�LhnLnK��L�K`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   � ���������  ��� ��٥��/���� 2à Z���Iw� z������� ��� ��L��`�������������_^FNNEzz#W4W2Yw� ��� Vé���ԅ ԩ
��� Vée��Յ ��L�ө(H� � Z� I�z�����e����������C��������`e����h:м`��� ���Jjj(**HJ~�~�~�~�J~�~�~�~�hJ~�~�~�~�J~�~�~�~��ж����`            x   �   ?�  ��   ��   �� ��� ��?� ��� aÁ� aÃ� aÃ� Ã� �Ç� ���� ���� ���  ��  ��� ��� ���  ?�  �   �        �   �  �               � ��������  0�                   p   | |  | >  ><>  <><  80  ?0  ? g�� ����� � |p 0w� 8�����~s�  s�  � 8��������g   w   �   �  ��` /�p x<x |x|~ <x|g <y�g�s�c��`��`� � �?  �   �   �    @      xH�Z� ��  � '� �ϥ� �	� � E��e��E*�z�hX@xH�Z,$ ,% z�hX@���؎	��H��H��H��H M�h��h��h��h�� 2� �ϩ � � ��	  � 0�  ��ύ& �
L�� 	
 !"$������ �%�6�K�`�n�n؇ؕح���������ٽ)�� )���^�`��`�]�Lڪ�c�L�۠�^�:�^`� ��J��F�]�
�	 �ֽL�׽�+� �� )�%� )��� )�����^� �� ��H�b��^�r �h�ٿ��
��`�]�
���ݜ�������
���օP��օQ�]lP � L٥Z)�`� )�� ٥]��`�`� �]�
�)�Lح��^8�ɂ�����^`�^iɂ����^`�L٦]�
���
�Lٽ
��?�
��@�^�Lٽ
��/�
�� �^�L٩��^�  �Lyة��^� ٥o�`��o�LXƩ��^� �Lyؽ
���
���^� �Lyؽ
��?�
���^��@�^� �Lyؽ
��/�
���^�� �^� �Lyة��^� ٥o�`��o� LXƩ��^� �L�ؤ]��r��s��^��芨�]�
�g�kȱg�l`�i�mȱi�n`�]
��k��l�� �^�ȱ^�ȱ^H��^zL���   �������]�
�`�)�Y�)��X��B� ��^���a٠ q^ɂ�*ک
���� ���� �^�@��� ��^������ �^��^�Y}cّ^�Z)��Y�dX�YX�]�
� �!�`��^� �]��@��b�I@�^�]�r � �`�d�L��dpdqdYdX��^�����Y�p������X�q���@�b�� ��^�s ٠�^�:�^L�ڭ�L�ڜ��



���b��� ۥf���q� ��)���d�`�L�ڭ)�L�ڭ�' ��JJ)����
�b�)��	�����^��ڪ��� �)	����ۅP�ۅQ�]lP 
����K�P�c�v�6�K�6�Kاۭۧۧ)�� ���d��	� ���Z��)�����^`�L٢ ٥o�`�"�o�LXƢ ٥o�`�"�o�LXƢ ٥o�`�"�o�LXƦ]�c��^�
� �^8�Lؠ �^iL�`�^������ �^��^�Y}cّ^�Z)��Y�dX�YX�]�
� �!�`��^� �]��@�  �  �b�I@�^�]�r �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �^8�ɂ�����^`�^iɂ����^`�L٦]�
���
�Lٽ
��?�
��@�^�Lٽ
��/�
�� �^�L٩��^�  �Lyة��^� ٥o�`��o�LXƩ��^� �Lyؽ
���
���^� �Lyؽ
��?�
���^��@�^� �Lyؽ
��/�
���^�� �^� �Lyة��^� ٥o�`��o� LXƩ��^� �L�ؤ]��r��s��^��芨�]�
�g�kȱg�l`�i�mȱi�n`�]
��k��l�� �^�ȱ^�ȱ^H��^zL���   �������]�
�`�)�Y�)��X��B� ��^���a٠ q^ɂ�*ک
���� ���� �^�@��� ��^������ �^��^�Y}cّ^�Z)��Y�dX�YX�]�
� �!�`���& Lp�-���a�