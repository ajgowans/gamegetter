$'0$�Z��)�0��;� ��z�`)H�;��M��h �z�`���������6HZZll��|���������� ��@�� � �,���8�@,���8�,���8�,���8���������`�0d���
��� �� ����� �� ����� �� ����� �� 䁈��������`�	��
��
���� �� ����� �� ����� �� ����� �� ���������`d���
��� i̲	) �� ����� i̲	) �� ����� i̲	) �� ����� i̲	) �� 䁈������Ь`�	��
��
���� i̲	) �� ����� i̲	) �� ���� i̲	) �� ����� i̲	) �� �������Ь`�Z�
� ������z�`H� ��Jh� � �J��J��JJ�
JJJ��J������ �Ϊ�D��H������ � �e� �e� �`�    ��� � � i̲	)�&� ���L�����e� ��� � �� L����`� ��H� � �h ���`��� <��FLD�)���т��:�]�p�Ӄ�   @S��   @SEO��   @Scepn�
�   @S%%ENN
-	���   @Scgpl��   @S��   @Sb&h)l0QQ0
o
)h&e.	�R�0�0�!�!���   @Sbk
qh
'	�I�J���   @Sjie
	o

-	���   @S��HZ�
��Hυ!�Iυ"�ڲ!����Ȁ� � ����!��"���zh`HZ�
��Hυ!�Iυ"�ڲ!����Ȁ� � L���!��"���zh`� � ����`� ��`
����e����i ���લਅ���` ��l� H�Z� ����� ���� hHi�� � ��� z�h`d�����`x Ԅ��X` #�� � � � `� � � � `�@�� �� � �����������`��`�چ�
��W�-	�{�����s��i�� ���h��W�-	�^�����V�������)���C ΄�٦�}���I

�ڹ`�� ���� ��i� �� ⅊������	@�� �� 	@� ��0LP�`H� ����� ��d��)J��j)���� ��������J��j����"����e⨥�e㪀��e⨥�e㪊J��j�h`W�W�X�W�h�����ֆ��Ɔ`��
i� �� L����W�I�-	�	� � � #��� ��� ���( `�	)��	�� �� �� �( �`��i� ⅊������� `���������`��i� H ��� � ���  �����h`hLԄ����	 �� �( �* ���L��


�� ����� ���������t������ ������`Hک��� F���h` @��v
�F�F��o/�R"�ʢ|X7�����zdP=+����Ǽ������}voic]XSNJFB>:741.+)&$"                                       ���9 9 9 9 5 5 5 5 9 9 9 9 5 5 5 5 9@����@L@LEGGG@L@LEGHG@LLLEGGG@LLLEGHJL@��6��0�6���H��@�6��0�6���H��0�H���6��0�6���H��@�6��0�6���H��0�H���H��@��	��<7<7>7>7>7>7<7<79;<7<7>7>7>7>7<7< A<A<<7<7>7>7<7<<>@A<A<<7<7;7>7<7< ����HTQOHTQOGSQOGSQOGSQOGSQOHTQO@LOQHTQOHTQOGSQOGSQOGSQOGSQOHTQOHLOQHTQOHTVXHTQOHTQOGSQOGSQOHTQO@LOQHTQOTQVXHTQOHTQOMYXSLXVSHTXST��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� H��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� H��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� H��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� 6��� H��� H��� H����ЂC>>C>>C>C ��ЂOJLNOJLNOSO ��� 6��� H��� 6��� H��� 6��� H��� H�� ��$�����������0$�	0$�0$�0$��	��9@5@4@9@����9@@@> @A@@�� H��� H��� H��� H��� H��� H��� H��� H��� H��� H��� H��� H��� H��� H��� H��� H���H��@�H�� �H���H���H��@��������������������������������������������������������7�	7�7�7���0�	0�0�0�1��������i����!� 	� \ 'q 2!"4VDEh��h�ۻ��������������������������쇾�Ez�Fu  Q                            #42#VeVf��w����˽���������������˪��ۘ�������������������������������������������������������������̻��������˻�̻�����������ffvUDC332                          "#324D3DUUUVfgffwwgxwwwx�ww�ww��wwwwwwwwvgwfgvffffgvgwwwwwwx����������������������������˻�������������wwffeUUTDD3333""""""""""""#333DDDDUUVffwwwx���������������������������������������������������������������˻�������������������wwwwwvfffffffUUUUUUUUUUUUUUTEUUTDDDDDDDDDDDDDDDDDEUUUUUUUUUUUUUUUUUUUUUUUUUeVfffffffffffffffffffgwwwwwwwwwwwwwx��������������������������������������������������������������������������������������������������������wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww��                ������������������������������������������������������������������������������������������������������������g�@�KV�������o���  �   `    ���(���������������@�0���P���������             �PJm�~���������������������ٶ�
p\_��I�P                       ?o�������������������o�u� b        # @(� @          8��������������������������W�B�a       ��<P�R����)"�?��Tf����������������������&�@              $ %Sl������̞��)�50F��X��������������������o�d��Q                @�n��������������������{猃z��4sWRfGA aEf����W�h���v�6Tc�8TFr$&eVTVGC�k���������������������eW2 0            E8GU>���������������z��G��X6=U4q6G�S�xF������G��5K�1b Q3B#5F�$�3xuh�W�EGu�������ܬ��������������ʗ�cU       4!��e�����x���ݚ���������}ּ��ic{e~�3f�uId�X�x�y{v~ۅz�gxw�y����W���ggGde#Ev%dGSTFggtifkhf����������������ۻ���8CfT3$1tTSTGBx%TJe�eewsw�V�xdytxY��������������������tFC3   10SWf����̻�쬺�ʌ����ewFg4r$"%2V2eGdh��z����̽�������ܺ����wVvT%TDER2D32UcU6cxww��y��������w�j��g�w��v������̬����������˪�v�44#       !DdXx�������������껩�v�WwfvdvFvVwgwy��y�j���xvvFwDfWuwV�v�x������̫�˻����G�WeT5DVDFefV�v�����۫�ܼ�ܺ�����xwvfVfwgewffwhvw�f�wx������g�wvh�x���������v�wehdVVeF�Wxv�y��˹���������ۛ��efD3       35Txx��������������ʺ���eeEcED5ETFvfvy����������xx�fuWUeUFfWfWww�y������ܽ��̺������gugeUFeFTTFffxw�x�����˼˻�����wuUUDD3B"""4CUUvx��������������̺���xeUUDB4"31#3DDTVUWvVwvgx��������������˻������x�wudUTDTDDUEfwhh�x���������������xxwgwgfgWgww���������������������������x�x��wfwfUVTTETEDUVffy���������̻�̻�����wvuVdUDDUUCUVVgx��������������y�wvwufefVeffgww�������������������wwfvgfffVfvfVfvww�wx���������������wvwwgwvwwwwxw�w�����������whvfEVUVeeVfwww���������˼������ufUTCDC3DDDDVff����������̻��������wffTeVEEUUUffw�����������������wwvffVeUeUUVUWgxx�����������������wvfeEDUDDDTUEUfvwx������̼�̼�����wfeTD332"#333DEffx�������������̻�����fUTD4333C4DEUVfgw�����������������wwwwvfffffgwww����������������wwwfffUUUUUUVVfffwx�����������������������wwfffffffffffffgwwwx���������������������                �X�����wwwww�wwwfUUg������eVx����vUUg����wvfy���vfg����C4X�˹�Dg����TUx�����eUfx��w�������wfffx���uEEg�������eTEW�����w��uFy���eDFzͺ�gx�vEh��vTV���vfx�wvh���wvx��x��TDFy������Uf���Vxv���x��dVwwgvvfw�����Eh��vx������uUx��vgvUW��vx��wFx�����e33H�����vy��UDX�˅4w����v3"5h�����few�y����Xww���eff��˔�ۨwez޸eh�uVxx����uffeUgx�ͨfVfV����fg��CV�ʇ�U4h��ʘ��fewwgx��fx�w����fUV�ܧEhx�fT5i�͸eeh���gfVX�ܤ %��˗x�CG���w�ݹvUi�v�w�v�w����eW����wxgg���DE����uDh����Dh�ˆUUX�̦Vgv�v�ef��ۖUT4Y���CDh���C$�ݓk̗w��y��Bj˪�dVuW����3E�ubk��bz��ˉd$����RG����B#|ۖ�DW��tV�˅ev15��˸d5X����x��x��fdTh̸vSEy��gvVj�؄EWg�gTgz��s"H��16���̦3Y���ʗefVw���Dg��x�fh��w��dz�ɗe!7�˘�ywT4���tE�������SVuey���w��͹efi�wefU�h���wwDh���S$e��d5���fh�̘"2W���u"2[ݺvUW���wC4�̹eF������cEB5|ڗ�����t5W����eVEdW��ey���wRl��A $|�Sy��fhvy�tWvY���B5�ۇVU���CBY��fUUh����3�������Vz��QE�˷x�xcDG��xdC"J���!Y�숈46���S���et6i��UW�˗w��3B#l��BY���2He4W���eBW���f5H���wz�yxeI���1"J�ݩx�vS"{��a3f���eE#K��0l즉�QZ�뇉�Dh��Uw���BE����4 ޺r4f�e|�y�B7�y���� ���i��Dk����1��}�tz���B����CW����44W��c8���˃%w�Di�܇Gz��|�g�eD"Z���a!z�ˇ4"jͬ�wvffd����aJ�܆I���1X�ۨh�gcW�ۘffgwyh�����wug����v���x���uVy��w�w���www����wwwwwww��x��������������������������������������������������������������vffg������wwx�����wwvx����vfg����vT25���ɅC3F���c ����sF���  ����SG���s  ����CY���Q  |����R #���� ����V9���R �����`����a �v�ɴ����l )۔��S+�l�� �x��d
�ڻ� ~�9ڠ��_˙�P  U��_�3��*�ֻ�  ��F��9yQx틘� i�~tB�T��j�0 l˓|�!jyB���fT  f��t�w0j�c��D4 ����Z�S��V˫�3!��sfK�3$�����vC2�߶b��dfy���feUUTBj��s"%���ff���fVfwveVw���eUfx��wwx��xvffwwwwwwx�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwxwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwxww��w�wxx�wwx�wwwwwwwwwwwwwwwwwww��x�x�wwwwww���������������wwwwwwwwxxxwxw���wwwxx���x���w�wwwwwwwwwwwwwwww�x���x���w�xx�wxw�wxwwwwwwwwwwwwx������������������������xxx�xxww�x����������U��Jć%h׳u�Le|gwH��=�eDV���x�uG���vVf�g��w�wveWy��wy��w��wwxwgwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww                )����wfeVfgwx����������������weT3""3EVx���������˻������fT2    5x�����������ܺ��vUC"       #G�����������ܺ�vUC!        $V�����������˨weTD3332#2""""""334DVx����������ܻ��vUDD33333332333DDEUUUVw�����������˩�weUDDD33334DDEUUfffffvfffgx����������̻���feUDDDC4DDEUVffgwwwwwwfffffx����������˺����wfeUUUUUUUUfffgwwwwwwwwwvfffffgw���������˻����wvfUUUUVfffwwwwx�x���wwwwwwwwwwwwwwwww�wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww                郈w�x��������������������x�geVUVffefgw����������wfvVefUeWg���˻��wVefe�h�w���ͪ�{��vDDVf�h��f�YgwVfVtDBCUW��������ݪ��xv�xv�Dd4�Xx�����{���z����6rs3E7ww��ww4S'T��{�~�ۯ��HbeV����ʦt21 3v�tu2�U{h����x�t�{������쪙fsevgfTd5wdT#5Td��uuU�EFg���̻�xwfWv��̭������zhjh�v$T%e�{�v�eDRduVwz����v6w�����ږ     6Y���ͼǨz{������ʉ5!  6X�������hiYuc41E(Ugv���G" 1W�������ʘc!"4GEVs�(UZW�z{�ݻ٩��z�uH&USdS%Duy��m�˛ث��YVwIT�2    19��������t         S/��������0         ��������         Z��������         �������0        
��������         ��������        �������         �������A        �������         ��������        �������        ��������         �������P         A�������          �������         V��������D        ��������w         %z�����Ys��˾���0        "5x�ʛ��vuVFSaA"34ETD5%TTE4S3B@!2B!24&5CB2345DS55DEDUTdeV4332CUVGUeefWFDDC%$#22##44DSTDDDDTEEEDDEEDTDDDDTdeUEFFfgVEUTdUUVUUVddE64RcTE5CcUGETdTE44CTEFUeUUEETUDDECTDDTdeUFEEDCTUVETUUVVfeefVVUUETTETUEUUUUUUUUFETTTTTUUUUVUUUETUDDEEVWVTTEEUTUVVffeUEDTeeUTTEUeVVeefffeUEEUdTDEEVeeUUUVVVVUUUDUUUVVevffeUVVUTTDDUUUUVeeefGUeeUUUUUUUUdUEDTdefVVUTUGGg���ywveTC31"222#$H����˾�ʆT        &�����۷��i�S       \����휉��B        3�������רVB         )������ޜ�tA        d���������vB       #Dx~��������U     3EGW��fgh������ɚxeC22355UefffefVeeWWw�����yx��wgedUEEEDUUUeefVVUefgwwwww�xxvvfVeeVefffeevggffuvgffeeVVeffffvwwhgvvgggfvfffffffgffggvvwggfvfffefffgfvffvvwwgvvgffvfggffffffffffffffgwwggggvffeffWfvvvwgggfvffffefggvvvwwggffffffvwgggwwvvvvffffggwwwwgwwvwggfffgggvwgggffgvwwwwgggffffffvwggwvvvffgfvwgvvvggwwwwwgvggfvvwwwvwvgfffggwwwwgwwgfvwggfwwfvvwggwwwggvwwwwwwwvwgfggfvwwggfvwgvwwggwwwgwwwwwwggww�������wfeTC223#2 T����ɩ����C       ������ff��ws"      ����������ƃ        ������Ǩ|�w0        ����������A         ���������t1          �������ۗD   !  &��������܇S@   $4DCRU99��ܿ������ɦeD"224DUfx���wfUfggw��yy����������wwwwwwwwwwwffffwwxx���xwwwwwwwwwwwwwwwwww���wwwwwwwwwwwwwwwwwwwwxx�wwwwxxwwwwwwwwwwww���wwwwwwwwwwwwwwwwwww�xxwww�wwwwwwwwwwwwwx��xwwxxwwwwwwwwwwwwwwxxxxwwwxxwwww�wwwwwwwwwwwwwwwwwwxxwwwwwwwwwxw�xx����w�wxw���wwww�w��x��������w��wwwwwwwwwwwxxx��xwww�wwwwwwxx�������xw�wxwwwwwxww�xxx��x����xxwwwwwx�wxxwxx���xxx��xxw��wxxw��xx����xx�������wwwwww��xxx���xxw�wwwww�wwwwwwx���������veT3!  ���������wUSv����uB  {�����ok�wC��}Jd`    ~�����m��GWwgEDB    �������廗�tDSSUU1    ������ٹ��u21"4EDC     �����������d3#4ETT4  ��������ʷ�E$!1CEFVv�xWTSC#$D�������˚xvtdU55Uf�����wwffffgwx��������������x��������x�����x�������wwwwww�����������w��xx���wwww�����������xxwww�xxw�w������������ww�����xx�����������������������������������������������������������ww������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������x��������xw�������������wwvffUUTCC9N�������wveEEv������vD  0Ǯ�����ɗSB4F������vB  ������ݬ�wS34Hy�����vC!   o�����ͺ��e43Dfgx����weSAG������˙wuTDDUfw������wfeUUUVw��������������wwxx���������wwwww������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������wwwwwffUUv���ۺ����wfefgw�������xUB  0���̝�ɺ�ucE5Tvhz���ܻ�vB Y�ﮫ�͜��U4BTFV������ɖc0   ŝ���ͽ�ʚVSD%4ehz���ݼ��tB  @ƞ���ͭ��zF3$5fy����ۻ�vdS3#"22d������                a�����������������������������������������������������������������������������������������������wwwww�����������TDUUVxw����vh��ܨu#DV����eDF�ެ��tC��w��p)���g�tEX���{� !��ۘu3d8͗W��`]�ۻ�dVC}��(�0G���ۨh�I��!�aa��Ψfye���*�1"|̞��F�G��Bݥ4C����sXv�Ȁܨ�Xu���4�|�W����3�i��d86߄`{���2����t`^�	ɚ� �8��S�� ݭ�` n��ˤ O�P��b Ά���0�� |������ o�p'�����o� �� �O�#����β �p-@��0W��i�0�V���h���� ~�`o��� ���ɷ�v	�O� 	�|��{P |fP���`���դ ���?� (P���i0 yhs�r�c���Ă��K�_�@'c���G Xz��W�egn���` w�zf��`����D 'x��{�g |���S 0wj�G��p	����0 'U�tkؘ ����" 0tJ�6������� &�B[������  @`+�%���o���p  D�"J��
����  00=�%��Q����` s�#Yj�?����  X m�6��'����@  ��Dv=������  � ��GC�.���� L�
�Ur?d����p � �eg�����   ���VpmJ����P  ��Fu�����d   �`=�hPz����0  ,��G������3  � ncx2k�����  M��G�&�����  5� }E�2o����@  l��gs7����� F��7vC�����  E{`'�wd=�����  g��GgT�����   Vh@G��u����`  frzWxi�����   fVV�w������   e@&kf�������   vCf�i������   TV{g������� �0h�z������  2 f�h������P�&i�������� 2' f�z������1r 6i�������P t6f�������� Q`Fi�������1� Fg�������r HRRBVz�������3�1U4%h�������S2YRDBg�پ���Ϥ4%�!US&y̋�̼�CSiR%e3w�Ƚڛ���F7�3WSGyڋܙ���EtxS6uDw�������ugH�DgTX�ٛˈ���Wu�TGuF��������ewh�UwUx��������gv�fhvW��������wwhvf�ex����y���wwwfhvh��������wwwvf�V�����y���wwwvxvh��������w�www�g�����x���xwwwxvy��������w�wwx�g���������xwww�w�����x���w�wwxwx����������www�w���������x�wwxwx����������wwx�x���������x�wx�w�����������ww��������������                a������������������������������������������������������������������������������������������������������������������������������������������wwwwww��������vgvUVfx���vg��˩dDDg���vVv��ʗwRF��ۅCEy���eVwcY��t#Cy���TVww�e��5d�ͻ�TW����t2&����U����UbGw�ؿ�5��͹Xt2Gv��ϦW��ͷ9�UEu���uW��ʂ8W�vu���Ew�˷AVjڈV�}�X�|̄f[׈(���J���C
�~�tz��md��0o��D@6o����a���@7��a��	���Y��I�_�ٟ�t ���_ �pP\t�%tS���� �"@�W�7������o��	��~�
�2����<�����P��p
�}��� }� I�� �3���� �w x� �'�͞�� u���Ia��W���k��� ,y`m�r[g���� yw 6��P�������t h��R�����1$tQ���7����740z�f:�����U Io�vz���'�a �o�w���� '0�Ϧ�����7 f  d�x�����`r  y;�x����#P@ �_������ &  	���x����" C {f��x���r0@�=��x���2 0�چ{���#  ��w���0  �G������#0   	�M�w����#   ]��i����3 ���vz����   ݘ�W����B   Z��Y����! �ۍ������!  �ʞe�����  i�ȻH����A  �ݸ�Z����   �ݚ������    J�ۊv����b  {�ٚG����#  #�͹�h����!  7�ܩ�y����0  %+�̘�{���"  Sn���v����  a���wW����2  (5���gj���10  h˟�e����  �>�ބv����#  ����Ui���Q2  \Qگ�7|���"  ���I����"  ���a�����  +�=������R  m`���	����0 ����N����  ���@�����   ;�������`   �po������   $� ��q_����  )���AϿ���  ]���5����p  u��?�e,����  ��P��d��׷ x���u�����  9z���h��zq"xz�M�xz���z@4��c��y�꽷�!DH��E�w������TZ��8�x����xrU�w�k���ۚ�yR6V�wu����Ɋ��3gh�wg�x������Ewz�wh�y�����tFw�vvy�������dWw�fw�����x��Tgx�gx�����x�vVw��w��������vg��wx�����w��vg��vx�����w�wfx��g������x�wfx��g������y�vg��vx�����w��wx��w������x��wx��w������x�ww���w��������ww���x�                ���)�  ��a�  ��E�F�  X�V�    ��    $�1�B�      ��  �#�    ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                     0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �q�r �� ��� � � � � � � � d�d��ߍ& `�q���D�r���(�}� ���v�w� �  ����� ������� �  ���}�}�x� ��报�Ņ� U��r���(��� �� ������� � � �  >�日�Œ�  �`�s�t�vȱt�wȱt�xȱt�yȱt�z)
�����{����|Ȅsd}d~�x� �"��t�u� �
�t� �d���ds��`������ȱ���ȱ���ȱ���ȱ���)
�����������Ȅ�d�d���� �� �r �� ���v�w� � ����� � `������ȱ���ȱ���ȱ���ȱ���)
�����������Ȅ�d�d���� �"���񒅁�񒅂� �
��� �d���膌d���`H�Z�y)?	@���y*��%����~�{��z)@��J�����Ȅ~�{����~�zd~��Š�� ��z�h`H�Z��)?	@����*��%����������)@��J�����Ȅ������Ƌ��d���š�� ��z�h`H�Z��)?	@����*��%����������)@��J�����Ȅ������Ƙ��d���� � ����z�h`� d�`� d�`�󒅎�����d����  � >����r` �� /2�   �

		�
	�    ��  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                �U�U�ݪ�U�U�����? ��(?�V���� ?�50ڰ�0�:��k��,683�+֜5�� ,�8���6\� ��5+�3�8,6�� �8,��'ڜ��5 l��ck� � 0 �?�觲|y�� �    0 � � kc��l�+>��m=�?     �88 >�:���   l2�༃��p
Ю �     �Оpj��� ,�,:  � ���:�>6�9$ � ���;�9��� ��
 6�9�  �0�w��7�4�    *"�"""      �"� "�      *(* *(      
"""""
"      
 
 
                                                                                                                                                   ����  ��                    (
�$�)�
��                                                                                                                                                                             ��                  �
�(�(�(�(�(�
  �H�����*  �
�( (�
� � �*  �
�( (�* (��
  �(�(�(�* ( ( (  �*� � �
 (�(�
  �
�(� �
�(�(�
  �*�( *�$�	��  �
�(�(�
�(�(�
  �
�(�(�* (�(�
                                                                                  �

( (�
�  �                  �
�(�(�*�*�(�(  �
�(�(�
�(�(�
  �
�(� � � �(�
  �
�(�(�(�(�(�
  �*� � �
� � �*  �*� � �
� � �   �
�(� �(�(�(�"  �(�(�(�*�(�(�(  �*H�����*  �* ( ( ( (�(�
  �(�(�
��
�(�(  � � � � � � �*  �(�*�**"* * *   �
�(�(�(�(�(�(  �
�(�(�(�(�(�
  �
�(�(�(�
� �   �
�(�(�(�"�
�(  �
�(�(�(�
�(�(  �
�(� �
 (�(�
  �* `����  �(�(�(�(�(�(�
  *("(&(�(���
  * " & *"�*�*�(  * �(��
��(*   �(�(�(�*�
��  �* *�$�	�� �*  xd آ�� 8�x n� A�X )� �� �� )� �� � �ˢ
 K����آ�� � �� )�� D̥ �ɢd D̩ �� 8ʩ��% � aΥ D� aΩ �% ��dd&d$dd�  �d�$8�<��$��#8�؅# �˥#�%�&�ɀ� �ȐL�ƭ   � P� k� ��L+�L�� ��
 D̩  �� D̢�� <��P D�L%ǥ#JJJJ������JJJJ��
8�e�����  ) ��J�����  H)��)h)��# ��� � <� K̭  )����  )��� � #�`���L������ ����  � �Ǧ� � ��  �̢2 D��� �ˢ D�L�� �˩�� <���8�����ذ9� D̢�� l��������  �� D̩  �� D� ��2 D�L�ũ  ��  D�L�Ţ � ����e���Z ����ʈ��� D�z�Ș8����	��`� 0 ��i����� � ��`�ZH ��d

&
&
&��i��� 
� y7΅�L�i �hH



�� �}Vȅ�}Wȅ�`��@��R�ȱ�R�������hz�`�������hz�`  0 ` � � �  P@���  ` �  �������0 � P�p����@�  � �@  �������� ���@�`������ �  ���� �p�� `���@���@�� @�@��Q��  �� {˩ (����\��X ��� � <��  ��< D̩ � ����#i ؐ���# ˩  �d$d� ��+��  �ɥ�  �� {˩ (������  ���`8`�( D̥#�C��� <��#� �8��#إ�  �� �� {˩  �� D̀ܢd D���i؅����L�Ţ�� <��� <� )��� )��d D̢�� <��  ��� D� )�L��H �ˢ� l�h� �˩   �`�e��e��i ��`�'H�H�H�H� t � � ��������#��h�h�h�h�'`� � � ���`H)
������������#� Z���)����~ɀ�L�ʱHȱHȱ�hzH�)�� ��@�!�`�:�)��h�
 ����g�� ����]ʀ��)��h�
 ����JȀ� ����@����)��h� ����-�Ȁ� ����"�Ȁ�hh �`hhHJJJJJq�� &�����LY�hi�LY�H� ���� ������ {� �� ��h ��`��ZH !����� !����H�8� I�i�z��H�8� I�i���� i̲	�ɀпh��H��h ��z�`��� �˥ �˥ ��`��� ��`���# ��`��� ��`HJJJJi0 ��h�H)i0 ���h`HJJJJi0 L�h�H)i0 L��h`          #    � � �@�� �� ��������� � dd`��d�	� ����� ʎʎʎ`ڢ D��` K����`H�Z��� ������z�h`Hڢ �������h`��'��#Hd
�

�	

&
e	�	��
�e	�	�
i�
h`` ḭ�H�	)��	h	�	$%0�H�Zd

&
&
&��i���
y7΅	�L΅
� ��	�Ȳ�	��0��	�Ȳ�	��`��	�Ȳ�	�����	�Ȳ�	�����	�Ȳ�	����	�Ȳ�	��
� ��	�Ȳ�	��P��	�Ȳ�	z�h`H�Zd

&
&
&��i���
y7΅	�L΅
�� ��	�0�	����	�1�	��	i`�	��
���z�h`` ḭ�H�	)��	h	�	$%0�H�Z



H�
y7΅	�L΅
�� � ��	Ƚ��	�0���	Ƚ��	�`���	Ƚ��	�����	Ƚ��	�����	Ƚ	��	��
��	Ƚ��	�
� ���	Ƚ��	�P���	Ƚ��	z�h` � � � � � � � � � � @ACDFGIJLMOPRSUVXY[\^�Ȧ�Z ��H� � �h ��z����`� � BI�� B��� K�L~�ʩ�� � �8� i�
e��8� ie��?�e�z`Z�d��ϊ8����ʼ � �� �,�� �!��� ���z`��z`� ���z`��z`��z`H�� �-�� �!h�� ���z`��z`� ���z`��z`h��z`L~�b�y�����G���>Ѡѵ���X�c�n� LEVEL GET  READY !                    GAME OVER                     TRY TRY AGAIN.                      SECRET BONUS         SSSNAKE    COPYRIGHT 1992.    B.I.T.S      LICENSED BY   BON  TREASURE     CO. LTD                           WELL DONE      LEVEL COMPLETED                     BUT YOU HAVE NO     TIME  BONUS                                             WELL DONE      LEVEL COMPLETED                        TIME BONUS                        CONGRATULATIONS    SUPER SNAKER.    YOU HAVE BEATEN      THE GAME.       KEEP SNAKING!           PAUSE                              OUT OF TIME!                      PRESS  START  TO PLAY.PRESS SELECT FOR SWITCHSOUND ON.OFF    X 1    X 2    KILLS HIGH SCORE SOUND   ON SOUND  OFF    WELL DONE!    NEW HIGH SCORE                                                                                         ���                                    �P�                       ��        �T��  �?                   |@       �T��� ��                  �:       |P����: ��                 �Q�:       �����: G��                 p���      �Q�����: ���  �?          ?  0���      ��������� �G�        ��  ��      G���������  p��        p�  L9��     �Q���?   ��   ��:        0�  L:�� ?   p���>    ��  ����    �   0�  L����   ���     �:  �>��   G  0�  Lp���   G��      �� C���  �Q9  0�  L09 �  S��       �� C�  �  ���  0�  L: � ���:       ��: S��   C� 0�  \L: � p��       ��� �:@�   � 0�  \��� 0��        \��:�	\:   �: 0�  l���� ��         ��:`*0:    �� 0�  �j�p�  L�:          ��:�*09    L�0�  �j� �  L�:          �:L:�.p�    0�0�  ��:�G:  G�       ?  \:L:����    ��0�  ����  S�      ��  0::����  � �:0�  ���V�  ��   �? ��  0:0:@��� �� �::   ����   ��  ���� :0:P���A�L�L:   ���:   �� � T� �>�G0:@����0��  �   �� |@������0:P��G��:���    ��    ����������0ꀹ�Ñ��: ����         ��������:p��� 0�@���p�o� ��jA�   P  �������������>00逻��0� �� L��j ��? @ ���������� ��0p��?p�: ��0���� � ����������   l��	9L:P��0������4@TQ ���������    ��L:LT��������:PED  ����� ���    ��)������  ���:`U  ����  ��     �@���f�: �    �XU�  ����   �� ��? <�� �YL: �:     Uef   ��   \�: P� �� �fL� L:`f   ����         p�:�A�� ��? ��	L�0�Yff `�f�         0�:p���������L���f�������         0�:0��_�F���  �����������V         0�:���Q�~�: ���: ��Z ���          �:L:  ��A�{�� |�Z� �@�������         L�:L:  `�U�~9�����L: �  ��         L�:\�  ����6����p��    ��   �     G�:p�@��f�~������� 0�          9     S���� �������� ? ��        ���    ��������������?  ���������� p��   p�� ��: ����.   � ���� 0���   �� ��@Df�~��   ��^ ����^ p������A��  _� U��{� @�o�	�l�_�o� ����j ���   p�ef���{�������������� �����VU��: ����������n��������  �������� pP����~^����O�  �^�O��  \������� 0i����������o��_`毹��o�  𩪪����  p��������n�����������������   ������  ���>��F������o�������   𫪪��    ��l�Q�~����o���^��O��    ����       ��A�{������_�o毹o��_�o               �t�U�~鞿�������������������     U     �������{n�o�������G��   dj   �}��f�~꾷^���O����^��C�G�C�G��   ���������������o�_�o毹o������  @TU�9u�������������������������������     T�LM�������o�o�����������     �s�Gf�~�����o���^�O���S�G�S����3W��{n�������_�o毹��o�_������     03Mgf�_��������������������������DDDDDD4Mu�����~n�o�o�������G��G�������������_�o�O����^�S�C�S�C�GD����O����������������_�_�o毹�����������ӧ�������������������������������UU5y9�s���F������o�o�o������G��G��GD���;��{�Q�~����_���o���^�O���G��WU���O����A�{����������_�o毹��_�k��k��WU������g�U�~���������������������������UUuy>O睛�����yn�o�o�o�������������CM����f���~^�o�_����_��N�S�G�S�Gꫪ�~NM}��������������o_������������j����������������������������������������~>��o Q���n���o���SS�_�����G��G�Z����yD�E�~����_����TO=�z��O�_�G��G���U���T_Q��{����������tC}z~�����k���[��=uߕ]def�~����_�T���SӞ�������������Uս�tze���������SS}}M�Է����UUUUUUUe�u�T��Umf���~�����N}S��S�t���_�eVUUUYU�eu���^U��������}��:�P�^SMwz�ＹVe����UVU���We�������������ԥ�~O}������UY��eUV]�ӝWfm��F���=�ާ�T_����ӟ?�T3��UUe�WeU}�Խ_Ud�Q�~�S����_���:���4��OU_ED��~Ue}NS��U��A�{?SM��>��^z?�44�L3Ms�e��UV}N�y�_]e�U��4MM��C���^�W?5�LM��uE@���WU}O�y�������4M�S�~S����z���M�O��] U��_U�4S�NS���_��OMSMSM�����NMOS3�T3]E@D����Z���4SSs���T9S}SS�����O�P�O��OWQe������MS��y�O�t�S�S��y�G���sN�4M[EDU��z�L=}�ԟ�P=��~SM�G^z饗�t�>MO=gUUUf��������95���3���P��������z���SMכYU����NS�9M�T?������������?���S�Ukffff����^����O��4u^��:��ꪮꪪ��O��M߭�����Z�w^�w�M3՟��y�������������NSu�jf������V���z��S=u���^�UUeUU������w�SS����������U�����������A�WYUUUU�������S}�ջ������ZUU�����  ��_UUYUUeUe������}ӹU�������YUU����    �_UYUeYUeUUU�������U������ZUUYU���  @UU�UUUUU�UUeUU�������eU����jUU�UUU��  UUUUWUUeUYZVU�U�����7�UU���ZUUUUUUUUu  PU�WU]UUUUVUf�YeU���7M�UVVUUUUYZUUUfU @U��}U�UUVfVYUUUUU��7MM�UUeUUUUeUUUVU� UU}��UUWVfUUVieUUUU�NM��UUUYUUYUe�YUU @U��G_U]UUU�UViUYUV��SOSUUVUeYUUUUeU�  UU}��tUuUUUUVYU�YUU�~�LMUfUUU��UUUU� TUU�W���W�UUUUUU�UU�U��:�OeVeUUUUUUjUu @UUUUUUU�_UWUeUU�UVeUU��:M�UUUUeeYVUUU U�UUUUUUUU}UUUVeiUU�U���SMUUU�UeUUU�UPU�UUUUUUUY�WUUUUUUUYU��{�SUY�UUUUUUY�UU_@UUUUUUUe��UUeZ�UUUUٽ�:MUUUUUVVeiU�@UUUUUUUUUUUUUU�UUUUUUUYu�uN�UY��U��eYUuPUUUUUUUUUUUUYiU�WUUUUUU���MMUU�UUUUUUU5TUUUU�_UUUUUUu�vt�UUe������SU�UUUeUUeU5TUUU�zUUUUU�Օ�A�����S=O�SSUUUVU�UVUU��_U���_UUUUUU[y����N55MMMMS}UUeUUU�YUYm�����Z�_UUUUYm�]��S�O�SMMM�UUU�U�UUeeu�oi������UUUU���_��NM�4u��S�T�UUeUYUUU���������UUU�[�G�N55՜z>MSSQ�U�UVUUVU5y��G����UUUUU�U�S�O�wz:�S�DT�_UYUVUUZ54��C����_UVU�Y�UMM5uz�:5M�U�UUUY�UUu�t�OG����{e�e}���W�O՟�w�O5}@DT�WUVe�UU��_�������UU�V�_�_:5�yz��9�w Qe~UUeUUe��U�������YVV�Vyu�:5u���y�� @T��U�UUVe��UU������UYYWWzz�>�_z�w�9� Qe�WUUUeUV�UU�?L����ef֕�����Suz��WN^� @D��^UUeUUU�U�?\�o���Y��׫��T����Wޫ Qe�{UUUUYUMW�����Uye�f��U�_��G9䑗�� DD����VUUUUWTQ�^�����C���Q����� Qe����Z�UUu���wE��Wf���~�P�G�U^y����@DT���Z�j�]Ֆ�ߕ�ꕙj�C��Wz����ꪫQe������ZUU_������ze��:�Pz�W���������DDT�����UU�o����_����^�����ꪪꪫ�QUe�������ZUu��?�������Kz�������������DUU�����jU5�����������ꪪ����������UUUf���몪��U��O��_�������������������ZUU�������UO��O�����������������ꪪ��UUef����������L~�M���꿪��������ꮪꪪZU���������ꪪ�O���_��꿪���������������VUff����������U��UU������꺪�����ꪪꫪVY������������kU}U������������������ꪪjUVU�������ꪪ[U����WUU�������������VUUU�����������VUUUUUUU�UU�������������VeUYV������ꮪ��UVUUUUUUUZUUUU�U��������UY�UU����������Z�UVUUUUUUUeUUZUUUU���UYUeUVU�����������U�UUUUUUUUUUUUUUUUUVU�ee�VUeU���������Ve�U����������������UU��UUV�UZU�������jUVUUOO���O��7��T7�=�e�UU�UUeU�U�������jUY�UU�t>9��9�w�����M�UUe�UUf�UVe�������UUUU�U�}������w������UUUUUeYUUVU������Ue�YZUU�y������w����9��UUe�UVYfVUU����zWUUUeUUi�����~�w���y��UU�UUUUUU�U��ZiYiYVUU�U���������������UUZUeVUUU�YUUUUU�UUUUVVUUUUUUUUUUUUUUUUUUUUUUeU�UUU  �˜ d� �����҅� ��^��  ��<� �������(����� �  )����i�) \̥i/����2�d�@���âd�2�  )����H K̈��  �� �������(����� �  )�����D \̥i/�����̀C�ic��ʠ �������(����� �i/������d�@���ѭ   K�)���d������  )�����ɀ�`�'I��' � )� �ˢ��  �̠ �����  �̢ �̈���	 <���� �˥ �˥ �ˢ��
$'� l�d������  )�����ɀ�` )�L�� D̥'I��'� ����8e �!�� �!�� ������)`�V���IӅ�{���� d��dd'��`���  � ���#  ���& `�h��������������������������������������������������SUQc3Cc"c2!!37egVfWWwV�X���{�������TL˨�z�������ٙ����X���wfgSn��d���w�������κ��߻����d~ٶh�{�Ȧ�޼�˽�����ׇ��T�ǆ\�̺��������Ȭ��ʨ���C��u~���ɍ�����������ʻ��uK��e������������ݻ��ˬܼ�T6��Cm��خ��̻��ݷy���d%�ޖV��4Vgu7�Y������w���UuR��S%h��!'t!�R[��c$���c7�bL݇fh��1"�;��s#���C'��D���SFwa��vi��ECc�!J��R&��B9�لW���!!�rj��B$����e8��tz��v4�ۇwy��c3��!8��!jt�cDl�3{��R��V�̧B��R���BL��<��骼�˩�R��U���b~�b���C+���i������#���y���b��!]��s$����쪜�QN��f���t�� +��~���X���z�an��U���P��
����!�욝�߸��!o����� ��%���m�a-�쨧��C����r=�{��!8�1M��$x��1��[�� ���x���Wg1=�����2 ��!��L�1��tu��t
��8��1h1����rEx!=�v�� 
��J����	޶Vv���1��@z����)��14����67�������q80����c&v M�#d�� 
Α [��&�a��Vg��v!����a #ͳ ;ͦ!5� l�qEw��K߁ ���7� M�sF���f ��H��AU�� *��1Fv m�A5gʴ k�1���H�@�wu��e 	޴j��!t�[��W�m�qVv�� [�Q��G�Q	��He���!��)��PG��I��@7�@��f��Aα \���� ��eH��A ��Q���am�!��b����Bwkݣ ��
��Q|�0-��U��� �����1�1��{̨sI�0=�H���1 L� ��6�� ���r6��! l�q���'�0��t����ib��x��$̔ JͶ �� ��dq9��" ��a���9�q	��gG�ܖA ��@���:��S���Ri�l��4Fݶ J�a k������1��0�� 8��1��κ�����x1��Y��1&��	ޘW��܅�A��I��1xޡ8��a(�P	Φ%#��A ����Q:�q [ܢ�� )�a (�����̩�k�م�j��!'ʹ��톇q��G��ai@��E�ʄ�� ��SC[ݱ �Q )ݵ��	��A��R ����a}�A.�ʨg��wb��`���|�Q^������yu�q{��I�p>똹���yf^�j��H̒x��VS�J��!7̵�˚g�ݧUA߷��P��1Nݨ�W��e1��A���Zܢ��Uk�B�u��1��A-�ڕW��dA.�qK��H��^G��T ��1��Z����ez��u1��A$��$��������c�����p���y���eA��(��`��1o�ʧ����f�S)��17��!^�ʨh��vB�Q;��G��1��E��0 
�s)��1&��q����Q�s:��A&�����T}��Q�*��Q%�����e���s����'������w|��t��!���k��+��f6��~�1���h��a��Q\��A���Q%���	��DE����1=��!y�� ^��TI�����!������@���V���A�S=��`h���N��w{���1��@���������v���r��ޱ8~��1��tE���!�s+��QI�����EG�� �]��!y����DY���^��"y�޴��"F����A,��1Y���
��#%���<��1Y�����3F���#�����(���!��a$~�� 1��������@~�#l��1$f� }��0x�����G���$1~�������@��${��@#S�]��!g��o�A%{��U�<��Pg����5}�$R>�������R!��y��axA.�#������t1��!F�� $@n�!������u!��1G���Ut����D��̨0��BW|��!6c-�"���3y��A.�r���25�p߳@;��i���Sn�s7���B6�E�TA;��{���vS��5��ޤF���G!���v����c��dh���Dg�A��b���9���v!��Fy��sT��#���h��s����Vj���z��̪��遼>��f���u���a��bF��Em��!N��wy��vx�u�FS������f!���7���WX��1��tH��#F!^�0&z�"��T4{��vz�﷚��b��SM���z���e3_�!4Z������%���uH�!��C|���V��a>�$���i���wb��bW|�Ft�$:윒z��Ȇf5�݄Y�ʆ3��a�ʂ+���Y���S/�i��!#{s�y3Gܜ����ɖXC��W���ʙ����b���7���BXqn�TX��tUB�U(작W�ܘ�Y���SF���v��a�Y@^��j��6R�2g��aFb�7ی�w���uyS��2X��u���1�XP<��9��CgR.�UI�ˆTe��Q���Fi��wVwc��3j�̵V���A,��I��Dgv϶vuY�R#3.�"L�#f��eT��P��Ey��R5�ʄ���z�ݥVi���vf��QV���~�G���g���vA��s6��V���UVA=�d5���2W�v1� '�܄E���h�� ��uh��4�ژB ��a'�ۓH��n�0Iδv��R�dY��Bh�ܧ4b�S~�Ry��dDd!��BX��bg�� ��1&{˒z�T"�!;��SH��Cz�6�Xh���d�xxb!�D|��Sh�ܗUxx4��V��ܕW�˨d ��R,��Vz��eFT~�BHg��x��do�c��E{ܹfW�t�HX����gxxuA~�@9�ʄ%x��UFd�C$���Ri��vfv"ބ1]�ti��uUyd>�t8f��&U��T2��19̺tH�˗gy��U2��dx��egwS��bYh��%g��e31o�1�ʆF�˘fx�Q>�D'޻�V�ʈgw�d�fs�y��Vi��uU1.�3�˨E���ww��!��s|۬�W���wwvS	�G'���dg���ffs�E%�ʪu�������B>�u;���f���wg�t ��cxw��Eg���WgR�D)���ew��wh��R�vW�z��Ux��UfeA=�TX���Uf��vVwvA<�Vhw��Ufx�wUgvR&�Wfvx�tUwwveffS&�Vfwx�uegw                $ L:�H�Zح' J� ���$ �	J��%  ��z�h@���# `�`$ L�H�Z����$���� H��
z�h@�	L���	` _� <� _� <�L_����B���  ��� � �F� � �G� �ߍ& ��" ��t ���d@��A�� � �@����A��� ����� X�ߍ& ���D ��  �� �S��U��T� �L���M�M�K�L�J t��M�r� ��M��d�N���O�M�M�K�L�J� �S��T t��O�O�O�K�N�J��T��S t��O�D� �L�� � ��M�K��T�L�J� �S ���Li�L�J t��N�J��S ���N8��N�J t��N�T� �L���U��T��S�L�J�J�K t� �� �� ���2 ��� ��xd `H�Z�S
�� ��@� ��A�T�P�U�Q�K�R�K����V����W�JJJ��@%D�V�@i�@�Ai �A�Q�Q� �Ȁ��P�P� �
�R�U�Q�L��z�h`H� �D t����Dh`H�Zd@�@�A� � � �@����A���z�h`H�Z�/���� ���� ��z�h`H�Z�X�B�B�P0�B�B�C� ��C .�z�(h@H�' )��B�E�# �$ �% h@�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L �LD�L\�L8�������