���� ��d� �������Ʌ������ǀ�Ȁ ��������兦���� L����	���������� L������������� L� ��8���P����JJJJJJ)�
����H���H����������zh� � ��  ) ��  )��  )�С`����������d�  ����LK�*    ����� �? �? ��� ���� ���    ������ 0� 0��            �UUU�  � 0�0      �   0    �Z   � p� pUPUUUWUUUCUUU    �UUU: p� p�\��W5W���sU�_�   �kQ��� p� p�\5 \5W  p� p�   �Z���� p� p�\5 \5W  p� p�   �����  p� p�\5 \5W��?p� p�   �E�    �� ��: \5���:�� p�   �Q�     �� �����:���:�����   l�>     �� �ꬪ��:���:�����   l�     �� �ꬪ�����?����:   l�     �� �ꬪ���  ����   l�     �������? �  ����   l�     ������?   ��������?   l�     ������?   ������ ��   l�     ����?�?   ������ ��  l���?    ����?   ������ ��  l����   ��� �?   ������ ��  lQ���                        �UU�>                        �V  �:  �? � ��� � ����   �jUUA�  0� 0�   0   0    ����  0� 00   �   �    ����  p��UPUUUWUWUUUU      ��  p�pU\��W5WUW�UUUU     ��  p�\� \5 \5WUW�U�U      �  p�W5 \5 \5WU5W�U��      �  pUU \5 \5WU�W�U         �  ��� �: �:����Ϊ        ��  ��� �: �:����Ϊ��     ��  ��� �: �:����Ϊ��     ��  ���: �: �:����Ϊ��     �F�  ��� �: �:�Ϊ�Ϊ�� �����Q:  �ꬪ����:���Ϊ��� ����j�>  ��������?�������� lUUUU�  ����?����?��������     �  �� ������������� �ZUUUU�   �� ������������? ������>   �� �� ��? � ���� ������                       ������                        68��E�                                      � ��     ��
 ��?     ��+ ���     ��*���� ��  ��*���� ��+�����
 ��*�����
 �

�����
 �o������ �o������ �o��ZUU
�� �o��VUW��� �o��U�_��� �o���_���� �o��UWU���  �o��VUU���  �o��jU���?  �o�������?  �o�������  �o�������   o�������   o�������    o������?    o������    o������    o�����:    �o�����
    �o�����    �o�����    �o�����     �o����     �o����*     �o����*     �o諸�
     �o�ꮪ     �o����/     �o����?     �o�����     �o����    �o�����   ��o?���   ��o? ��   ��b� ��   ��b� ��*   ��b� ���      � ���     � ���     � ���      *           �           �                                                        ��          ��  ��     ��
 ���    ��
 �    ��
 ���    ��
 ���>    ��
 �Zj=   �����ZY�   ��� ���ۻ   ����ꪪ�   ��ۿ�����   ���������   ���������  ���������+  ����������   ���������  ����ꪮ��  ��������/  ����������  ����������  �ۿ������� �ۿ�������  ۯ������  ۯ������  ۯ������  ۯ������?  ۯ���*��?  ۯ����
��> �ۯ����
 �* �ۿ���� �* ������� � ������  �� �ۿ꿫:  �� �ۿ���  �� �ۿ���  �* �ۿ���/  �
 ������     ������   ��������   ���ÿ���   �������   ���� ��   ���� ��     �  ��     <  ���      ?  ���     ?  ��
     ?  ���
     .  ���     *           �           �        (c)1992Thin Chen Enter.  Push START Button Stage: � �I�@�J��I����J�J�`����
�[��
��
��
d���
����
����
 �� A���
�����
���⥤i<Ť��`

�� ��� � �����`� �/ ���
���
`���
��
�@�]�<��8��
 ���Ii0�K�Ji �L��
�����K�I���K�Ii0�K�L�Ji �L����
���  ��
�a�1�]�-�D ������IȑI�� ��� �I�Ii0�I�Ji �J��ߩ��
� ��
�_��a�Ș j���
�a�����
`��
`��
���
`��
�M�]�I��8��
 ���Ii�I�Ji �J�Ii0�K�Ji �L��
�����K�I���K�Ii0�K�L�Ji �L����
��� ��
�a�1�]�-�D ����ȱI��I��'��� �I�Ii0�I�Ji �J��ߩ��
��
�a�����
`��
`



}"��K�#�i �L�J��� ���&�eI�I�Ji �J��K�I��`(�(� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 ���  ��� � � � � � �� � �( ����ÅG���H ~��@�LdK�� �K����L�L�`���
��
���� S���)���
���
��
)�S��
��L�Ə��
����
�͏� =���
�ԏ��
� ��
�ۏ�i =���
L�@@@@@@8  0@P`8@@@@@@p�����Т ��
�	��
8���
�����p���
�	��
i��
����������
��
i��
��
ɀ�Ly�d���ɴ��  ����  ����`

������
�����
�����
�����
��
��
��
i��
��
��
��
��
i��
��
� ��
��
��
��
`	
+,)*78'(56%&34#$12!"/0 -.                   P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*������������������������������)���
�`��
��
����
��0'� �����
����
����
����
Z ܔz�����۠ ��
����
����
����
����
�Z Ĕz�����ة ��`��
��
��
��
��
��
��
��
���
��
 ����
JJeI�I�Ji �J��
�



eG�K�Hi �L�JJJJeL�L��
)��
��
��K��
��K��
�
.�
.�

.�
.�
���QI�Iȭ�
QI�Iȭ�
QI�I�Ii0�I�Ji �J�Ki�K�Li �L��
�L�`e�Ť��`� ��
���`H)�����IhJJJJ�J
eJi@}���J` 0`��� P���@p��      
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ������������������u����� t����������M�������H��^&�G% �����������w�^&9G
u� �+������t;���� t4����j�5�wRP��M�������������j�5�wRP�N��������������d
���~���P���+���+�����Pj����P����P����j j �HO��>.  u�9���u
���� t�� V��WPj�W�����>  tW�I��t���� tǆ�� �^ǆ�� �V���� t�Eu���� tǆ�� �:ǆ�� �2�Et���� tǆ��	 �ǆ��
 ����� tǆ�� �ǆ�� ���� t���� t	�������ǆ��  ����������P���+���+�����P�6~�6��6��~����P����h� j ��K����� tZ���� t$��������������M��������������N��/j�5�wRP�z������t��������QP���w������H��N�^��&�u ��������P��w�y��FFt�~
u�h������v�v�~
u� �+�P���F��V����F�@u�<�����P�v�v�o�����P���F
- t	Hu�� ���Eu&����h	j j j ���w;F�uVhF	j j j ���w�����v�vj �s�F��V�=��t���VW�v�����P��F��V�V��W����Pj�W� tC����P�v�v�o��v�����P����j�W% P��F�+ҋ��Gt	VRRR�'�w����h	j j j ���w�F�;F�}�=�����h@P���~� u�(��Et<�F��F�����h
�N��v��F�P���w�F������E����8Gw�u�O��g�����hj j j ���w��������h	j j j ���w�F�VhG	�v�j j ���w����h�v�j j ���w�F�9F�Y����hj j j ���w)�������F�;F�~����h�F�HPj j ���wVhj j�����h�F�+���Pj j ���wW�_�.��FHtHu�� HHu�� Hu���V��W����VhH	����h	j j j ���w����P����j Q���w����P������h����P���-��P����P������������RP���w����j��&�����tA�F
 ���� ~����hj j j ���w+���Ht�F
�����h �v
����P���w���������P�������~�2��6hje��V��WPj
�v�W�v��V��WP��V��WPj
j �W�v��V��WPj
�v�W���Vj �W�t�a�����h
�v
�F�P���w����P�~��EP�o�� t�Eu����P����F�F��E*��.�������;F~� ��������w����P�6x��M�������������PP���P��K��d
����������� t����������M�����������w�d
��������~;F�|�����h�v
j j ���wVhj j�������wj�FOw�Āu�Y������FP�twV�FP��w����P�F��+�P�F��+�P�Q�R�=wV�Ԩw����Pj j j ���w�t����P���w����u��(w����u5��󚗁w;�tǆ���߁��� u�����P����������w�u��V��WPhh����P���w����P������� -�6
Vh������v
Q�6`j h-���P����  �.  ����j j j �'�w�-��N�^��&�G������P�v
�4�N�^��&�G����;�u�k������6�j �������������Pj����J�~
 tj�FOw�}qǆ�� ����9. tP�. ����h����h	j j j ���w����P����P���w�t ��������Pj �'�w�����]�w�~
 u���  �P���w���j�FOw�|j�FOw�}	ǆ��  �v��^&�w&�w&�w
���^&�7&�w&�w
������;���t� �+������9��N�^��&�G-�r- v�S�>.  t� �� $��F�����&9Gu&��u�)�  ��<��^&�G�F�&�O����VhH	P����P�������w����P������P�����_��u�r���UUUUZ�5QA*RԒ�A J���Y*�[����������R�+��jm�����[��P�(�mZ��U�յj��$�*���￾�k%&R�R"PH"�ZU[[)JBB@   �R     A@   %*�W�DQAH�!Q  ���     � �R�Uu�֭����B�
�J�H����UR�� �$�ER��EQQ$H  "�������)
   � QJI! @      �P         @   
 
�E�DQAH�!Q  ���   
� �R�UU�֭��z�B�
�*"H����UR�� � �ER��DQQ$H @"�������)
  � QJI!@B   @ �P        @  
 
�E��                                                                                                                              5JUUUUUVʪ^�T$P @� *$EU�U����������U"
��ݫ�������T���U���Z�]j��*�T�m�uuv�����ID�R�� A%T�JT��  D
E @@ �  
  �   
B�X%@T�J�D       "$E5U��ޮ���]��"��T�*������$��)��H��M*����UUUT�����@@�@��  T�JT �                   @��P-@T�J�D  � �"$EU��ޮ���]֖"��T�*����$%� �)�H��L"���-UUUT�����@@�@��  T�JT�    @    �     @ P�P�                                                                                                                              D�UUUT��5UQ��J�D!*�@ɺ�Uww����������U��kUw]�ߺ�l�PJ5Zvj�ֻz�WV�RI"�i������j�IU*D�*!@�UV���H�   @ RQH    � �  
@�,�K� @AA@��%P�B     $ �� eU�5���[ꭺ�A
��JUUUZ��D�@JR$���"�E P	 � ���UUIJ
 @*@   Q��@       P        �   @ D� %BAAH��%P�B�@   $���e�5ݵ�Sj���A
��JUUEJ��D�BRJR!���"�E P	 � �ҕTTIJ
B*@$   %Q��@      P@     �  @ J"��                                                                                                                              *�����UWM*J��DT  @   �"���[���������� *J�����������J�J��֭��׻j�U�"�(�k�u��]V�$���)@� �%%UV�) �    !J�        
D  @UT T�U�(�(�(!H
B��        "*J�[[�koz��{j *�����U�����H  B���(�*U*(�U �(R�Uj�U� � !    � DT�(      JD           P D�Eh(�(�)!H
B��      "*B�K[�kmj��+h *����������H B��� �*U*(�U�(EJ�Q*�U� � % "$ � DT�(     JD         P D�M(�                                                                                                                              *��UUUU��I�UB) �  B�"%L����������{����U�խU[���{��H�T�ս�Uv�UUV�)T�I)7_���Z�IEJ��R
	 IUkiIRiJ B  (�!   �   � �J�T�"� T@�@�B      !  D��*��Z���mz�֡�UT�
�UUU+"%�AUKUT�QD� D -UV���R�HDJ��R    IS)%	B B       �              �  J�P�"��T@�@�B   �!! D��*��X���mZ�֡�UT�
�TUU+"%�AUIUT�QD� D �%UV��"R�HDJ��R   IQ)!	B B     �       @      �  J�R��                                                                                                                              $�iUU*�JV�$�R�H�JR�jUn���������	����ծ����V�)!U�.�Zۻ���UQD�$�J]�����֩"RIJD� !�UJ����    $�� P     �   �(�*��$�)UQ�B��       
**UJ������Km�	ƨ����Q*����L�  D��R���+T�$@JʩUT�D  H �   B��(�       �$         �     ��$�)UQ�B��@     �
**QJͷ��6�Km4	ƨ��(�Q*����D�  D��R��)�$AHʩUT�D   �  B��(�     @�$        �    
���                                                                                                                              )JV�U�*�5��%�)     @AJI(�$��������o%�E��-U�����v�T�JU*���Um�l��UR�T��߷wwZ�JD���"��D E%T��T���   �H�       @  PD����BB � ��P        @ � �����v�m��[m�
��% ���*�*�D��"T�4j�D"�PD*�UUU�J@��"�     D�"�       H�                @��*�BB � ��T	 H     @@� �����v�m��[m�
�� �*�*�"�D� �"T�h�D"�PD*�UU�JD�R��� @   D�"�	 �     H�              � @��*��                                                                                                                              *SIj�UUJ%*� �    $!RR��T������������*��ꪯn����ګJ��j��oV�֫T��-&�T���]��Y)I)J��(JU�K��� A    5*�@@� � 
� "A
"ih"J�UJ! �         (DR�mWz���w�v��"	U(�j�Z��T�i ��"VʑJJ�)P�%$ *�UT�� 	  
cJ��       "�@      �   @
IH"(J�UJ! �     (DP�-Uj���U�V��"	(�*�J���T�) ��"J�JB�)@ �%$	 U*�T�� 	!  
#J��    "�@@   @B�   B@
IX�                                                                                                                              %-U*�JR�UJD�(D"@ "I�%�Z�o������߼�%@J��Uu����kv�T%R�uO���T�RJ���P�+w���kj�BJ)*B� �"�Jt,)D   ED�       B  �T��*�$E  H " HD         H �	R�m��W��zݴ 
��� ��V�+JԔDPIQ*�T�R�B
��  )
�R��Y �  B)"   �P!       DD            � D �"�	$E  H " HD @      H �	R�m��V��jՐ 
��� $�V�!JT�DPIQ
�T�P�B
��  )
QR�#I � �B)"
 �P%      DD            � D �"��                                                                                                                              *��Ҫ��,���T� @  ITR�d(T�*�{���������"H�[j�׮������ �UV�Z����j��RU
�R
V�}�^��,����ED� ������(! @  �	)*�    �*�  *(���d ������       B$ T$"%*�k����իm"@

��(�R����Y(� !TFT����J��P�P �U%T���"�@    ���@       		
       �     �$ ������    @  B� T$"%*�k.���թm"@

�
(�R���U(� !FP����J��PH�Q �U%T���"�@@   ���@ �    		
@      � @  	H�$�                                                                                                                              %+%*IUQ$�        �$�IE)J��߿�����������ڵRSZ������UU
*�����[]Z�J�IT�%QM��kmڪ�!�D�2�"RUjU*��$  @ �UD       "@��B�V�RSX!Q Q �            	(���������v���T�B
�����MT�(���eTITPB�  QL���)H� �D� � BI*
       
T@        @  B@ �QH!Q Q �            �	��������v���P�B
*����ET(���%TITPB� QL��I)H� �D� � JBA*
B     
T@        @ �B@ T�QH�                                                                                                                              JJZ�V�j��RT@@ $� %�)")Jim��������ڮ4���J��[���}��SU[{km��ꪫT���*H%+~ݽ�WJ��U)��D�  ����UUPX �  $!�)  �D  	J�  *� 
UUP R�T* D         �("@D�Un�o{mmګZ*�
�J("�Uj��ZR� E
SIJ��B��  @T�%J ��D	"@    �(�Q@P �      �)          *� EP 
R�T*
D@     � @��("@@%Uj�m{ilʋZ*�
�J"�Qj��JP� E
SIH��B�� T J@T�%J ��D)"@$   �(�Q@P �    ��)      !(   *� EP�                                                                                                                              *��J�&��J�A	 @I $R�IJT��]���������JB�/oV����־��Kj��UV�^�u��J���RD��Jն�V�ڪ(��%JH�"B�)UUJ��  � 
j�    $ D@UT�Z�
��
"��@�              B��UU�����U��
B�*�R��%Z���Jh��T�V)%$�H���  �J�d�U�J(�!    �	��      
*D           @ UT�J
��
"��@�          B��UU�V��U��
B�**R��%���Jh��T�V)$ �H$��  �J�$�T�J(��   �	��     **D          @ UT�J�                                                                                                                              )*MU"X�%P	     J�A$���io������t�����RQ���������*�j��ʮmkuUUUT�(U�mV�j��BTT�J!@  ���UHRT   �T�       A@  )@��UR� 
P"(          @$ �)J�_k}V��mԐ��R�P���Z��� �J����I"�UP� 5YR�H��B� @  �*�Q@P       �        A@  ( �R�$
$P�(��      $H$ �)J�[+UV��mT���R�P���J��� �B*���I"UP� %IR�H��B� A  �T*�Q@P    @ �       A@  ���R��                                                                                                                              "��HIC*�   �"I P����QW��������{�%�^�uL�m���nꪪ�B��u��i�Vʪ�R�EEJ������Z��IIRT*�"$U���UT��  �$�@     �� �J�Uh ��  A          � �%QMU���W�kkR���U�IU*�Z�*��@$)"��!RT@��B� D �E%T��J$ �@@BP   �D��      $E@             �DH �� A�  �     � �%QET���U�ikR���U�IU*�J�*��@ ) ��!R@��B� D�A%��J$ �H@JRB ���      $E@        �   T�LH�                                                                                                                              *T����PH�!  �  ��"��,UU	*���������rHV]�*�%W[����jR�Zʵ��U5,*���!*�okj��A!���@ IJ*���%PB@   	( @     *b!$@H!	*�* ��� @            �!$E �mn��V���pHBZ"  JիUSU"�JJiRJ���$ �$  *�J)*�! !�  @  	H"�"� @       	         
@ $@ @	"�*���H@           �!$E �-n��V���pHBH" �JԣQSQ"�JJ!RJ���$(�$B *�J)*�!%�  @ �	H"�"� I �   	         
@ $@@	"��                                                                                                                              $�J$B� � 	"  )A%%2J/k�߿���k���P�=[ꪨ��WޯkV֕%%V��5UUUJ�J��%R�J��֭j�H��T�T�HRR�UJ�J
    $	J��  � @ 	   J�
%N��P �H                 % H�*ݶ����j�D��*RȊ�U5T��RL� ���TPD@�@ �� T�ʥ(�H  (�D  @TAHJ       B�@            B�J*U �H         �    �% RH%*Ֆ����*�DA�(RȊ�T�*RD� ��%TPD@�@�� T�¥(�H (�D  @TAHJ      B�@       �  B�J*U0�                                                                                                                              )(��*� �  @@ !@��I*�RD�Un����������E$+�UT	[v����ު��UU�}n���j�UJ��H$�J��Z�U�R�)D�i ��UV����     !�       T  V�@��Q$T   ���          @ �	(  ʫm��mn�l��D$	�@	*j�UUL��PD�U*E��*B
�H J�%)E  	@�@   ��� �       �            � �A$D(� ��H��       @ �)( J�i�]m*�L��D$	�@	"j�UUL��PD�U*��* B
�H J�!)ER IB�@��  ��� �@    �       R   � �A$D�                                                                                                                              $�B @ �@RQ!	 R�HP����۾�����w�R�].���UV��ݿwuک"��{��j�R��R*4H�Iomu��UB))T! 
R��T��!D �  �EE+@      " � !J�V�           @      � �������{[�տ[� H*T�@RR�UUUQJ� �))Q(*J��@  @*�T�(   	   B"%R�!        E"@            ! J�R�$      @�      ��������{[�յR� H*�@RR�UUQJ��))Q((B��@ @*)T�( @ 	  B"%P�!       E"@           � J�R��                                                                                                                                �	@� "    �B��P�""�	 �'�������wݥ� �;�UR �m{wkݶ����UUZ[�R�����B�$�!#jګWT�RR�ʤU"�@�J*�UIJ�D    )R�  @ @   @J@	h)J��              � �    � *������T�e� �@ IKkUj�&  �TJ*�@�*A $ JJ)D�@�B Q    �D�H
       R�            
@( @($             ��  � "���Բ�T�%� �@ 	IkUj�&  � TJ
�@�*A�$ �JJ)D�@�B Q  D �DHJ      �R�           *@H� @($�                                                                                                                                 � ��R�(�I$H%TU$��%*m����������X���URZ�߿��m�T&-Uj��U�WUT�T!) T���T�R���I*�D( *�UUV�RH�      �H�         � BER�P              �	  T$"�!"J��u��kk����H���5T����h� "	UB�QA%UT�@  @d�Ġ   
 @   S
         �            � �P            �)  T$"�!"H��U�mkk����H���T���� � "	UB�PA%UT�@$@$�D�  
 H  Q

�       �          � �P�                                                                                                                                "   @�D   ��I(H�HI"BT���������t�/{V��}u�[�ڪ�H�*����j��E)R�JBD�"�UUU�� (��D��� UV�R��!  �MBU   @     " �T**X                �	  @�   ER�{�w[�\�EWT*��@ �UUUV�ʤ� �**�TH � @  @ �U��   "@�     RIP��       EBQ            "  @((H          �    �	  B� � ERZz�w[V\*ET**@ �QTR�ʠ� **�TH � @ @@
 �U��  "@� @ @R)P��$      EBQ        @   " PB)(H�                                                                                                                                 EQT�JT"�@�(��H��*��������h!޴�����V��_�J"�����6��T���J��K��U**J*A(�!PJUj�UU��     (�        	J 	�R�           "�@ ����VֵZ�Z�� ڐ�����B�Zժ��H� �"��R�� ��
H� 
�DL"	!@  
QH�E$       �             H �R�  @ �  @! "�@ �(���V��Z�Z��h ڐ�����B�ZU���H  �"��R�� ��
H��
�DD")!@ 
QH�E$ �    �            H �R��                                                                                                                               �� @  ����֊��%%)%*�	Jn��������J&���W�j��u��������e��T�+T�T��)!�U�UQ�EE	JT�*���VH      JJ�           � (RIM(        �   ��D

   J*U�^�Uj�
%`"�R� UT�U)T���(�ID��*@(@    �!Q �     ��R       B*            �  RI( @   �  � @��D

 �  J*�\�Uj�
$ "�R� UT%U(T���(�	T��*@(@    �!Q@��     ��R      "B*            � RI%(�                                                                                                                              �Hu�"Hu��Hu��-- u�Hu�W-1 u��Hu�Hu�Hu�(-a u�8Hu�EHu�N- ry- w�aHHu�- re- vrHtf-W u�HHu��Hu�	Hu� 	- u�	Hu�	-�u��	Hu��	Hu�
Hu�
Hu��	-` u�
Hu��
Hu��
ǆ��  �#Whjd�Q9>u�KW����P�(w���uǆ��  ����u�����	�����+�������W�����17�u�Wjh������������w��
j�FOw�}�6hjnj j ���w��
W�����
h�h�6`�� '�F��V��6`j j�h�h��6`�� '�F��V��6`j j�vh�h��6`�� '�F��V��6`j j
�VWj��&�F��tP�u�wh�hS�6`�� '�F��V��6`j j,�!�60h�hR�6`�� '�F��V��6`j j�� �60h�hR�6`�� '�F��V��6`j j�� �60h�hR�6`�� '�F��V��6`j j� �42tIWhh����P���w����P�W����P�2= u�uW���	j �I�����u�t	ǆ��  �����������������Ph�������u������_���� u�8	h�h��6`�� '�F��V�����~�6`j j&�6RP�;&�	�6`j j��h�h��6`�� '�F��V��6`j j��Wj��&���tWj��&�����u�Pjj j j ���w����h	j j j ���w��������h��pu� �+�Pj�j����w��qu����hj�����RP���w�jW��W;t^Wj �W�����tNP�x������������h
j �F�P���w�^��������&�G@t����hj j j ���w����������jjj j ���w����j j j �'�wWhj jW���j�FOw�}�6�  ���>� t	�f
 �h�
���>4  t	�6�  ��>  u+���6`j(hZh� ����6`j)h�h;���j h�hZhA�]�wHt�Aj j j �o�3h�h�6`�� '�F��V��6`j j����>Tu�&�V�L�M�60h�h  �6`�� '�F��V��6`j j�6RP�;&�����v��v��� '+��F��F�����}��>"  t>�6`h� hZh� ����6`h� h�h;����6h�hZj4�]�w= u�6�6L�6V�
���>&  t�P�6`j7hZh� ����6`j8h�h;����6h�hZj�]�w��6���
�>Tu`�&�V�6`jFhZh� ����6`jG����Ph����VA P����Ph��Z���
�6h�hZj4�]�w= u7��60h�h  �6`�� '�F��V��6`j j/�6RP�;&= }�o�&   h�h�	�6`�� '�F��V��6`j j�6RP��	���tX�6j ��w�6`jHhZh� ����6Vj ���t,�>&  u%�6`jKh�h;����6�h�hZj�]�w�>� u���6j��w�6������  �j����@t@�6j�p������tm= t(= u�����h�h;�\ ��6`jPhZh� �?�h�h��6`�� '�F��V��6`j j�<��6j�^���6j�g������u�
��(= t�= u��Wj��&�F��u�	PhF	j j j ��Wj��&�F��t,PhF	�Wj��&�F��tPhD	j��Wj��&�F��u�PhG	�Wj�W%  �F� �9Wj�W%  ��h�h��6`�� '�F��V��6`j j�b���5��F� Wj��&�F��tPh Vj �v��W�9>t�� Wj�v�W�6h j�-�h�h)�6`�� '�F��V��6`j j ���h�h�	�6`�� '�F��V��6`j j!����> ��أ �F�h� P���6����P�(w�6jj �����������wW�~�6j j j�'�w� �@\�B  ���Wj��&�����u�uWjWj�W4 ����P�W���� t)Whh����P���w����hD	j ����j P���w�����j j j �'�w����%  �F��,�>4 ��أ4 �F�h� ��> ��أ �F�h~ P���6���P�F� P�������PV�~���% P����Whj j j ���w-A PW�  ��6
h'���6
h&j�FOw�|� �+�P�r��6
h(�f�ǆ��  �����㋇&����ى��������|�ǆ��  ��6jgj j k�����������09���|��K�W��ǆ��  ���������}�����㍆����؋��;�&t�W��������W�~�� �F� h�
���6h$�v�hp�<W�t� �6j|h� h0��� �F����F� ��6`j|hZh� ����6hZj j j �  ��^h�hP�6`�� '�F��V��6`j j-�*������09���|��k����������;�w�d ;�v��6��+���Pj j ����~��F�F�t�v��v��� '� ^_MM��]M�         �����N����F�V�V��>  t+
�V��6
����PP�v�Rj���  �>  u��6�F�P��  �F�+
�F��v�F�Pj�k  �V�0   �vj���  ���>�~
t�~
V�u,�~
V�u�F�F��^���F�V�F��V��^��F�&�? t
��+��F��F��v
�v�v�v��v��4���FFt�v�vhf��  �u8����6
j��v�j�[  �F��tPj��  �u��v�PPj���  �ՋFFt�v�vhP���  �t�u����	��r@ �6
j��v�j��  �F��u�JPj���  �u��v�hPPP��   ���v�v
�v�v��u��~ t,�F�V�<�>�F
�:=�r=Ms�:��� �~
 u�� � �F��   jsj j �y	`�F�� �� �>� t	�f
 � �F
s �v
�v�v�y	���t� �~
st�2�@���>D r	�6D���  �v���  �s�:��@�B  �$�~
 u\�>B u�>@Yr�>B u�>@�w
�v����4�v�j�P�6�j j j ���  ��v�6
�v�v
�v�v���  �+��^_MM��]M�
 X�EU���؃~ |U�~u+�^&� u[&�puT�6�6�jj &�7��  � �=�~ u�^&� u*&�pu#�6�6�j ���v�v
�v�vh6���  �+�MM��]M� U���V�F�  �9Fu�vj��vj
�   �F��u+��Phj j j �T  �F�� �@�� �@��  �<�A��<�A    P    �         � ;`=H ;�=    ���  ����    n#    P   = �        �      ;�AT;�A   ��� ����    n0G     P   ��          ��     `=�A`=�A��H/h�:46�)l �$P�$ `          46�:2 2 � > �S�=�A��=�A��`:H/h�:46�)l �$P�$ ` � �        l �)� �Q      �=�A|�=�A�        �$l � �$ $         � �� �          �=�A@�=�A���:46�)l �$`:H/hP�$ ` �      �:�>H �:�@  � j8~� jt>�A�t>�A�#   �  P   g         �      �:4?H �:�@  Cj�~Cj�~�    �#   �  P   h         �      �:|?H �:�@  � ~8�� ~8��    �#   �  P   q $        �      �:�?H �:�@  C~��C~���    �#   �  P   i         �      �:@H �:�@  � �8�� �8��    �#   �  @   j <        �      �:T@H �:�@  C���C����    �#   �  P   k           �      �:�@D �:�@  �p � �p � �    �    P    T         � �:�A�:�A��H/hP�$ `46�)l �$                �@�A� �@�A��`:H/hP�$ `46�)l �$ �r[�v���x�~��z�
t��F�t���B���@�A� �@�A����W�Z͊��F��t� �RȋN���FǊ��RʋF��tA�R�_먊F�
�ty��� �ΰ����})�_^�f�]M� i( l(?pl?e( V(?pV?!  �<�A
 �;�A 




 
p � `   !p!0 q�F� ��~O~U�^�G�F&�G�F�� �v�F�  ��7
��ts��� ��F�V��F�'��&�O����&�q����(��F�A� 3��:�A3ҋL��\�+�s��+ы|�߱�|u��� T�V���D
+ǉF�2�N��~����v
�F���K����
tQ�^��|ۀ� �� �ۈ^Ɗd�D�~�v���ub�~�}t"�m��P������������n����X��p��9u+tF�~�u�����������$? ����?�� ���u+�ފ�X���ދ��E(= w�= t�= t���E*�^�����q�I�i�nċ�}(t�i �^ƀ���"���"�
���t�}(u�ފi.���Ոn���u�f��^�.��1��@t3�3Ұ��F�u5��䰀�vȄF�u�nĳ�� ���� ���� ����� �F������
�y� t����.����
t�.��1�Nŀ�F��� tV���2�
~�"�:��
�yE�~�Vȁ���ӉVʺ�."�  .2�0 $�� ��.��  �ΰ��F���f���F����I��t��Ę2�2�2�0fĈV�v݈NՊfĈf��F�U�F�+�'�ؚ� ��ڍ>������=����FĈ�2�6�l2�6�\�^��ŀ�w
����.��6�\��
t)�nƀ�
ݗ3�.��� �6�D��.��� �É6��2�������v�N~���Э��+�~�vK�N����^�"�2�ڋ�"݊�ʸ������˻ ����̀�uU~�P�F�� �X��2����u"�3�FN:��:��:��:�ډv�II��;����#ъNǊ�#�#ىF�^�= �#�����~�P�F�� �X��u#�3�FN�Ć�;��;��;��;��멺�����FՆ��F͆��F݆���F�3�Ú� �P�� ������3���X�� ��ú���ú����#���!GG������!GG���#�1GG���#�	GG��Ë�#���Ћ3�#«���Z͊�Ë�#���#Ћ3�«���Z͊���В�3�#�3ë��ø��=3�=����[+�s��69
 w69 v6� �����6�
 6� 3�� ����                        GetKeyString Esc Backspace Tab Enter Ctrl Shift Num / Right Shift Num * Alt Space Caps Lock F1 F2 F3 F4 F5 F6 F7 F8 F9 F10 Pause Scroll Lock Num 7 Num 8 Num 9 Num - Num 4 Num 5 Num 6 Num + Num 1 Num 2 Num 3 Num 0 Num Del F11 F12 F13 F14 F15 F16 F17 F18 F19 F20 F21 F22 F23 F24 Help Clear Break <00> Prnt Scrn Num Lock Num Enter Right Alt Home Up Page Up Left Right End Down Page Down Insert Delete Right Ctrl Acute Grave Circumflex Umlaut Tilde Cedilla �     % * 0 6 B H L R \ _ b e h k n q t w { � � � � � � � � � � � � � � � � � � � � � � � 	 &+5>HRWZbgmqv����������*6789:;<=>?@ABCDEFGHIJKLMNOPQRSWXT`abcdefg 	
 !"#$%&6%&'()*+,E58EGHIKMOPQRSFTV\789E:8;<=>?@ABCD5634E:9	�'`^"��~��FFGHIIIJKL��EU����VW�~s�  �� �F<Vt<5wHr��uA2� PS�  �2�
�t/� PS�  ��Āu< v�^&�&�G � � �����
 ��F��u�a���/ �	����� �W�Yu�+�O&���t����� W�Yu+�O&��>  r-P�  �6 P���@�Xt�B�~�^2�PWS�@�&2����.����~3ۋN��
�tC��2�O���_^�f�]M�
       X�EU���؃>.  t�6`� +�RP�����6`� $���MM��]M�U���V�v��WPj
�W�F�P�x�F��V��vh�vj j ���wk�	�v�&� �F��v����F�^��]� U���vh��Y��u� �vhl�Y��u7�x�? t�F�^�?.u��?.u�F�	&�? t�F�^&�?.u�&�?.u�F�^&�? t)�^�? t!��-* t�- u�F�F�ڊ�^&8u��^&�? u�^�? u� �+���]� X�EU���؁�V�v�e��~ t�v��WPj
�W������v��WPj �W�����u�� P�x���������vhj j j ���w����ǆ��  �#�vh
P�F�P���w�^�Ķ��&�@@t3��������9���vo�~ t��vh
P����P���w����P�������P������F� RP�o�����P�e�����P�v�U��t��vh�v
j �������w�������^MM��]M� U���
�. 9Fty�F�. �vhj j j ���w�F��vh�v��F�P���w=��u;�t;�vh�v�j j ���w�t �d
�~F��F��v�F�Pj �'�w�F���v�]�w��]� U����F�F���?	t�F�^�? u���+F���]� U����v����F��v�v�v���F�P��K��F�F�`�v�F+F�P�v
j j j �v�v�j j �HO��F�@)F��~� ~6�F�@F�FP�i��F��v�vP��K��F��^�F�F�F�~� u���]� X�EU���؃�WV�^&�G
�F�&�G% �F�&�O�N�~ t�tQj�5�wRP��M��v�j��v�j�5�wRP��M��v�j�5�wRP�N��^&�u��v�j j j�Ì� RPj j j j j ���ǚHO���&�@�F�X�+����^&G�F�>.  u�9F�u	�~� t�� �~
�uw�Ft�F@t�F
 �Fp�_�F
 �X�v�?���^�^���F�� �Ft�F
 �-�v���t�F
  ��v���t�F
 ��F
 �F�^���~ t�~� t���F���F�  �v��F�P���+���+F���P�6~�6��6��F
�.~P�v�h� j ��K��d
~F�� t�F�u	�v����v�j�"N��v��v��+���+F���P�v�v�v��z��v�j�"N��^&�Gt�v�Ì� RP��w�~� u� �~ t� j�5�wRP�z��F��tp�F�V �~���ڥ����v�hj j j ���wF�F��^&� t�v�h&�GHPj j ���w�t��)F��v�F�P�vꚈ�w�v��H�^_MM��]M� U���vh�v�F�RP���w�vh�vj j ���w�vh�vj j ���w��]� X�EU���؃�V�^&�G���F� �~ u�j�FOw�}�F� �j�FOw�|j�FOw�}�F�  �d�^&�w���F�F�^&9Guz&��u�?�~ tP&�w��% �F��QPh
&�w�F�P���w�v��WPj �W�F��u�� P�x�F�V����^�&�@% �F��v����~� u�� �~� t�v�j��&�F���F�  �~� tt�^&�w��W;F�uc�^&�G=��tW&�wh
P�F�P���w�^&�w��WPj �W�F��teP�x�F�V�F� RP���F��v����~� u;�v��WPhj j j ���w�^&�w&�w&�w
��Z/;�t� �+��F��v�v�����~ t
��P���w^MM��]M�
 X�EU���؁�(�~
�u��vh�v
j j ���w�����t�F9u�h�~ t3�vh
�v
����P���w�v�v
�M��u����P���up�/�v��WPj �W�����u�P�x���������vh
�v
�F�P���wĞ��^�&�Gu�GP���u�������� �������vh�v
����P���w�v����P�(w����PP����P�>w�~ to�v��w�������� tǆ�� ����Pj�j��w�ǆ�� �����5�wRP�z������t��������QP���w������H��v������w��v����Pj �'�w�v�]�wMM��]M� U����F� ���F��u+��*��  �F�P���w�F�
 hB j j�+��V��t�P�x�F�V��v��F�P�(w�v��F�P��w�F��V��^�&�G&�W�F�P�v��v���w= ����^�&�G&� ��V����l��X�P��^�Ph ����V���f�P���@�F�F�j PjB����\��tJ��f�P��V��x�F�V�F�HHRP�l���V����F�F��v��X�Ph���F�t�z��v�h3��V�j j ���w� ��]� X�EU���؁�@V�F�  +��F����vh�vPP���w�F�j�FOw�}f�vh�vhj j j ���w�F�Pj j ���w�F�j�FOw�|�vhj j�j����w�vh�v��v��v���w�vh�vj j �Qj�FOw�}�~� tǆ�� �=�v�vj�!��0�~� t�F� �#�vhj j�j����w�vhjj �v���w�~ u�v��WP�~�v�FP�tw�v�FP��w�F�P�F��+�P�F
��+�P�Q�R�=w�v�Ԩw�F� �F�2 �F�Pj j j �vҚD�w�t
�F�P���w�~� �F� ��N暗�w;Fta�F���(w�~�u{�~� t#�vhj j�j����w�vhjj �v���w���� t�v�vj � ��vhj j�v���w�� �~�t��~� t�S��F�P�v��vښ�w�t�<��y��vhj j j ���wHt�4�~ t%�vh
�v����P���w�v�v�S�% �F��w�vj �W�F�P�x���������vh
�v�F�P���w����P��������F� RP�o��^�Ķ��&�@��% �F���@t�v���� �p�v����~� t�F���}����P���t�F�������P���tS�F��hB j h� �+�F��t?P�x������������P�M��������� RP����P�o��v����F��� -��F��� /�vhj j j ���w�F��tv�N���wP�v�v��v��v����P����F��V��~� t�v�G���~�PRu�~�NTu��  �vΚK���~�FIu�~�LEu�v����vΚ_�v�w�t�vj����  �~ u�v�w�t�v��WP�~� ^MM��]M�          U��F*�=| t:w(,"t4,t+,t,,t#,t��|��~,t��t,t�~ v
� ��F�+���]� U��WV�vV�������~��ހ�:u�G� ��^_��]� U��WV�v����<\t�<:u�| t�D��F�< u��^_��]� X�EU���؋^�? t��F�^�? u���\t�\�F��F�^�?\t��vS�o�MM��]M� X�EU���؃��F�F���?:u�\u�G�F�F@�F��F�^�? t
�?\u؉^���^�� MM��]M� X�EU���؁�V+��F���������P�vh������P������P���ǆ�������^��?\u����\u�^�G ǆ�����^��? t�:u���% �F��F���� �F�P��������u)�F�������Pj�
��u���������  �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                8    �     U                          ,    �   PUU                         8    �  @�UUU           P        QUU ,    �  UUUUUU          TU         hU 8    �   @UYU�         @U�        @U ,    �    @P	          hUUU      @EU 8    �                  UUUU    @TUU ,    �                  `�U�    TIUVV 8    �                   %T*       �P� ,    �           U                   8    �         QUUU%                   ,    �          hUU%                   8    �          @UU%                   ,    �         @EUUUQ                  8    �       @TUUUeU                 ,    �        IUVV�JaZ                 8    �         �P�*                    ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �       ���                       ,    �       �Y�*                      8    �      �jVf�                     ,    �      jVU�Y
                     8    �     ��UQUi)                     ,    �     �ViT��                     8    �     �UU PT�                    ,    �    �j�EAP��
     ���            8    �    �VE U��     �Z�
           ,    �    �YU  PZ�   ��Zj�           8    �    hU  @i�
   ����U          ,    �    �U  Q�e*   h�YeU	          8    �   �f�U   ���   �U@%          ,    �   �Z)T    Z�
 �jU  �          8    �   �� @Phi* �Z�EQ         ,    �   ��     T�V� �jJ  @	         8    �   �e    �Z���@  %         ,    �   jeT    QUZ����   �         8    �  �jU    @�V���  Q         ,    �  �fT     PUZ�VJ   @        8    �  �V  @ @Aei�UY   D	        ,    �  ��VA    P���ZZ  @ %        8    �  ��T      @��   A�        ,    �  �i      @U��jT    P       8    �  jZ     D�Y�@    P	       ,    �  �fQ     PQZ�F      @%       8    �  �iT      D EZ�
      �       ,    � ��ZEA       U��) @  T      8    � �VVQD       T�V�       T	      ,    � ��      @TQe�R     %      8    � ��EE@      @@T��J      @$      ,    � �VFA      DP�V�
     @�      8    � �VR       P ET��*   @  T     ,    � �eQ          UY�)      @	     8    � h%A    UiY�@     	     ,    � j)      ATT���A      $     8    � ZP     ���       �     ,    ��ZYU    @ @@E�V�j @    P    8    ��V� @E@@D@A EUYj      D    ,    ��Z�UUQ EPTUUUTPe�PTTT
    8    ���DUT�EeEi�UjUe��T�F�UUU�QQ
    ,    ��VT���Q�U����V���V�Z�����     8    ��eU*(U��(UJ(V*(�**(f�(    ,    ��f�F�"VB�b�B�"J���J�"�A�� D     8    ����*(j*h&*h�*��*(�*�    ,    �j��R
�R��R
�R��R
�R��B     8    ��f"��  �� "��  ���"��  �� !�    ,    ��U��$���$���$���$���$���$�       8    ��f)�$�(�$�(�$�(�$�(�$�(�$�       ,    �����%���%���%���%���%���%�       8    ���"��% ��% ��% ��% ��% ��%       ,    ���!�e	 �e	 �e	 �e	 �e	 �e	       8    � ���U��U��U��U��U��U       ,    �  @VU
@VU
@VU
@VU
@VU
@VU
       8    �  `Z�"`Z�"`Z�"`Z�"`Z�"`Z�"       ,    �  �TU�TU�TU�TU�TU�TU       8    �   �� �� �� �� �� ��       ,    �          T@  T       T       8    �   P     PEU    U     PEU      ,    �  T                            8    �                                 ,    �      @           @          8    �        PTU          PTU       ,    �         T     PUU   T        8    �              @U           @   ,    �             PT                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    � TU                 TU         ,    �   TEA     @U         TEA       8    �      D  PUU             D  P   ,    ��       UE     @ @        UE   8    �&                UQ               ,    ��                                �8
   �
                                ��                                       �                                                                                     �        �        �        �     " ��  ��" ��  ��" ��  ��" ��  �� � �� �� � �� �� � �� �� � �� �� ��� �( ��� �( ��� �( ��� �(����
���������
���������
���������
�����������+���������+���������+���������+����~���_����~���_����~���_����~���_�����_�_�W�U��_�_�W�U��_�_�W�U��_�_�W�U���W�U�WU��W�U�WU��W�U�WU��W�U�WUu�}]�_UU_u�}]�_UU_u�}]�_UU_u�}]�_UU_}�Wu��WU�W}�Wu��WU�W}�Wu��WU�W}�Wu��WU�W]UW���UU�U]UW���UU�U]UW���UU�U]UW���UU�U]UWu�����U]UWu�����U]UWu�����U]UWu�����U]U_u��_��U]U_u��_��U]U_u��_��U]U_u��_��U}��}��Uu�U}��}��Uu�U}��}��Uu�U}��}��Uu�U�UW��Uu�W�UW��Uu�W�UW��Uu�W�UW��Uu�W��U�}�UuU���U�}�UuU���U�}�UuU���U�}�UuU�W�U]w�WU�W�U]w�WU�W�U]w�WU�W�U]w�WU�U�U]w��w��U�U]w��w��U�U]w��w��U�U]w��w��U�W_������U�W_������U�W_������U�W_������Uu�W�u����Uu�W�u����Uu�W�u����Uu�W�u����W}�W�]�W��W}�W�]�W��W}�W�]�W��W}�W�]�W��_]U_W_UW��_]U_W_UW��_]U_W_UW��_]U_W_UW��  �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �     P                           ,    �     T                          8    �     U                          ,    �   PUU                         8    �  @�UUU           P        QUU ,    �  UUUUUU          TU         hU 8    �   @UYU�         @U�        @U ,    �    @P	          hUUU      @EU 8    �                  UUUU    @TUU ,    �                  `�U�    TIUVV 8    �                   %T*       �P� ,    �                                 8    �                                 ,    �           U                   8    �         QUUU%                   ,    �          hUU%                   8    �          @UU%                   ,    �         @EUUUQ                  8    �       @TUUUeU                 ,    �       TIUVV�JaZ                8    �    @   �P�*          P        ,    �    T                 T        8    �   @VU               @U�       ,    �   UUU)               hUUU       8    �  @UUUU              UUUU      ,    �   ZVY	           U  `e��       8    �   �jh          TPUU   )�
       ,    �                 VU�            8    �                  �              ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �    X                            8    �   �j                           ,    �   �j                           8    �  ��Z             `             ,    �  ��ZU            ��            8 @  � ��ZU           ��            ,    ����VU           �jU            8    �U���ZUU          ��jU           , @  �U���jUU         ��jU           8 @  �U����UUU      � ��ZUU          , @  ������VUU     `U ��jUU          8 P ��U����VUU
     jU���UUU          , @@��U����VUU    �jU����VUU         8  ����Z��j�UUfY  @�jU����ZUUU         ,  Ph��$��ZQ�YUV	 U�������ZUUU        8  ��E��V�UeYeU�U��V����ZUUU
        ,  �B�VifY�VUUUUYU���V�����UUU        8  e�ViUfU��DQU����Z�j��jYUUfY       ,   T���E�UUjUT��j��V�PeZZYUV	@     8 @ �TEYUQUUdTTX�Z�B�UePUdYeU�    ,T T�UUQETAUeQ@�@�  fQh @ TYU)    8Q@Q�U@ @UB   @�@
PTPUPUE�T   ,@ �      P      P  � UT T   8P @�    P                @ET   , @ �               @    T @   8    � @  @ @  @ @  @ @    ,  �  @    @          @    8 @ �@    @    @ U  @      ,  �           P@        8  � @     @    @ @   @     ,@  � @     @    PT    @     8@  � @     @    @P   @     ,@  � @     @     P@  @     8@  � P     P    T@  P     ,P T�@ T T@ T T@  T@ T   8  � P     P    @@P  P      ,    �  @  @   @  @  P   @     8 @  �  @  @   @  @  UA A   @     , @  �  @  @   @  @  AAA   @     8 @  �  @  @   @  @  @ P@   @     , @  �  P  P   P  P  P  P   P     8 P  �  P  P   P  P  AU TP   P     , P  �P    P    PPU  P      8  @� @ @  @ @   U@  @ @   ,@ @�    @     @    @      8  �     P     P     P   @   ,  � P  P   P  P   P  P   P  P    8  P �    @    @    @       ,   �    P     P     P         8   �@ @  @ @  @ @  @@U     , @ �P  P   P  P   P  P    T@@   8 P  �T  T @ T  T @ T  T @ P PA   , T P�   P    P    P    P 8  P�   P    P    P    P ,  P�T  T P T  T P T  T P T  T P T8 T @�T  T @ T  T @ T  T @ T  T @ T, T�������������������������������������������ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ��VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU�VUU媪�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ�ꪪ����������������������������������������������������������������������������������U�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[UU�[U�����������������������������������������������������������������������������������ꪪ�ꪪ�ꪪ�����ꪪ�����ꪪ�����ꪪ��UUU�VUU�UUU�VUUUUUU�VUUUUUU�VUUUUUU�VUUUUUU�VUU�UUU�VUUUUUU�VUUUUUU�VUUUUUU�VUUUUUU�VUU�UUU�VUUUUUU�VUUUUUU�VUUUUUU�VUUU  �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �     P                           ,    �     T                          8    �     U                          ,    �   PUU                         8    �  @�UUU           P        QUU ,    �  UUUUUU          TU         hU 8    �   @UYU�         @U�        @U ,    �    @P	          hUUU      @EU 8    �                  UUUU    @TUU ,    �                  `�U�    TIUVV 8    �                   %T*       �P� ,    �                                 8    �                                 ,    �           U                   8    �         QUUU%                   ,    �          hUU%                   8    �          @UU%                   ,    �         @EUUUQ                  8    �       @TUUUeU                 ,    �       TIUVV�JaZ                8    �    @   �P�*          P        ,    �    T                 T        8    �   @VU               @U�       ,    �   UUU)               hUUU       8    �  @UUUU              UUUU      ,    �   ZVY	           U  `e��       8    �   �jh          TPUU   )�
       ,    �                 VU�            8    �                  �              ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,    �                                 8    �                                 ,  DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD����������������������������������������YUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����������*                  ���������������������?                  ���������������������.                  ���������������������.                  �����������������ꯪ/                  �������ꯪ����������+                  ���������������������.                  ����������ꪺ��������:                 ���������������������:  @             �����������������_���:    P        P  �������_���_���������_   � P   � �_�����������_Z�_��뗥PZ P���PZ P� ���_Z�_���תj�����i}��i����jA��j����jA��j�����i}�����Zj������Zj�����Z�����V���j�������j��jiiY��Z�jii���Z�jii��VZ�jii���Z�jii���Z�����j�������j�������j�������j�������j������j���Z���j���Z���j���Z���j�Z�Zi��j�Z�ZZ�������������j����������Z������������������������j��������������������������������������������������������������������������������������������������������������`mdfv8�^�jEv7�bmd8�f�v�v�&�amefv8�_�jEv�cme8�g�v�v�8``xآ��� IՅ �I� �-d ��� �� ������ ��Ս ���� � �� ��L� �� �ߥ��� (�L"� \�d� �8���i
�� ������� I���d�dd���	�p�
 ��dddddddddddddd'd(d)d*d?d@dE�d�F�dH }� }� }� }� N� ��h:��J�B������ �� N� }� )� � �� �� �� @� v� M� �� �� �� (�� �0�0hL�ĥ��8�����`��� ����`����������	���,���Ņ� L�P �����L��            Game Over             �p�� ���L� �ũ���������	�������Ņ� L����
�� 8� �� ��P �����`            Stage:??              �J�8���� H��d���������8��嚅� f�d���������8��嚅� f�hɠ��`����P�����xH�P���� [�h:��`��
��
��^�����ɪ� D� �ƭ  )����
����
��
���` ��)i�� ��)?i���P���01����������� ���� ��):�� ����	 ��)::�������`d������ ������` ����}�����}���ɠ�Z��	}�����}����x�C�
}�	��	� }����� L��)
�� ǅ��!ǅ���JJ� ǘi/���Q���ȥ�Q���`^` < � ��  )�� ���  )��� ���  )��� ���  )���`��������E
��E�F��F� )����`��L9Υ�L~ͥ���nLȤ������ǐ	d�#�L�ϥ)
��Dȅ��Eȅ��������LȼMȢ �����d��J���������dd`�ȴ��dP   �Hȅ��Iȅ��������PȬQȢL����Jȅ��Kȅ��������RȬSȢ �LL�T�zɮ��*,	(	(� �?  � ��  �*���  ��� ���kY ���kY ���j�. ��몾. �*뫪: �&�ZU) ��vu% �6���- ���uu% ���UU� ������ �껪��������િ�������������������������������������������������������������������������������
���������������������������������  ��   � �   ? ��� ���� � �?  �* �?  �� ��  ����� ���� ���f �����= �*���> �&���� ����� �6���� ������ ������ ������ ���� �����: ઺��� ������ ������ ����������������������������������������������������������������������� ������ ����� ������ �����< ����< ����  ���  ���  ���  ��� ? ���  � ���  ��   ���    ��*  � �
�� ��? �*�� �; ���� ��� ���� �Z� ꪬ� �Z�躬* �ڶ��/ສ���������������VU��?����]]��?���j��?���j]]�����jUU������������������ �������? ������� �������  ������
  ������
  ������
  �����  �����  �����   ��﫺*   �����   ��着   ����   �����/   �����/   �����/   ���?   �� �?   �� �?   �� ��  ����
  ����  � *     � (     �*  �   �� ��?   �� �;   �� ���   �� �Z�   �� �Z�  �* �ڶ  �/ສ�  ������  �������
 �������/ �������� �����������ꪫ������������������?��������?��������?���������������
��������
��������
�������������������� ����﫺* ������ ����着  .����   �����/   �����/   �����/   �� �?   �< �?   �< �?   �< ��  �� ��
  ����  ��
     � 
     ��d��}�������ͅ��
��L�                       ��* �<    ����^  ������V	  �������:(�������������������������������������������������������?���������?�?������������?�� ������   ���ɀjɀje����ϐ��υ���I�i ɀj� �ϩ����΅��������	�$�L� �
 �? �
 �+ �� �* �.��� ����*�����+�kY��.�kY.��
�j�.����ꪾ.�����뫪:������ZU�������vu��?��������?����uu��?����UU������������������ �������  ������?  𿪪��  𿪪��   𿪪��   𿪪��   𿪪�*   �����+   �����
   �����   �����    �����   �����  ������  ������  ��??��  �����  ����*  ��
 ���  ��
 ���  loru��Ѕ��]���8��鐅���� ���'������8���0����� �����`� e� ��"d#��$8�	� JJ�r8�
�"�odn Q�v�%�w�&`�	���
����L�ԥ
�s�L�Х�L~Ф�Z�� ��z��LqХ
)�L��ƠƠƠƠ�L��ƠƠƠƠ�L�Ф����e	�	���e
�
�s�d�s�
�L�� ���������������������������� ���� 	
d�	)i
$0i�L�нх��х��ѼѢL�'у���W���'Ӄ���R� ����4�������_�?WW�]UU�]AP�WqS5_Ve=|�U U0 �* �Z1 �[ � �� �~1 �^ �*5      4    ����4������?�}}�]]?wUU=wA=_�q5Y��UV�U �
% �V9 �V �:4 �* �.4 �� �n1 �j �
    ��4 ��>����4�����w�7�_]��UUu7�Aup5M�7�UU� WV�P�Y=TPAU}@Zo] U�k5 T�� @��6  ��  ��6  ��  ��u   5\   4  @ ��$ ��>����$�����w�'�_]��UUu'�EEup5M�'�UU� �Y� \V=T @U}  ZoY @�k% P�� P��& P�� P��& @��  ��e   5X   $  @ �? ���������?���?����wUUuwAu\�M�|Y���UV= X� @��PU�P��P��P��P��@����^  �T @T �� �����������U��U��U ��W�W��_U	�U	 i ��  �V  �V  �Z@�nP�� �� ��  Tj   T   ��  ��?  ��� ��� ��_� ��_u ��_ ��}� �uY ��U�  �WU  �   X   V   W  ��k  @�k P�� P��  ���      T     �? ���������?pU��pU�� U��0���T��?`U�?`U�@i�  �
  �
  �. @�~ P�oT����  �� @�       ��  ��?  ���  ��� _�� ]�� P�� S}� e]� VU� U��  T�  �%   �   ��   �V @�[ P�z  ��  ��  P  @T      ��8�������`e
�
�s��s�
� JJ)���ԅ���ԅ����L��R� �? ���������?���?����������������*��p��5P��P��P��P��P��@����^  �T @T         �� 0�?����������?���?���������������꼪���*�>@��@Uj@�j �^ �^@�j  	
�����`�	��
i�����LL�  �բ �բ�0`)@�Aڵ������"���օ��i �ک� �z�8����t��L��`����������������)?����u�ɠ�tL��ڵ������m���օ��i ��� ��`   <����������>�����?0<  0  	
 �� !� ��L٢ �'�'�'�'`� )�` ���������
���`��Lש�Lש�Lש�Lש��' ��)i�7t/ ��)?i0)��+`��'� 0����`)��`����H���H�
���ׅ���ׅ��+���/���7JJJJH�7



u3�3hu/�/ɖ�	�i�zhL�hht'�i�L������Q؁�PT���������?��?������������@�o  �  �  @   �* �>�������/��/����������տ�����������/���# ����� �* ���
���:�:Z���Z���Z���Z���Z���Z���Z���Z:�:Z���Z���Z���Z���_���   �    � ���?��<��������������?��?�� �  P   �   �
 ��( ��� ��� ૢ ૪ ૪ ��� ��� �U�U�_ �   P  ��'� �����`�+�^�/�_��b�c�	�`�
�a��d��e��f�gZ ��z�`�'ɂ�L|��`�  ٢ ٢ ٢�'0`�  0٠ 0٠� ���`�+�^�/�_��b�c� �`� �a��d�e��f�gZ ��z�`�Z� L�z���� �'ɀ�Ɂ�Ƀ�'Ʉ�=`�d�L���
eF�F�ɐ�ȅF� �'�i�L���;�+�<�/�= �٩P�7�8�9�:`8�/���/`�;�`�
�d;�L���;�<���=��� ���څ����L�     p�j�j��V��P:d@
o @d ��@	�P��:�Z�p�j �1  �   I� ��L���>�>)�` ���(�`� �?�?`����������?� �A���C`�  �ڢ�?tJ�5�A��ɐ�(�C��� )��A��)
��
ۅ��ۅ��i
���L���?`�A���C����1� )��C�C��)���H��H��)��ۅ��ۅ��i
�zhL�`V?�i
�L��"�B�b�Bۂۢ��ۢ�  E  V �p�vw����g��f< �  E@Vp?�|�v�����g|�f0 � E@?V����v���p�W�������;���/���>�
�T��P�* / ��;���/���>P�
�P�*�?�
@��;���/�+�>��
�?�*�� �  �ۢ�?0`�A�^�C�_��b�c�	�`�
�a��d��e�f�g �ð`���`�0`� ���"��� )��n܅��o܅���� ��#e��$e � ɠ��%e!�!�&e"�"ɠ�`d�L��vܶ���6� �? ������?��?��������������������?��?���� �?  �? �����o��0��4����o@����������o@����?��?0����� �?  �? ���������?���?����WUU�  �  �WUUի������?���?������ �?  �? ���0����?��?o@������������o@������4��0��o��� �? ��`��`��`�  ) � /ޭ  )� 8ޭ  )� �ݭ  )� �ݭ  )�O�  )�]`�	i���LLީ��	�
���
�
��p��
`�	i���`���	�
���
�
�s�N�s�
`d�
�s�A�	�	��9��	`����
�s�*�	�	ɐ�"���	`����`���%%0���
�` S�L�ޢ���� b���`��^��_��`��a��b�c��d� �e��f�g �Ð�������d����� ��	LL�`��=�9� �^�"�_�	�`�
�a��b�c��d��e��f��g �Ð��` ߥ )�`������ D�L�ߥ )�`��`������������ 8�:� ��L��d��  �� L����߅������� L�F�  ��H� ��h ��F�`������߅�����	��LL�Time:             Time Over             ������ 8� Z� ���* ��z����`��H)�&  � (�h�& `��H)�&   �h�& `Hژ��]
�h�Qh�P`�l�m� �lH
�� ��\�!��]� ����`l\&�4�B� �l� �����`� �l� �����`� �l�( ��������l`� �O�� �O��)�� ���:� ����"�� � � �( ����`dO v�!�:�����(��O��` ��O��`�(tO���!����Lv����X�Y� � �X�P��������]� �Z������`�a�b�O`�O�`�`��L�����a��a�`� �`�bm��a�]�
�Z�	�Z�� L��d㪵P�V�Q�W�`� �V0L�����L�����L������ �]����� l�V�bm��a l�L3���� l�V��V8��V�W� �WL3����L�����������}h㨹��V���W l�L3����- l�VH l�VH��}h㨥V���W������h�Wh�VL3����' l�`�`� �V�������Vi�V� eW�W�`L3���� l�VHȱV�Wh�VL3����2�`�)��:�� �� ��V��!�`�ZL�� l� l�L3�����`�`�)��)��� l�`L3�ɀ�(逼`�

��*��+��,��-� l�`L3�`����`㨹�� ��� �� ��  l� �V��!�`�Z l�`
��V�P�W�Q�`��������`�_��\��\�L�� �T���� �_L���� s�T��T8��T�U� �UL�

� s�T��!�\ s�	�( �
�) ��)�* 	�* L��   �V��W`�T��U`H���
�hJH��m�hnn���`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   �������������8��墰I�iƔƔ��8��声I�iƕƕ���日���������ė�L�0��Z�������� *���e���8��咅���e�����e���z���`Z�������� *���e���8��哅���e�����e���z���`Z�������� *���e�����e���z���`���O�H�� L�)���JJ��W�1���h=S����` U��0����?��������������� ���^�_�`�a �奓8*��� *����m^�^��m_�_�d���
&�m`����ma���������� ��8���^����_�������`���aƔ8�^�`�^�_�a�_�`�a��œ�Ly�`��Ŕ� 楓��������e�ɠ��� (�8���ɠ�ׅ� (�`��e�ɠ��� *�8���ɠ���L*�`�n�o� 8�nH� �o�h`H�nEn�n�I�i�hI�i ��$n� 8�vH� �w�h`H���v
�whJH��ew�whfwfv��v�w`�oEsH$o� 8�n�n� �o�o$s� 8�r�r� �s�s ��h� 8�v�v� �w�w� �x�x� �y�y`� �y�x�v���wFofn��xer�x�yes�yfyfxfwfv��`�n�oEo�oI�i��nI�i 8�(I�i`�n�o� �Hn�*�o��o�h*��`�oErH�rI�i�r$o� 8�n�n� �o�o ��h� 8�v�v� �w�w`��vJ�w�pn&o&p�p8�r��p&v&w��`�qEsH$s� 8�r�r� �s�s$q� 8�n�n� �o�o� �p�p� �q�q ��h� 8�v�v� �w�w� �x�x� �y�y`��vJ�w�x�y�t�un&o&p&q&t&u�t8�r��u�s��t�u&v&w&x&y��`���;���;�` 	$1@Qdy����n�o��r��s�w�v�n&o&v&wn&o&v&w8�v�r��w�s��w�v��**Er*�r&s���FsjFsj`��8��
��i
�n�



n`�n�o��n���o���
�o�n���n8&v&w���v�w`    
  ( P d � � ���@�E�n��o��p� ��p�n��n�o��o8&v&w&x����`        
    (  P  d  �  �   � � � @ '  N @� �8��@� 5�z R�r�z M�s��r V慘���~H�s V�8嘅����*�~��s V慘��h�r V�e����e��*�`�{ R�r�{ M�s�}�r V慘���H�s V�8嘅����*��}�s V慘��h�r V�e����e��*�}`�| R�r�| M�s�~�r V慘���}H�s V�8嘅����*�}�~�s V慘��h�r V�e����e��*�~`I�8i@�@�!���"

JJ(�I�i )?����(�I�i � `�� `����` 	"%(+.0369<?ADGILNQSUXZ\^`bdfhjlmoprsuvwxyz{||}~~8��倅���偅�8��傅���僅�� ��������������F�jF�jF�je�����)��e���������F�jF�jF�je�����)��e���Lf륍����F�jF�jF�jF�je�����)��e���������F�jF�jF�jF�je�����)��e�����e�����e�����e�����e���`�)�r�JJJJ�s��)


8�r�n��)�J8�s�o��)


�p��)�J�q��enfv8堨jEv.�nep8�r�v�v� ��eofv8塨jEv�oeq8�s�v�v�8``H�ZE����e����嶅��  E��� �� ����z�h@��+� �� �����m���� � � � �`
�
m�� �g�������`�,
� � 8� � 
�@@ 
��<� ( �  �S����P�  ���� �l���?�  �����  � � � � � � � � � � � �Ʌ��& ���d��?���n�n��� ���@&��@&�

���I�� _���L�� ���@�������4�'�����0e���� e������` U����


 L�
e�����`��X텪��텫` 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]H� ��hHJJJJ ��h)	0�:���H�Z��Z��Z ��z��z��z�h`8� d�
&�
&�
&�ip����e���� Z���� ��� � ���0e���� e���z����8���~�������`���H򅘦��H�F��	F�*F�*L6�F�*F�*F��	F�*F�*LI�F�*F�*F��	F�*F�*L\�F�*F�*F��	F�*F�*Lo�F�*F�*`        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d�  �U�LQ�� 8� ���������������� ��LT�`d�d�� Z�� ��z���Z歱�ƭ ��z�����`H 8�栥�I����hd�i��
&�
&�
&�
&�e�����e���� ��� ������������0������1������`������a������������������������	�������
���𑪠����櫠��� ������!������P������Q��ƫ`��������� d��C����� ������(���'e������0e��������`����.���n�������n����`���� 8� �����Ę���e������0e�����ƙ��`�? ����`���n`� �������������� �� ��L���?�n��� "������.�.�����n�n��� ����`��d�
&�
&�}�������e����e����nJJHJJJe����溼��n)�ȹ��������������d�h)��&�&�&�:��ڽ.�� �����ȥ����ȥ����ȥ�����e���������`�����.���n�������� L�nJJe����櫽n)
�����������d�
&�
&�}�������e����e����nJJHJJJe����溼��n)�ȹ��I������I������I�������h)��8&�&�&�&��i���H� i��ȅ�hi �ɐ��ڥ��å��ĥ��ť� �� ��1���ȥ�1���ȥ�1���ȥ�1�����e������0e������e�����ƼЫ�` ?�����������������         ?���������                 ?��'�M�y�l� � �� ���Ļ��`� d���d�)����
&�
&�� ���Ļ�楜) ��`� d���d�)����
&�
&�
&�
&�� ���Ļ�ड़) ��`� d���d�)?����jj��j)�� ���Ļ�奜)? ��`���`�ɪ��Õ�` @� @� @� @�        ����� ���@�����������L����  ��� ��� ��� ��� ���0e������e�������΢�� ��� ������� ������� ������� �������  ���0e������(e������e������Ч`��F�������F�������F�������F�������F�������F�������F�������F������`����H�


�hLE���� ��� E������ E������ E������ E������  E��0e������e������в`��� F�����F�����F�����F�����F�����F�����F�����F����` ����Ť��`��E�M  e�*��E���e���&�E���`���A���  :00*00)00*0( * ( * + * + * ( * ( * &( * ( * + * + * ( * ( * (���  &0)00(00(00)%#%
%#%� 0 %��H�����  6()(()(()(()(()(()*()(()*  (    (    (  )      (    (    (  )    ��  30 �O��!�������  8  00&0&000  00&0&000  00&0&000  00&0&0000  '0 ' 00  '0 ' 00  '0 ' 00  &0 & 0��  $0 �(����<�o���  :
 � ( )00( ) ( ) 00  � ( )00( ) ( ) ��  %0 $0	0$00$0"0$0	0$00$0�v�������  :�  �  � )  0 �  0��  '
00
00000�         ������  :$���  7$
�����  8  00&0&000  00&0&000  00&0&000  00&0&0000  '0 ' 00  '0 ' 00  '0 ' 00  &0 & 0��  $0 �(����<�o���  :
 � ( )00( ) ( ) 00  � ( )00( ) ( ) ��  %0 $0	0$00$0"0$0	0$00$0�v�������  :�  �  � )  0 �  0��  '
00
00000�         ������  :IO      SYS           (� ��  MSDOS   SYS           (� �  SACHEN_HO  (          fA      COMMAND COM            (�& �  WINA20  386            `��x�$  SMARTDRVEXE           @jY�  RAMDRIVESYS           @j�F�  EMM386  EXE           @j|~^� VSAFE   COM           h�t�,  MOUSE   INI           �Q�P   MOUSE   SYS           @j�qx�  VSAFE   SYS           h����{  PE      PIF           �I�6!  PE      EXE            `�/  PE2     BAT           i(\   PE2     PRO       �@�& L��������