                      	     �      �      �      �      �	      �      �     �     �     �     �     �     �     �     �                                       �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                         
           �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                  
          
               �      �     �	     �     �     �     �     �	     �     �     �     �     �                                 
     
     
     �     �	     �     �     �     �     �	     �     �     �     �     �                             
          �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                        
               �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                                   
     �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                                   
          �      �     �	     �     �     �     �     �	     �     �     �     �     �                           
     
          
     �     �	     �     �     �     �     �	     �     �     �     �     �                                      �     �      �     �	     �     �     �     �     �	     �     �     �     �     �     
                       
     
     �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                       
               �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                             
          

     �      �     �	     �     �     �     �     �	     �     �     �     �     �                                
               �     �	     �     �     �     �     �	     �     �     �     �     �                                      �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                                      �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                             
          �     �      �     �	     �     �     �     �     �	     �     �     �     �     �                                      
     �      �     �	     �     �     �     �     �	     �     �     �     �     �                                             	
          �	     �     �     �     �     �	     �     �     �     �     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     H�� �@�� �0�� � ��� ��� � �t ���u �u �r �t �q  [ϭu �r� /��u �� ����� �� /��� ���� ��� �u �u �r �t �q � ���  [��� �� �� �r �� �q �� �� � [ϭ� �D0 /�� ��� �� ����� �� /�u �r ��� �t �q �  �ϭt i�t �q  [ϭ� �q � �ϭ� 8��� �q  [ϭ� �� /������  /ꩀ�d  O�x��  ܜ� hLv� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       DDDDDDD         DDDDDDD         DDDDDDD@         DD@D@D@DD         DDDDDDDD         DDDDD         D@DDD@D@         DDD@DDDD         DDD@DDD         DDDDDDDDD         "" " ""         """" "          "" "  ""        ""   "    ""    ""   ""         "   " "  ""    "    """  "      "  """          "" "" ""         333333333         3033333         333 3333         3333330         33 333         333330330         3 33 33         303033030         33303333         33303033         333333333                  UPUP          UUUP UP         UPUUU         UUUP                   U    U    P   UU  UU    UU                UUUUUUUUU         "  " """         UU "" "   P     "  P  UU     P  """ UP ""         """"""          """" """          "     ""         """""""          " "   ""         UUUUUUUUU                  ff`fff         f`         f                                                      fffffffff         """"" ""         "" f`""         ""`""""         """" ""         f` " f       `  " fff ""         """"""          " """"""         """ " ""         fffffffff         3333333         3033333         33030333         33  3330        33 w 333    w    33  w3          3 3333030         30303333         33303 33         333333333                                                                                                              �   ��        � �        ���                                                        ���������         �������         �� ��� �  �  �  � ��  ��     ��  ����  ��     ��  �� ��  �  �      � �����         ��������         �������         ��������         ���������         DDDDDDD         DD@DDDD@         DDDDDDD         DDDDDD         DDD DDDD@         DD@ DDD    ``   DD@  @D   `f   DD   D@         DD@D@DDD         DDDDDDDDD         ������          	���   	�   �                      �����	���         	�    �       	��                           ���������         33033333         3303333         33330333         333033033         33333333         3033333         3 303330         30303333         33303033         333333333                                                                                                      wpwpwpwwp         wwwwpww         wpwpww         www  wp      w  wwwww w         wppp wwp    w    w wp  w     w   wpwp  wpw          w wwp         wwwwwwwww         ffffff         f` ffff           f f`fff         fff`ff`f`         f`   fff  ff     f   fff  f`      f  ffffff         fff`f`ff          f`ffff         fffffffff         "" """""         ��  � "   ��  � ""   ��"         """ """          """ ""  �         " "  ""         " " """          """""         " "" " "          ���������         D@DDDD@         UPU @U D   U   P U  UU    U   U  D  UU  UP         D@D DDDDD          DD@D  D          U  DD@ U  UP   @ UP UD         D@DDD@         UUUUUUUUU         ���������         ����	� ��         �� ������          ���	� 	�         ���	���	�           �� ����         ���	�����           	� ��	�         ���	�� ��         ���������8�`�����؎ �(�P�x���ȏ���@�h��������0� �	���$�-�6�?�H�Q�Z�c�l�u�~���������������ƀπ؀�������� �)�2�;�D�M�V�_�h�q�z���������������ˁԁ݁�����
���%�.�7�@�I�R�[�d�m�v����������������ǂЂق��������!�*�3�<�E�N�W�`�i�r�{���������������Ã̃Ճރ���������&�/�8�A�J�S�\�e�n�w�����������������Ȅфڄ���������"�+�4�=�F�O�X�a�j�s�|���������������ąͅօ߅��������'�0�9�B�K�T�]�f�o�x�����������������Ɇ҆ۆ���������#�,�5�>�G�P�Y�b�k�t�}���������������Ň·ׇ����������(�1�:�C�L�U�^�g�p�y�����������������ʈӈ܈���� �	���$�-�6�?�H�Q�Z�c�l�u�~���������������Ɖω؉�������� �)�2�;�D�M�V�_�h�q�z���������������ˊԊ݊�����
���%�.�7�@�I�R�[�d�m�v����������������ǋЋً��������!�*�3�<�E�N�W�`�i�r�{���������������Ì̌Ռތ���������&�/�8�A�J�S�\�e�n�w�����������������ȍэڍ�������  � @�� �` �@�� �`	 
�
@�HPX`hpx�������������                                                                ����  �����c�V�c���ci��cZi�����                                ����ZUU�j@��@��@�j@�ZUU�����                                �����UU��V���Z�
�j�R��TU�*U����                                ��������UUUU    UUUU������������                                ����  �����cffʣ���cffʣ���cffʣ���cffʣ���cffʣ��ɣ���  ��������*  ��*(�bUU�ZUU�ZUU�ZUU�VUU�VUU�VUU�VUU�VUU�VUU�ZUU��j������������������������ꀫVU��VU��VU��VU��VU��VU��WU��  �;  �  �������������RUU�RUU�RUU�R �R �RUU�RUU�R �R �RUU�RUU�RUU�  પ����\_�5WP�P� � � �WUQ�\Z�%��

                              �*(       �*(              (�*       (�*       �* �V�`UU	XUT%XU%VU�VU�VUU�VUU�VUU�VUU�XUU%XUU%`UU	�V� �*  �* �V�`UY	XPe%Pe%Tj�V���VY��VV��VV��VV��XY�%X�j%`UU	�V� �*  �* �V�`UU	XPU%�j%h��VVZ�VVU�VVU�VVU�VVU�XY�%X�j%`UU	�V� �*  �* �V�`UU	XP�%Pi%T��VU��V����je��Ue��UZ�X�U%XUU%`UU	�V� �*  �* �V�`UU	XP�%P�%���Vi��V���Ve��V�i�Vf��X�U%XiU%`UU	�V� �*  �* �V�`UY	XPj%��%Tj�V���VUj�V���VUj�V���XUj%XUY%`UY	�V� �*  �* �V�`�j	XPZ%PZ%���VYZ�V�Y�V���VfZ�ViY�X��X�e%`UZ	�V� �*  �? ���������:��:��諪
諪�諪�ꫪ�ꫪ�ꬪ�:���:������ �?  �* �V�`UU	XPe%PY%TZ�V�V�V�j�V�Z�V�V�V�U�XeU%XYU%`UU	�V� �*  �* �V�`UU	XPY%�Z%���Vej�Vf��VZ���UU��U��Xje%X�Z%`UU	�V� �*  �* V�  P�  P$D�@�P�P�@�D�P$�   PV�  �*      �� �WUpUU5\UU�\ �\ �\=��\ �p5��? ��� gf���?��� �       �? �U�\UUWUU5W @5W|5W|5W|5\�@����� �� �g� ��:  �?  � � ������������_U��p5@5_UU5\��7_�5z��UU ��   �  � � ������������_U�@5�p5_@5\WP7\}��p���UU �� �?   �? �W�pUU\W�5\��5WUU�kUU��_�p��s�\}}5�UU _�  �� ����� �? �W�pUU\UU5\W�5W���[UU�k}}��s�pڜp6��_�_������:��?<  <�  ?��� �� ���3���?|U�?|UU=|W=|W=�W3�UU W�  �?  p  �?     �  �  ��� �� ����w��WU�wUU�w�p��p���p��UU W�  �?  �?  �? ���������:�
0+  諌2꫌2ꫀꫪ�ꫪ��
�:���:������ �?  �? ���������:���:���+��諯�ꫪ�ꫪ��
�ꬢ�:���:������ �?                 �  �  ,9  l:  �:  �                          �   �  �   �   �   �   �   �  �  �  �  �  �  <                            �  �  [9  9  [9  �  �                   � ������>;�����)�b�/���Z�<�������0�� � ; < <   ?���_���eY�וV׼��>lUU9\AA5_AA�s1L�s1L�|1L=pP��W������:���                ?���_���eY�וV׼��>\AA5\AA5|1L=s1L�P�p�V���?    � ���=�Ue��U��U��WUV�WU��������pU��p���|e0��X�������� ���=�Ue��U��U��WUV�WU�������\U��\���\�0p�U5��� \-  �? � �|���gYUקVU׫�U�W�U�C�U�C���P��3SU53Sj5Tf5\Ub��� x5  �?     � �|���gYUקVU׫�U�W�U�C�U�C���3S�:3SU3Sj�Y=_%V�������        ?���_���eY�וV׼��>lUU9\AA5\AA5|1L=s1L�P�p�V���?���        ?�����몪�몪���?���:��:�2�:���2���
�������?���?���_���eY�וV׼��>lUU9\AA5\AA5x@v1L-z1L�pP���Z3����?      ?���_���eY��eY�|eY=\eY9\eY5�eY:���.����UU�sUU�UU?���:  ��     ��  ��> ����������������:,���:+����+���ꫪ��ꫪ��ꫪ��ꫪ��ꬪ��:����:������������ ��>  ��   ��   �  ���� �*����
�����������:� ���:� ���ꫪ���ꫪ���ꫪ���ꫪ���ꫪ���ꫪ���ꫪ���ꬪ���:�����:��������������� ����  �   ��    ��   ���  ���� ���� ���� ����������������������������� ����� ����� ������������������������� ���� ���� ���� ����  ���   ��   ��  ��� ���?�����������������?����?�����������?����������������?�����������������?����?������������ ���? ���  ��              ��� ����������������?����?���������������������������������������������������?�����?��������������� ����  ���   ��          ?    �?    �?    �?    �?   ��?   ��?   ��?   ��?   ��?   ��?   ��?   ��?   ��?   ��?   �����?�����? ����? ����? ���� ����  ���   ��   ��  ���?  ���� ���������?�����?�����?���  ���  �����?�����?�����?�����?�����?�����?���  ���  �����?�����?�����? ���� ���� ���?   �� 0  3  33 ��� �  ��� � �� ��� 0333 0  033033 0333 ���� �  ������� ���� 0333 0  0333033 0333 ���� �  �������� ��� 0 3 0  003033 0 3 ��� �  ������� ��� p 7 p  p 3pw7 p 7 ���� �  ������� ��� pww7 p  p 7pw7 p 7 ��� �  ������� ��� pww7 p  p 7pw7 p 7 ���� �  ������� ��� pp7 p  pp7p7ws7 p7s7 ��� ��� ��������� ���� ��� ��� ���;����; ���; ��� ��� �������� ��� � ; ��� �������?  �� ��� ��� ��� �����������������������                                              �? ��00 ��?�?������0� 0030 �������� ?00�0 �������� � �33 ��?��������?� 003< ���� ���� ?0030 ��0�� ��� 0� ��00 �������?���?                                                                                          �?�               ��               ��                ��                 ��                 00                ?� �       �d������ ��� kĩ7��s 
������� �ũ��v��2������ �ũh� y����~��4������ �ũh� ���	�� ����8� �P�����! ũ`���  � �ĩ��  � �۩ �	�d��h �� tǩ�	`��� �&����e 轀��f � ��eȩ �eȭu �
��� �eȩ �eȑeȑeȑe` � 7ĩ��<��4������ �ũh� ���	�� �x��8� �P�����! ũ`���  � �͜� �� 
�����e 轀��f �� �e�� �� ��ޜ�  ����c  �`��� � �	����(���x� ��� kĩ��0��>������ �� ܩ��(�h �� t� ܈г��	��� ��� `�� �s �0�
8���8�
�8�i�� `��� ���d  O� �ܩ	�� �o i
�o  �� � �ܩ��  �� � ��8�o �
�o �	��  �� � �ܩ��  �� ܢ <� ���p i�p ���  �� � ���p i�p ���  �� ����` 榜�  7ĩ-����:������ �ũ��F��2������ �ũh� y����Z��4������ �ũh� ���0��x��6������ �ũ0�����8������ �ũ�� ���t� �  ɿ� I������� �� �� �� ���  � ��` �� � ���� ��� ��� �t� � �ĩ��  �`��  ŭ�  ŭ�  ŭ�  ũ  �`��  ŭ�  ŭ�  ŭ�  ũ  �`�H�e ��f �N�g ��h ��� ���x��
��  ��  �� ��L1� � ��i����  � � ���i��
��  ���	��  �  g��  �� ��L1��x��	��  ��i��
��  ��  �� ��L1� � ��i����  � � ���i��
��  ���	��  � g��  �� ��L1����L=� ܩx��	��  �  �� ��L1��i����  � � �)�ɠ��i��
��  � � ����� ���� ��� �d�r ��q  [ϩ���#���	��	� ǩ���<������ �� �`��d���� �  ���\ � /� �������� �  ���= � /� �������� �  ��� � /� ����� ٪����e��g`ڊ
��k��k� ��`Zڭ� 
��k��k� ��z`�� �
�� �� �| � �  ��a���e��g� ٪�� ����� ٪��g�� I�� ����� /��| �� ����� �| ͦ Ш�| ��� �� I�� �����  � ��` 7Ģ �2��� ٪����ei���g���朻 ���� ��� �d�r ��q  [� ��` 7ĩ7��P��s 
������� �ũ	�� �x��8� �P�����! ũ`���  � �ͩ�c  �` 7ĩP���s  �ŭ  ���?����s � ��8��s �����s ���i�s �P���s  �� �ĩ��  ܀�`H�Z��� �� �å�� ��� �  �����  �Υ ��z�h`� ��I�����(���� i0�� �� i �� ����` 7ĩ-��
��:������ �ũ
��2��(������ �ũ��P��*������ �ũ(��d��,������ �ũ��x��.������ �ũ-�����0������ �Ŝ� �� �� �� �  ���L{�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ^�n�~�������������������.�>�N�^�n�~®¾�����������.�>�N�^�n�~ÎÞ�                                                                                                                                                                                    �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  HZ�H�@��m��������8��HJJH

�zh8����m�� ����ɪ�8��i0��i ����h�zh`H�i0��i ��_�����8������h`H�H�H�H�H������ k�h�h�h�h�h`xH�Z�ڮڦڦ� ��8��JJ�8���� � ����� ����h�h�h�h�z�h(`Hڭ  �� �������%���h`��������?_ow{}~���������������������H�  ����h`xH�Z�ڦڦڦڦ�
��`���`�� �â �  n�- �� n�- ��� Ā��iɠ���iɠ������h�h�h�h�h�z�h(`Hڪ)�JJJJ Ŋ) ��h`HZ� ��$�#�0i��:8�0��A08�7�i �Ȁ�zh`xH����L��Z�H�H�H�H�H�H�H��H��Hi�H�i �H ��8��JJ�8�����m��i ��������?������6� ��ȭ��h�h�� �������� ��m��i ���hh� h�h��0�� �����������ݬ�������
�h���h�	��h�h�h�h�h�h�h�zh(`�� �2��.HZ�Z�Z� ���������
������� �h�h�zh`xH�Z�H�H�H�H�H�H �à �ȍ���-�i��i �� � v�����m��i � ����h�h�h�h�h�h�z�h(`� �#��H���hH�Z�ڦڠ �������Lt�L}�L|���� ~Ȁ����LWȥH�H�Z�
�������������	8������	�� ��������*�e��i ��e��	i �	� �������	���8����	��������
�8����������������8h���h������
�������	��������h�h�z�h`ڦ
����	��.������`H�� �� h`�  � `H�Zx�H�H� H�H�H�H�H�H�H�H�H �Ì�JJ�NN� ����:����:�ȱ���:����:��8�����h�Hڭɀ�
��8�
���e�ȱ������e�������� ����+� � � nʍ �� �3� m������ n�ڮ� v�����
������P��r� m�����m ����8� � �8� �	� �m ��H n� v�h��,���� nʍ �� �� � n�ڢ ��� �� ������ �L,�h�h�h�h�h�h�h�h�h� h�h�(z�h`Z���z�`Hڦ��	���Q����h`�ڮڮڍZ�)���="ˑȱ�=%ˑ8����Z�JJ�����

������	��
�M��z�

�����JJ����z��ȭ�h�h�h��h`?���H�Z�H�H�H�F�H� �

�ȱ�z��Z�H��hHڍ ǭm����m����hhh�h�h�h�z�h`��d % 4 O B 
 z  0 7 p 
   � � ���7�kĺ���ŀŕ������t�~ȕȤȫ�n�v�)�                                                                                                                             ���  � <� 7ĩ  J�L �� J� 7Ģ��� �� � ��  <� 7ĩ(�� �c  ��� ��	 ���� �� �� �� �s ��c  �s ��L׬ �� ҫ�� �� �� �� �x ��y  xΩ �� ��u �P�p �v �t �{ �| �o ��  Gܜ�  l��# �� ��x �� 7��s L�̭� ��#x /魼 � ��� ��L{�L�̜� �d�� L�̭� �� }؜� x �ĭ� � Ǥ�� ���� �d�� �u �r �t �q  ~ӭ� �� ��XL!�H�ȍ� �ȍ�  �ĭ���θ �� /� /� /�ι �ݜ�  ���� /�h`�H�e ��f �s 
��X��g �X�i��h � J� � �g�e�����e i�e �f i �f �g i�g �h i �h ���Ωߍ& �� �� �� �2�� ��� �� �� ��  ����� ��� �s 
����m ���n `� �� �@�� �y �� �x �� �
�� ���  ��`�� �� �� �� �� m� �� �� �k �� �l �� 
��m�g ȱm�h �� J���g)���gJJJJ
���i�� ��i �� � � ���������� i�� �� i �� �� i0�� �� i �� ����� � �� ͨ �L��� �� ͩ ��k i�� �l i �� L��`H�Z�	썗 �	썘 m� �� �@�j � �i �r � ��i i0�i �j i �j �� ���q mi �i �j i �j � �� �
�  ���� � ��- �i��� ���i i0�i �j i �j �� m� �� �� i ��  ���� лz�h`H� �  [ϩ�� h`���  ��x�� �v  ��X�� �� G܀�� ���� ���� ����  G� /ꭀ �оx�� �x  ��X�� 0Lx���  ��H8� ���� �å�� ��� �y �� �x i
�� �
�� ���  ��h� l�X`��� x ���� �x X ��x�΀ �v  �� ��X�� �� G܀�� ���� ���� ����  G� /ꭀ � л��0Jx���  ��H8���� �å�� ��� �y �� 8�x ��� �
�� ���  ��h� l�X`��� �H�� ��� �x ��� �8��� �y i
�� ��� ���  �ΩH�g ��h �H���8���x� ��h�X��k ��l �k ���l ��x ��  s�/��� �����i0���i ����K� �܀��d� G܀����Ȣ�/�g�� �����g i0�g �h i �h �i0��i ����� � �� �� ����� �y  l�X /ꭁ � �L��`��� ��� �H�� �x ��� �8��� �y 8��� ��� ���  �Ω�h ��g x����H���8��� ��h���k ��l �y ��� X�k ���l ��x �࢜ e� e�/��� ����8��0���� ����d� �܀��K� G܀�� �Ţ�/�g�� ����8�g �0�g �h � �h 8��0��� ����8�� ���  l�X /ꭁ � �L��`HZ�� �� �� ���� ��� ��L����L�ԭ� �0�r ��i�q  �ԭ� � �L�ԭ� ��L����L����� �r � �L��8��q  �ԭ� � �L��L����"�r �0�8��q  �ԭ� � �L�ԩ� L��������C)��9�� �d��� �� �ܩ��  G� /�L�Ԭq � �L�Ԉ�r  �ԭ� � �G�@��<�� �d��� �� �ܩ��  G� /��q ��ȭr  �ԭ� � ��� �� ����� zh`HZ
��m�g ȱm�h z�J���g)���gJJJJ�� h`�� �� � �X ׀Y���UX�� �� }ح� ��C�  ���� /�7�� CՀ.�� �Հ%����� [ր���� }׀���� �`���  C֭� � �ܩ��  G� 4� [֢�� ��W�t � ��N��u  �ԭ� ��@ }׭u i�t  �ԭ� � ���ɭu i�t  �ԭ� � ��� �� �ĭ��� !�`���  C֭� � �ܩ��  G� 4� [֢�� ��Y�t ���Pȭu  �ԭ� � ��@ حu i�t  �ԭ� � ���ǭu i�t  �ԭ� � ��� �� �ĭ��� !�`�u ������ �	i�t  ��`���d  O� �� �ܩ��  G� 4� �ܩ ��  G� /��� �L׭p �P��y � �� m����p �d� ��8�p ��p  G� /����u ����� ��@�u i�t  �ԭ� � �- �ܩ��  G� 4� �ܩ ��  G� /ꭽ ��
�  ���� /�`���d  O� �ܩ ��  G� /�p �P��y �
� Zр� ���p �p  G� /�����u �u i�t  �ԭ� � � �ܩ��  G� 4� �ܜ�  G� /�`� �ܩ��  G� /ꭆ �� }ؠ��v �t �o �P��x � � �ЀL �ܭ� ��8�o ��o  G� /�v �.�� ���� ���� ���� �o  G� /� /��v �v � д�`� �ܩ��  G� /ꭆ �� }ؠ�o �P��x �� ЀF �ܭ� ���o i�o  G� /�+�� ���� ���� ���� �o  G� /��v �v �к�v �t �`HZڭt �� �p ��� ��%�� ��E� �o i� ٩��d  O� �؀'��#�� � ��o 8��Ο  ٩��d  O� ���zh`��J� !� ٭u Z��  ��z�� � �L~�x ��X�� ����L{٭� ��L~�� �i� ـ�� !� ٭u Z��  ��z�� � �L~�x ��X�� ����L{٭� � �L~�Ο 8��� ـ� �`��k��k� �`Z�� H�� �� �� �� 
�����e 轀��f � �e�� ���L������ɿ���	��0��0�0�ȱe�q ȱe�r ȱe�{ ȱe�| ȱe�~ �u �r �L��8�r ����| � � �q �0}8�q ��u�{ � �n��� �  �ܭ� �	�i�0���� �A�� � �.�� ��'��� ��� �{ �| �� �eȑe��eȑe�d�� ��� �� �  �ܠ �� �e��~ �e��� ��� �L�� ��h�� z`�  �ڭr ���r �r ��r �r ���r �{ �|  �ܠ �� �e�ȭr �eȩ �eȑeȭ~ �eȩ �eȑe`�s �0�
0�0��
������� `x�� �� 
�����e 轀��f � �e�� ���k�� �� ���ל� �� 
�����e 轀��f � �e�� ��3ȱe�q ȱe�r ȱe�{ ȱe�| ȱe�~ �� H�� ��  ��h�� ��� �� ��H����� �� �q �u �r �{ �| �~ �  �ܠ ��eȭq �eȭr �eȩ �eȑeȭ~ �eȜ} �eX`�  ������  � ��`�� ��� �� ͻ ��`�� �� ���`H�� H�P��  /�h�� h`H�� H����  /�h�� h`HZڥH�H�o ��p ��� 
��W��W���	 � �ĭ��������� h�h��zh`HZڥH�H�o ��p ��� 
��W��W���	 �h�h��zh`�H�H�H�H�� H�� H��� �z  0ݩ ͥ �" �ݩ ͥ ��� � �ͯ ��ͮ � �߀�~ h�� h�� h�h�h�h�`�� �y �r 0[�-8�r ��L�ݭ� �| 0L�ݩ�� �8��| m� �z �r��� �� �| 0�8�� �| ��T�z �R8�| � ��Fi
�r 0;���� �| ́ 0�(�y i	�r ���� �r 8�y 



m| 8� ���� `�� �H�x �q 0Q�x 8�q ��0L�ޭ� ��L�ީ�� ������ ���� �



m� �� �8� m{ ���Fi
�q �0?�{ ̀ 0�� ��0��� �q 8�x �	��� ���� �	



8� m{ � �À�� h�`HZڭg H�h H�k H�l H�� H�� H�� H�� �� �� 
�����e 轀��f � �e�� ���L��ɿ������ȱe�q ȱe�r ȱe�{ ȱe�| ȱe�~ ȱe�} ȱe�� �� ���� � �L ��������� �f�
�8��  �� �ڜ{ �| �} �u �	��r ��r �t �	��q �/�q �*��  �ܭ} � � � B᭾ ������
ɿ��  �ܠ �� �eȭq �eȭr �eȭ{ �eȭ| �eȭ~ �eȭ} �eȭ� �e�� �� ��L��h�� h�� h�� h�l h�k h�h h�g �zh`�� H�� H� �~ �j�~ I�~ �� 
��%�i�� �%�i �� �z 

m� �� �� i �� �z � �� v�������$�� i�� �� i �� �i0��i ��^���h�� h�� `HZڜ� �� 
�����e 轀��f � �e�� ���7���3ɿ�/��+ȱe�q ȱe�r ȱe�{ ȱe�| ȱe�~ Z�  ��z�~ �e�� ��� Т�zh`HZڜ� �� 
�����e 轀��f � �e�� ���=���9ɿ�5��1ȱe�q ȱe�r ȱe�{ ȱe�| ȱe�~ ��Z��  ��z�~ �e�� �� �М�zh`�} � �(�� �� )�ɐ��� ɕ��� �ɔ��� �)�� �o ~ӭ� ������R�� ͇ ��� ��  ~ӭ� ���:�� ������� �������� ����  ~ӭ� ������  ~ӭ� ���L䭆 �� ����} �� )�ɠ�L�� �歾 ɿ��������
�L�} ����} L䭾 ������� �i��� �b�� ������� �P��� �I�� ������� �7��� �0�� ������� ���� ��� ������� ���� �� H�� ���� �� � ��� 

m| �| �0�| �r �| �} L�����3�| � ��r ��| �� 
�� �| ͑ �| �} �
8� �| �} L����7�| � ��} �} � �t�r ��| �� 

�� �| ͑ �| �8� �| �N)��(�{ � ��q ��{ ͑ �{ �} �,8� �{ �} � ���{ m� �0�q �{ �} ��{ �} h�� �| �歾 ��r�� ɤ��r � ����� �]�r �Xɥ��r ������ �F�r �Aɦ��q � ����� �/�q �ɧ�&�q ������ ��q �r �q  �ԭ� � ����� `�� �0�7�l�	�1��%�� � ��r ������ L5�r � ����� L5�� L5�r �u ����� L5婔�� L5�q �t �
���� L5�L0婖�� L5�r �u �W�' �孇 � �I���C)���� )�� L5��� L5� 歇 )������ �� �m�q �t ���� L5���� L5�q �t �H# {�q i�t ��� ����� �/��� �( M��t i�q ��� ����� ���� ���� `�� �� 
�����i 轀��j � �i�� ɿ��� �� ����`�� H�q H�r H�{ H�| H�~ H�� �� �� �q �� �r �{ �| �~ �  �ܠ �� �iȭq �iȭr �iȩ �iȑiȭ~ �iȩ�iȭ� �ih�~ h�| h�{ h�r h�q h�� `�� ��.�q �t �& 6�� ����� �q �� 8�r ��� ����  c�`�� ��.�q �t �& 6�� ����� �q �� �r i�� ����  c�`�� ��& 6�� ����� �r �� 8�q ��� ����  c�`�� ��� 6�� ������ �r �� �q i�� ����  c�` �� +�`�� � �s�r �u �L*�q �t 08�t �!��V�{ �v N��t 8�q ��A�v �{ 9�� ���	��0�0��� ��� �� � B�
�� ���d  O�} `�� �� �� ��L.�iH
�����i 轀��j � �i�� ������ɿ��
��0L'�ȱi�� ȱi�� ȱi�� ȱi�� ȱi�� �ȱi�� �r ͚ �L'�q ͛ 0!8� ���� �'��L'�{ ͜ �L'魛 8�q ��� �{ ꭿ ��L�譾 ��*�	��� �	�L��HFL���0	�� �08��� �	�(�-� hL.魌 ����� ͈ �L'�	�� hL.� ��hL.魇 ͈ �L'�q ��!�q �q �r  �ԭ� � ��{ �| ���} L'魋 � �����r �
0��� �r � ��r ����� �r ����r ���� H�q H�r H�{ H�| H�~ H�� �� �� �q �� �r �� �{ �� �| �� �~ ��  �ܭ� ���� �ڜ  �ܭ� � �i��~ �ih�~ h�| h�{ h�r h�q h�� �� hL4�`μ �� � � t�� ̥`H�� �����
6m� �� �
008�
�� �� �� �
0 8�
�� �� �� �
08�
�� �� ��� �٭� �� 07��� �� �� �� �� �� �� ��� �� 0��� �� 0��� �� 0�ݭ� ������� �
�� � �β h`�� � �,�2�� �� � �Β ���� �� �� W��
�� �� ��`��  �ĭ���� ���`HZڮ� � ����� ���� ���zh`Hڪ��




�� ��)� �& �h`�8�`��� �`�i`��i �`STAGE  1$STAGE  2$STAGE  3$STAGE  4$STAGE  5$STAGE  6$STAGE  7$STAGE  8$STAGE  9$STAGE  10$STAGE  11$STAGE  12$STAGE  13$STAGE 14$STAGE 15$STAGE 16$STAGE 17$STAGE 18$STAGE 19$STAGE 20$YOU ARE VERY LUCKY$YOU ARE BREAVE$AND CLEVER$THE BUBBLE WORLD$IS SAVED$HIGH SCORE$YOUR SCORE$CONTINUE$END$GAME OVER$PRESS START KEY$HURRY UP$��������������������������'�0�9�L�[�f�w��������!AB>�6����,�n����4�v�����~����D���ȕ
�L���Ж�T���ؗ�\�����"�d����*�l����2�t�����:�|��� �B�|���|�����L�����t������آ t ���d���� � �����������  ��� � �� � �� �ߍ& ��"  7ĩ�� d
�� ~�L`�H�Z�  ��xL{�� � �� � �ε  z�(z�h@H�Z�' )��� � �ζ �� � �η  �ޭ�# �$ �% z�hX@� � � �  �� �� � � � � � � � �* �W �^ � ���X �b `H�Z� ���%�; � ��4 � �5 �  ��; �; �6 � �� ���%�H � ��A � �B �  ��H �H �C � )� ���X� ���� � �� � � �  P� ����- � ��& � �' �  ��� � � � >��- �- �( � �� �� r�z�h`� �� ȱ� ȱ� ȱ� ȱ� )
���� ��� � )0�" ȱ����X �b Ȍ � �  � � �L(�!  �� �� � ��! ��Ȍ! � ���1 �2�4 ȱ2�5 ȱ2�6 ȱ2�7 ȱ2�8 )
����9 ���: �8 )0�= ȱ2����X �b Ȍ1 �; �< �6 � �� � � �d )����� �>  )�`�> �?�A ȱ?�B ȱ?�C ȱ?�D ȱ?�E )
����F ���G �E )0�J ȱ?����X �b Ȍ> �H �I �C � Ш� � � �d )��@З��� �1  ��# �$�& ȱ$�' ȱ$�( ȱ$�) ȱ$�* )
����+ ���, �* )0�0 ȱ$����X �b Ȍ# �- �. �( � Ч�/  2�� ��$ � ��/ ��Ȍ/ �# ���c 
�����[ 轹��\ �[� ȱ[� `�c 
�����[ ����\ �[�$ ȱ[�% `H�Z� )?	@�K � I��-K �K �  ��� )@��J��K �K �" �8��" �� )0�" Ȍ  �����  � �  �K � z�h`H�Z�) )?	@�K �) I��-K �K �. �+��* )@��J��K �K �0 �8��0 ��* )0�0 Ȍ. �+����. �* �. �K � z�h`H�Z�7 )?	@�K �7 I��-K �K �< �9��8 )@��J��K �K �= �8��= ��8 )0�= Ȍ< �9����< �8 �< �K � z�h`H�Z�D )?	@�K �D I��-K �K �I �F��E )@��J��K �K �J �8��J ��E )0�J ȌI �F����I �E �I �K � z�h`� `� `H�Z�X ���%�Y ���X �^ �Y )?
��l��` �l��a �_  )�z�h`�^ �* �W `�_ �`�S ȱ`�M ȱ`�N ȱ`�T )
����P ���Q �T )0�U Ȍ_ �O �R �S � �b `H�Z�^ ���L�M �V �S I�V )��V �R �P��T )@��J��V �V �U �8��U ��T )0�U ȌR �P����R �T �R �S )�K �Y )����
�@����K �K �V �( �K �W ��* �W �O �O �N � )�z�h`H�Z�  �  2� �# ��! �/  >� �� P� �� ���� z�h`H�Z� � �
� � ��] �d )?�] �Q�� �K�] 
�����2 ���? ����3 ���@ �1 �> � � � �d )�����  )�d ���  �� ��z�h` �� � �� � �� � �� � � � �� � �� � �� � � �!�  �!� ��!� ��!� ��!� ��!� �!� ��!� ��!� ��!� � �!�     � �!� q�!� �!� ��!� �!� q�!� �!� ��!� ��!� �!� ��!� ��!� ��!� �!� ��!� ��!� ��!� ��!� ��!� ��!� ��!�     �} �!� � �!�}�!�T�!�.�!��!� ��!��!�.�!�T�!�} �!� � �!�}�!�.�!��!� ��!�     � ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� T�!� ��!� ��!�     � �
�a� �
�a� �
�a� ��a� ��a� �
�a� �
�a� ��D� �
�a� q
�a� q
�a� �
�a� �(�a� q�a� d�a� q
�a� 
�a� q�a� q�a� d
�a�     � q
�a� 
�a� �
�a� 
�a� �
�a� �
�a� �(�E� �
�D� �
�D� �
�D� �
�D� ��D� �
�D� ��D� �
�D� �
�D� �P�E� ��a� �
�a� ��a�     � �
�a� �
�a� ��a� �
�a� ��a� �
�a� �
�a� ��a� �
�a� ��a� �
�a� �
�a� �(�E� ��a� q�a� q�a� ��a� q�a� K�a� _�a� q�a�     � q�a� K�a� _�a� q�a� q�a� K�a� _�a� q�a� _�a� q�a� q�a� ��a�  �a� q�D� d�D� _
�D� q�D� d�D� _
�D� q�D� d�D�     �.�a� ��a� ��a�.�a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a� ��a�.�a�     �  �a� ��D� ��D� �
�D� ��D� ��D� �
�D� ��D� ��D� �
�D� ��a� ��a� ��a�.�a�.�a�.�a�.�a� ��D� ��D� �
�D�     � �
�a� �
�a� �
�a� ��a� ��a� �
�a� �
�a� ��a� �
�a� q
�a� q
�a� �
�a� �(�a� �
�a� �
�a� �
�a� ��a� ��a� �
�a� �
�a�     � �
�a� �
�a� q
�a� q
�a� �
�a� �(�a� �
�D� �
�D� �
�D� ��D� ��D� �
�D� �
�D� ��D� �
�D� q
�D� q
�D� �
�D� �(�D�     � ��� /2��     � ��� ��� ��� ��� ��� ��� ��� �� w�� q�� j�� d�� _�� Y�� T��     �     � _�� d�� j�� q�� w�� �� ��� ��� ��� ��� ��� ��� ��� ��� ���     �     ���  ����  �� ���  �� ���  �� ���  �� ���  �� ���  �� ���     � ��,� ��,� ��<���<�     � ��,� ��,� ��<���<�     � 	�!� !	�!� #	�!� %	�!� '	�!� %	�!� #	�!� !	�!� 	�!� �!� ��!�     � #	�!� %	�!� '	�!� *	�!� ,	�!� *	�!� '	�!� %	�!� #	�!�  5�!�     �n���A   (( '( &( %( ( ' & % (( '(      �J   �J      �   �     ( �
     ( �
    	
�
	�
	
�
�	��	
	�

		 �
	 �	

�	

�	
�
	������������������������:�  ��$�  r���n���  v���r���              h�z���F�����h�z���F���*��������	���3�Z�e�x�������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���
�