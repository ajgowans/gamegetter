                                                                             Q @i @� P&i�U @T ��e PQ  �  T                      @A@UFPX` JaPIPd�iH��� PUP�t@U  P               � ��T��R)dHAQJA�@�P)XQ�ReJ)
XD�  P �@� $  @DB���V@�TEP!Uh@EX� XU!U�RE��R Dh Z��P@%     @ �@  ` PV		P� BU% �$D � �TED�� I @( �@ A@    �    P   �   @  $@	  �  @@@      P   @PUUUUPd&P��PffP��PffP��PffP��PffP��PffP�������j  �� ����Uf����Uf����Uf����Uf����Uf����U��� �j   �  V
  Rf  V�  R�  V�  R�  V�  R�  V�  R�  V�  R�  Vi  R
  �     
   &   �   j ��P��j�V��j ��Y���� @YU `  @��                        �  %  �� XU L�V[� �j  �  �  �                               �  �
  )  
(  )  �
  �                                  �  �  j* �
� �� �
�  j*  �  �                          �  �* �Z� �����������Z�  �*  �              �
 ��� �����
� �
j @**  **  **  *j @*� �
��
������  �
                          *  �k  ��  �k  *                                              P  �k  ��  �k  P                                                 �W  �G  �W                                                        ������                                                     @  �  �  @                                          �  �	  )  
)  V&  �  �                                  `  i*  	X @� �� �� @d  �  �                      @  � @� �W��� P`P� ��U� m`  �  T           � ��/ �P�@x @@  -	  /  $.  }6  m    `� �5� PY        T @�W P?�?���� ����O�������P�@�W  T               @=_ P�������  < �?� ����P�@=_                 @=_ P���������  0 ��� �����P�@=_            @   �  5 @? ������� ����0�������@?  5  �  @                      PU @�j  �� �� ��@�j PU                                                            @   �  @Z  �P P
���P骪��                                ��  Z�  U�  ��  �� zU�nP���                      @j TP�@i�Z�j� 忖   � @��                       �  �� @�e �Z$@���j	T����  �u�	�V�@�                �  @�  � �z����       � ��� ���   �    ���� �z  �  @�   ��  A� ժ�@U����i   ��+ �� �Y� ��/ i   ���@U�ժ�A� �                     T  PZ @��P�J @��  PZ   T                                    U   �  �� P���� �  U                                �j  i��
A` 	�Q��V�xe&%��Y*������ ��               �   �  �Z  ��  (�  Z  �Z ��� ��� ���@�UUU��������   �  �i�������������z��D�����?if�_���_f�������ћU��O�z����_���w������  ��  ��  �� ff  GD ��= ��� ������9UUU55UUUfff���               Z  �� h�@���֥{��@�� � ��  Z             @�jf   �  �&  �	 �f �� �* �R�jfR�j�*  of  �  o  �   o@���           �  @�  � �z���� �T� ��U���� �z  �  @�   �                �  A� ժ�@U�����
� �Y� ���@U�ժ�A� �                    @�  � �j� ��Z���F  �]���� ��Z �j�  �  @�                    �  �j  j� �B* �� �Y�{�� �B* j� �j  �                       ��@T�@d %h@$�WP)h��+��j��
 �� ��               �_   �����IDDDdUUU���� ��� ��� ���  �Z  Z  (�  ��  �Z   �   �������Ѧ����Dt�OU�����_��w_���_���?ef�������D����z��������i����� ������UUU51UUU9fff��� ��= GD  ff �� ��  ��  ��             t  @  �  ԯ  ���� �AWeKg����  P� �jx  �   �   @  @�  T@��������j�	j��j�	u��$  � u� �� ��	 ��                   �  @�  � �z����mf �z  �  @�   �                        �  A� ժ�@U����ff�@U�ժ�A� �                 �  � �j� ��� ��j��VZ  P  �v  P���V� ��j ��� �j�  �   �    *   �
  
�  ��
 �A* �V� ]Z��SZ���� �A* ��
 
�  �
  *                � @d ��`` ��@	�T	�^}	�fI
��� �� �� @�     jU����P� P
�  �P  @Z   �   @                                    �� nP�zU��� ��  U�  Z�  ��                                             �   �  �j  `  )E   @V_ @~ ��U �ӕ �z� Ы� ��_  ��    �� ZE U h B� P� ���  �� �� T�~ �� ��+ �� �� �Z       Pj   PU T^ U\  A@A�U�QZ倥j�����@�Oj@��� ��� �o�  �j  @�   d   X �P  UT}@q*[UA)_eU!��F:���ꮺ����* Uj �                       �  J � � �R  �  h                      �  e @P��`  T0Q������^����@�n  �  P                                        �  Pf  �� @fV �YU dVU �UU fT                                �� fff ���	UUffUU��ETUeUU�ETUU                                                         .           @j P� P ip% �]	�S	 �& �% �_1 ��= �?  �  �  � YT@ V� Y� ֑* ��j ��i ��i �i Zo[ F�Z �� � ��@W�k�f��e�_UUTUU�RU�[KT�4-T�ҴP-M�@�4�T�ӤS=M�S�$*էJ�W�Ry��8uffl���uf�   �   �  �  �  �  �  �  �  �  �  �   �   n         UUTUU�RU�[KT�4-T�ҴP-M�@�4�T�ӤS=M�S�$*էJ�W�Ry��(uffl���-uf�UUTUU�RU�[KT�4-T�ҴP-M�@�4�T�ӤS=M�S�$*էJ�W�Ry��uff\����f�      i  ��  ��S`tDdpYC	��	Z� ��Q�Z����@�� ��   `�`��� IҤ MӤ��}� *�� �����j�I�D@ VU� if� ��
            M���e��Ki��F��V��Dz}*��)��)&�Z
 �
  �                  � �Q�fV��Q�fV��Q�fV��Q�fV��Q�fV��Q�fV��Q �V  �`�`��� I�� M�$��}�   �   �  ��  �` ��  �E �Q �E� �U� @Vk  �m���/e��oe�/%�e����Fi})Q�)T�)��Ze �
 �               @�@ ��  ��  ��  f�  ��  f�  ��  f�  ��  f�  ��  j�  ��  ��  @�@`�`��� IҤ M�$��}   �   0   �  �  ��  ��  m @[ @�  {D  }Q]Ի�.���oԽ,կw�� ��_d})�)G�)V�ZD�
Q��  u          �  $  h  $  h  $  h  $  h  $  h  $  h  $  h  �                  �  �) �� �� �����f���� ��  P*         ��o�7���_�畍 W�����d�d�`
�ŉ�`�������Li��抭Ŋ�d� y� 9� Q���	 �� {� '� �� �� �� r� ԗL��`���������`������(���7���U���F���d��`��������(���7���F���U���d`��7�o�"����o�7��d�d� ��)������ � &�` 	
  	
��`��)�`摥���d�`��
i����)����0e�����������
��p���q����� ��`������

���	��	�o��`)����������
������������ ��捭���LX�`������������������������������������ !�*+�45�"#�,-�67�$%�./�89�  ���������ɭ���ɭ�`�o������`������`����=���Ņ����70���7�`           ����������������`�s�t��
����������٘��ژ��������N���O�������(��7��F� �U������d��`   �� ��� ����ȘΘΘΘΘΘΘΘΘΘΘ � � �(Z�Px������������������ΘΘΘΘ���������	��2FZn�(<Pdx���� 2FZn� v v v�����������>�2�2�2�2�>�>�>�>�2�2�2��ooooooooooo����������������f�~�~�~�~�~�l�r�x�r�r�~�                ��
���������l `̚י �;�`���̚̚̚̚�����


 �ɀjɀjiF��ƋƋƋ8�
�`Ǝ��


 �ɀjɀje�ix����


 �ɀjiP��`��)��s接�



 �ɀjɀjix8�s����



 �ɀjɀjɀjiP��`�(��)��x��ƌƌ��

 �ɀjɀje��`Ǝ���)��x�ƎƎ��
e� � �ɀjiP����
 � �ɀjɀje�e��`��!�)�O���������8���`��i��`��8���`�����}󚅋��}���������}󚅋��}����` ���  ��� ��)�L ��接�


 �ɀjɀjix8厅���
 �ɀjɀji2��`����}K�����}c���` �����������  ����������� �����`��
���������l ����     ��������������������������م������`
��՛��֛�L�ۛ��      ����`�����Ɛ`����拐ƋƋ����挐ƌƌ`���n�`���!���` 4� d� �� �`��0`��0`������	�������"�
��@ vȐ���`��0`��0`������  ��ƫ�`��������	��������
�"��" vȰ`���o� �������捩
Ls�`��0`��0`��� ֜ƫ�`��������	��������
�"��@ vȐ捩
Ls�`��0`��0`������� �ƫ�`��������	��������
�"��" vȰ`���o������捩
Ls�`�_�s��ud��u�o�����v��`
  ���u�d� �� �� � ����`�����o��vɠ���ɠ�`���70Lڝ������v���(���� ��)i������`�����v ��)i�� ��)i������`����0`�v8��ɠ����v`��i�����v��������% ��)����������
��l���m����� ��`���o��`��)����������
������������ �঒��` �� Ϟ 9�L����0`����0`���v����	��������
�"��@ vȐ������`��0`����0`������  �ƫ�`��������	���v������
���  vȰ`���o� ������������ X��Ls�`��0`����0`��� S�ƫ�`��������	���v������
���  vȐ����� X��Ls�`��0`����0`������� ��ƫ�`��������	���v������
�"��  vȰ`���o����������� X��Ls�`d�d������	�o���������_�Z�
��^���_���b���c���f���g���_�V�����������������`     v�j�|�n���r� @�@H H� A}A}}}}   �ś�`�������L蠩��` Р枥���d� ����F� ΡLĠ � �� H� <�L,����������`枥���d� Р ���iɠ������� <� ,�L������������������������`����������������������` N�Lw���0`������������	�"�
��@ vȐ��`��0`������  ��ƫ�`��������	�������"�
�� vȰ`���o� �����������LX�`��0`��)�`��斥��F�`�_��`d������������ �`ٺ�|]> ��0`�_��`�� �ɀji@���� �ɀjiH����8���`��
i�� ��)i����������
��l���m����� ��`��������������������B�&�0�:�A�F�L�V�=>�?@� �� t� �� � K� ��L��`��0`���0`��������� ��
�	��
�"��@ vȐ��`��0`���0`������  �ƫ�`��������	��� ��
���
��" vȰ`���o� ��������������LX�`��0`���0`��� e�ƫ�`��������	��� ��
���
�� vȐ�������LX�`��0`���0`������� ��ƫ�`��������	��� ��
���
��  vȰ`���o�������������LX�`����o`��� ���
��� ����`��8����� � Jf���8����� � Jf���
&��
&��I�i����I�i����Ū&�)��l�` ��0`���0`��� ���
��� ᚦ���ɠ�� ��ɠ��
`�o�`��0`��
i����� ���
�� ��)������������_
��p���q����� ��`������o�`)����������
������������ �ঞ�`�<������o�M��d�d�d�d���������������d��4����
��`�ś�`��枥���d����o0����o0������������` Q� t� �� +� �� r� �� a�`$$$...8888$$$...ƥΥ �'()�123� ;<�����ޥ   �   �  ��  ��  �� � L� �� � L� �� �L��`��0`���M0`�������5��A�	��
�"��@ vȐ��`��0`���M0`������  m�ƫ�`��������	���5��A���
�� vȰ`���o� ����������M`��0`���M0`��� Ħƫ�`��������	���5��A���
��� vȐ���M`��0`���M0`������� �ƫ�`��������	���5��A���
���  vȰ`���o���������M`��0`��0�o�`������������	�D�
��� vȐ��`��0`��0�o�`������������	�D�
��� vȐ��`��0`��0�o�`������  ֧ƫ�`��������	��������
�"�� vȰ`���o� �������棩LX�`��0`��0�o�`������  5�ƫ�`��������	��������
�"�� vȰ`���o� �������椩 X�`���o�L��������� 
��¥��å��� ��`���o�L��������
��¥��å��� ��`����`��)����� ��)e��� ��)e�����������
��֥��ץ���� ����`����`��)����� ��)e��� ��)e�����������
��֥��ץ���� ����``���o�`���桥��0�d�`ơ��ɠ����`���o�`���梥�ɀ�d�`Ƣ���P����`��8��4��4`�4��8������ɖ�K��8������ɖ�=��M�o�`�����o�d��L䩠 � ������M�� i
�5�� e��A��`����d�����d��4��I�i����I�i��`���M0`�58��ɠ��5�A}[�ɠ��A`���5�o�M`��� ���i���5���A���M$�)����������
��l���m����� ��`���M)����������
������������ �ঞ�M���o�M`���M`�����P��d�d�d�d����������������`�ś�`�������LM����` Р�)?� r��)� x� ��枥���d� _� ��L��` Р枥���d�����iɠ�������L��` ���`���������� ᚥ�ɠ�����ɠ���`�������
��p���q���� ��` �� ��`��0`����0`��������������	�"�
��@ vȐ������`��0`����0`������  �ƫ�`��������	����������
�"��" vȰ`���o� ���������������LX�`���� �ɀjɀje������� �ɀjɀje�������8���`���
i����ɠ�������ɠ�������( ��)i����������
��l���m����� ��`����������`)����������
������������ �ঞ��`���������p���8��d��)���d���o�M���A��`�ś�`����0	�<���� X� ���)枥���d� ~� �� �� �`���M�o�`��i�5��i�A���M`���M0`�58��5�A}խ�A�5ɠ��Aɠ�`���o�M���5`������ ��i�����5���A���M� �%�))����������
��W���X����� ��`���M���o�M`)����������
������������ �ঞ�M`��0`���  �ɀji@���� �ɀjiB����e���`Ɵ��ɠ�`���d����P����`����` �� � T� �� 
� :�`��0`���M0`���������5��A�	�"�
���@ vȐ��``��0`���M0`������  �ƫ�`��������	���5��A��"�
��" vȰ`���o� ����������M����LX�`��0`���M0`��� n�ƫ�`��������	���5��A��"�
��� vȐ���M����LX�`��0`���M0`������� Ưƫ�`��������	���5��A��"�
��� vȰ`���o���������M����LX�`��0`��0`������������	�U�
���  vȐ��`��0`��0`������  X�ƫ�`��������	��������
�U��  vȰ`���o� �������棭���LX�`��.�)��(�()����������
��.���/���6� ��`�(�()����������
����������5� ���`��
��"�  ��  �  ��  �  ��  �  ��  �6�A�L�A�CDE�GHI�MN�CDE�GJI�PQ�CDE�GKI�ST�g�i�k�m�o�q�o�m�O�R�U���	�m���� m���� m���� m���`����M����LX�`��0`���M0`������� Ưƫ�`��������	���5��A��"�
��� vȰ`���o���������M��
�"���L�UU@ �,�����H  �]�޶�w����ݱrI?��_#'����?�q�����{�o�e�p�w��C��y�\�����!nPNlo�#�GN�A����ޗ "�-���"� ���P~B3m3�U!�X�K�������Cc=�������	�������u��ҫغ���B���u�!£�� �j���T�ymz�A�(V��R0��.��m�JVקKߐ�9�C�e5AM�F~�jh`�������+�{:џ69U��X1��6\��@#�.L`�*��{.F��Y��=0��3y=>��<e`1�3���b���b�t�$�-���sb%/$!w	a����T����#ll��������~���^2�!��/�!Jq���*5!}p5h4�=����"��+��/�Fop�]s�_0P�A��Y<����#FJ:aUf '��
bש�Ġ �C���#$#�U���� ,� ^w/1��m9Eg�Z���.[��dn"&� Y�½:S�m���	U��������pRӴ���9�4Q��ڠ����-��:��V��`����h�Ơ����la�!A>�-*���Z=������K�e*	t���n���K�j���tJa�"�VɄa2���O)2��ds�D
#u��
����o=RZ�L�=ϕXx$�C�FO��(%��C�uY d�l\�������1z�����v��2�W5��+�u�`�(a ����a���y�i튰��!�z9�	�r�e��N��S���� #��G�\I�ȀC,٥)�5u�k��h9���t�OI���v�i����0�F��L6�-�(0�8�WEs��9���a@Q�$j�Z��g�16����ր�l)���|�U@AM ��Ye߹]~� ���K�9�+�z�!PN�'�!D1�=>\\t��AQ����:�Y��­!�;(X�	��ѭ�z�Q��&�R�S렘1Ni�����Xw��;��C=�����ѿ��)_�?�B����B���b��� ����*���FC	e��Ж��� � B�K`G%Pҩ�Іp���E㚀�@)n
.)Y��3�H"�n�c�XRp�a8⦑\���+���V� ���������4�fЦ�r�)8������2� ��p$*>ą5�o�/�@�I,���Ґ�i%$� ��/ۗ �ʉP���"��i9^�����r����R?>w �S7�A ��=�/o_`
Ϗ�f�	��k> �6�uc-�Iq����PR(�)kNC�&�)��M ��>?�v `�2�t�Ѵܧ_-�{�� 0m��i��ku�C�K�;����$�i4��a 8	.Bu�r�{�칝�{�:��ݭN8���c�b��*��
��P���!C�u�p8��&����.�8Q�Q '��	$n������"i��	������H��6w��Ѱʺ��-$�y�ߠ�8p�ZDW��� E��%N�dDo�|�X�G1��.��1�Ru�]��F���H�{׮��׾�HÝ�/����Dhm�]Ye���y���"���\��^ȃ��w�3��\���by�\��#q�>O�.i��#�m��у�_\������\�:y���|Rd����EFv�U�>)44_^��*��[�jϕ�B�L�<����Z�e�$�S�󤀓Z�\;�I�H�b"��pp|Y�!�w�� i�>	.���$�v�ڲ�|����u+ć�E�]T��c�E�9Dm����;�8�x�'^vZ�W�,D(M়ו�(���N�$�ۻ���i,웭w�u*�ww6��n�'��""��$�5�P�	f�����ͿC[B5	iH�9l��WjL�>�ܭ�]@#���ؒ��В W[<�o}��X���UPjIHy_Q"��8������a*b�!�c���QD��$@�yE�=��I�$'�JI2���"6�^�1�O5� X�e����6�mmv��BCJ��یp}ϐ��׀��R�Pr��8�0x�� $��J�P�ӈ�P�l/DFx�h��H��a���,EbFQ�c�&��g.�@L�>.�M��X)�v�0�*I.��S$�${cLx�	�m������B���=�]K!u���9{{j�Tx��X���SC���H�<3��$��"�������7	������α�1�e���
��.ҋ6u}(�qfHŏ���-��/�*z��%�x���B��)�,-$+��g|�"���qP��"��#
����3p��	v�(��a�W�D/�d�k{X�fѦ�F
��U���*�FqH4�~��LӋ�T#�v�B��g�[R��0~�v�-�)L��H�+�]�.�D�S�!�0�١$x_Wu%w7N�e͎����bh�W���!�&�4	O�����л �Zє��8�F��6��e��K^I"I��rH&��	%�-Ė�J����oc���l�������fIW�D;�w)�o����n؋H��GH��l�_����?�&-�ؒ�EC�5�w�!Tl�דk��Z3���NIUB�,8��OG@�3��ķF2s��@�Sq��_I�E�ڗ�%����<�%{N����6)�^w�N�q�BI�:5y��&w�"T6�В�6�V����Z���~�%�K���},y@�@#q��f�P�p.�g�)6a4�T�8pj	R�z
4�[I�m(���N�	C���g\=���/+��6UN8��}euӱ�ʇ��|��Yg�]eE�d=7Y�������D�k�<�@��J$��|��X�-������V���[�#|��Q��b!�O��IlٻKF�y�Rq�]j\GM�Ix���5P����@y✲d����H�ⴿ��e��r�
{��tDk��0�Wt�)��Lޡ�Z5@)5���/��6�y���b^��0�3�⑫�A2kdʁ��m��4��bԺ��D��j&�MO�W�8��B/�X)Ba�Fy -8(]C�"%�l�P�7���7Bا�֒L$�Is���� A-��b�4锨�YDީ�Pm�UK�6z�lA��l�"�$t��F���9�D""	%�ˑ�B=��b����}��&`��h��q��{��v���a�8�����\B�1������$"�!~�/~�&�Վ��D߸���/�D�ǏOi�Dc�4P�,_1Љ�_<jM2o�Ň�FD�μ4��3���*��8�8��iQ��{~�H�$�ɥ#H��ؑ�H�g4���t�_�D����Q鹂y�=���'_�����/��$##D��F)&:� �}�0����N����=v���}`������B'���v@���d(��q��ш�L�u����T����"&�������t!�8�����"%�E���(�O���B"0<Y" ��\���� �YF�2$R���3�rx�����
 ��d���^B�~>�$�W p�H �~IC�$I�cc�&X�98F���b8�K�bX�xq���9r����V1̉�\N�>.$��P��H���G��"�IV%^�� P2��$����>=}X�����������w����J'�!��x�D��rt���0�,C�I:�݂ �$#	vۖQ��N�	R2]�We�gNB\p�&�$XK��);�ԡ��>ޫ��p�f��������@�?�D7���G��`�B�t��&۵΂�����`$ �C���R�_�ս�{���t i6��F�m��m�d�&e��d��p.d��%˙e��|���rq�/��.|�q������A�詒-wC.:��L؄)�p������ؽW����;l2ե>9��2��0-O��mn����J�U�]�n٬6�7�s�/CX��e-��>�����XLl��yu^-��*�m��H4�}�(G�Z�b�^j��ZG�$�[f͋	O�YV���K��3���@���_�^J��N�	Ȉ>J�p�������qC5��K�ưg��4�m���$^&]�k"�+��-J��J���Fqj}�@�.�V�J��������+����%7j��Ϳ�dV|"~������c���k�,l�C��搢��.���]���kD�h-P����n;�0�������\&����1J�_�c ����ۭjїӥJ���f%�0CX��J_I�]q�Iz� ���X��Zp?A�W�W~�26��b����?HV
4{��=fM��φf(�P�g|-�F;;;s�_ʰ����6��;e�4c"�yLS��/K��	�o�ۡ����F�����g�`��	}�0w�`���i��`�ժ�Я�5���+Jm�}��M�?�6#���X����2���]�7QM�?Km�k��av��0K�q�6�,�
2����j�:�b.e��x��@j/�%O���`�-s,_S� �i���
-��0�2�;�T�GQ}.���N�Dd�EY�A�E"<���PmЩ'�
�\�~|��T�Kb��b� m��*��(AϪ���b��yr�������-*�H���w!��1QύX����8%���QkL,���Е7pfX)�ϩ��v;rzq�򴔨V�������wa|�y� b7:�x�U��4��2�+ŏ��k�iy��Z��1j�UG)xи����.��-��kJ��6��e�?d�e/�k���T^�a�e¤�gc�(?�&�	n.i�}=%�2}�0dL��v���%~�;J\��{���yuGm��2#tl�*h�_�Q�)��D˚�tJ����2�����Ѵ�󴪏p���qρ.�U/Pjq8��Di�U����ʴ��4�W����J^�����w_�u;J��!i��\�%#͕��j x-%�P�������y�>�����Gp=|#˟�'9x��4���nz˅��@�y�M'?�>O����B�j/�i�)��u�k���gG�O�sM�T�)��Ŭx����Ŵ�a�`QA�OV)�me�,
��m9Cg��d��<��o@�q{A)ͽ��fźՃ.�@���f
9��$Q�n�f��j�`�M��`�\���n�֭_I���[y
���J��C	>����j>��f�<41���m4�@}�L;h
�_q���;��s���"/x����yM<��J�kѽ����V�XF�7urNA_5n�^+��(�8�f!B�z�6�.�����S�&y����R���IJ���Ź�jt�_����S����:p��m-�a0����k������S=����Jb]w�+bE_��y�F��E��ځy$v]��?k��ЪF�0�5�9���M;m���U쑽w	|�0Lk��gA�����x��w���E|��7�6V-b��	���v���|�O����x�ݐ{�仴Eu��p%_��QV'(�8�W\��:9���y����������b�dt�8`�5�.^VO��ZO�M�^�X�?�7�L�t@,��d�] C|�|v�*}P�È�|脱�/Pٳ6�"�}�b��)3x `�e���O*2.�爾_��ejn<���"k�k���zs�^J��(�W)y~J�s>��/^��-�H>1~"��o���%��������Pe�^8�1Qd!��8���iς �)82��^��Ł��;��ίD��<�0����^.39~�9!�HxUH�u���b���~��!��/δF#�����*D
��^�~���焽�0ߐ:������j���0[4���'��$��԰
�F7�0�<Ԟ~;jVP궒��"����5I��%�e�S�W�A�X� ��䮋�K�r�j�P��c�V v}`��1�v�ķ�p�_����J��x�_��y�����b�_�!P�����? ����,��_�T\y��iw1}b]s�^;�~���^S�f/y��^��ݡ�wY�/�l�䲹w����y��'��/��^�b��g��#����/6?"���Э��s�_{�/�t��,�{bR���-e������\3�}`�y̖3����%ʘ��������~%ꔽ�ï1}���@5=`����<��7�W�;^��+X,��޳���Goj��L�.�!�C�1�CP��um�AfIً-�ݏ�����y��.��HKp7y��,��N$������x^R�k���O�[3�/7�/a9O'�Ea��
Z!�I:N!8j��^O?���	y�;=>�|&������C}
?���3����Z���^� `�:Z�}�y�"i��Hp4�Y��t�5�^��,�F~@18�B�G�/�WΒ�1��j�C�J�QC��n.�5� ��W6���%�H������� X /�|S�	��㤿J�߈>w� n`����l9�/�.�w��3i���BKl,5̹A�/F����|���7�I`-�Ǆa0�	��Qt|E��_�η:�ר�%�g���Sx�Y���aa����5'��B֭��1x��B�[��������ry�u8���:�Ҫ��E����2z0�pAZ�N���Ix�Q�z?[��/=X��_��ۑ�id�"�.z���Ʊ��ļ�Ã���=�ĺA�7ĺH�B<�|r?������;�`E�t��4ۺρ�E�f �K�\�E��V���8�}������p �B8�u�$m�7m̙rx%�m�[���ܾ[��2e|��T�_��Y�&�1I��& 8u�e� �ύ]�'Q�/�1(D����7�pjݻ��F���8z�Ȏ8�W�8NȜ�^|?��ձ8*�j��6c6\���6ڧ:�E�]ֲ8A�$sB˄qh��U�G�8�ͭu����A."j^�p�iH_˯��r6R�� �ŋ$s^�g���l�OmBu��N+�
�F�@����*r���F�uZ�Q]��ݍ\<'>@��sW`*��f��v�ΤE�	�V�k�����sg"�y=b�t���z��Ө8 8�\��\u��X*�MZ�����?d�%�V#z�.NqSWU����I�q��\�7ɰ7���MMM=O9��#q��8C�p�F֨+�B6�==+>U�t�p[_��O�〨ɗ_�q�ih�h���n�?]wNO��l�#�����P���>`H<8N���pVݠ��T�cȚ��c����k�:�|Ff`��As9�+�U�9η)��:��ǡq�R�p0�V;k�K�̎9�wR��W=c��p��=�g),�ŗ�rM�.w�%��w��U�6�s9�ۜ���� ��*�w��s��Ӌ|G)����,k�U#q��)�d[�9K`���q�W!���@a�↸-����f'�qW%�F���p����f*�[����i����f΋kCF�ݔ�8y�|*[kx`��\l�8��q2��P8�"������>y�|�����(��~:��^�����:Z_�p*Sf1	Y��>q�x�. q�|oi:�A��6j���1��'���	ő����-/ApSU��h#����Z�pҳ7���n�t�ȉ#��+��!\gV��o0��f���%��'�.m]Z�W7���@p��'1��Y�C/�q���ߓ-��?�g���H��N|��c��s��pfom*$�W��4	� z�[V��	ƙ����	���ŉ�9��5��*a��Ȼ�߲�ͱ�r�<ƺ�99Qߞ\��"���]��БÝL���M�������S8֠���q��u=WMn�SS�.��D�7oV�Rz��9����7��Fg�%Ƴf�=��׋��|q��v��Bzn9����
�_��LLA�w�F_)�p���Sy�����Qjlr_ [Q:���x�a��"�c=��bx��o>���C��Õ��,O}�˧F,� w,؄q�oޣG���)���V�'����XŬv�g����Ue��rBG>��&+or��p��-U�}�32� E������K#M����y�.��Zq��·�s3Nn�n��0�(_,f9({�,�x�D���R��fj�����Ykr=�R{B�0��[��W�m�[]K6o�E��̥PAŷ��4ۏ^mE�Y��(��@��=�ښY��f9@˃�m�&��g��]Ds�t���AA��dyNdX�I�h"Ip�I��<�|����ݐ߿�|6޻z�of:��=c(��kG�o7�o�,��G9��{۹��	����Ѝ_��}'��"�q�g��Թ�+��*��f���MD�;�U�v���k��λ�3��kx��5����<��]�r߽l��Q�C�X(��t g�(W��A`0����(E��ģp�'oX������:I�נජ�OzPT�66�$5?�b�01����|�fnD�����	�QJ:��L�v��D<x%14tC�p{3-׷y�n�M*RL8��/�:�f�nFlJ)�G}� zG��ʡ&��
�	%�%y&�Jg\�9�����gi0�d �� �Z��1�	�9Q��o���&a��-Pέ�]��s/�e���Rs�9z�7��E��p],��=Kzn,�а�x	��6ަ���ht��R�}?%��է�P�=�6� �&Q���S���
nn����i]�{;j�==A�Jc5ŝ	��۪؝)�א�B����kS�+g��8%]��v��HrfF��ʇ��8%��&�x@�[�F�s�E���9��9��!�r�Q�R�x,ܶ^����s�KW!;��e� �2hͮ��j�����\���P�sH#�TK��B�\i�T ��w�ԫ����p	pYO�7��~��g��ny�� |����J>	��ޙ�Wr_����z:���/r怗˫.��@z:���U�}u��hO�E��������
���ܚ��믧�����r���ϡ�*_��d��*�B������3�
& W`)�x���^������ȸJ�L���	�ӆ�A�3�>�X`}�c��<�N��G o�]�c>c)�����KN#8"c^gO_�]bt�pL��#��9�q�r3��'Dq��;�A��	�bt��ŕ��9 ��}����+�sQe��8���\�$��E �/���m���fY.%���f��ƭ��Cmx#� �z2C���pU�pQD�8�I�pn��9�$����^��'��ݬ8��.��������Y" '�v= c����Ar��z	�7Ë��:� ���w*��{XG��O��)ڄ�8\ v�R�m�ɹ��!�8W�R.)�*^��|#�0Q@��K(b-�~���)XT5��x��8V�?r
��� a��iI�2��Y<Do�gJ:��^�v�>�N�`�G��r�R4ٌ�~R7�;M;F�	/��=u�8�	�RM9���ۗA5ڒLJu�	�f���a�[v;7+g�a�:���k)	k6te�7&*;N 9�Nq��.^�nmK�I����8>O �m��I�7<��bm��7����*��+	;�v_�u�����7ƅ�š��ĤߛA�G��m����N7q��/�8р�p���7D*_�īXG�����&(�5��Q��7i��n�9k~&�M�3�B�`�<8t����N�6�ws����� B��>�ů�щ���{���  !�[�ۛ�6�d�[�ݗ�.^�s&����Źd��_;��'s�O���I�!�R�㋓��*zӡ�l�b�vC�L�o<��V��˖H�r�z�O�3�Hzԥ�[`� ����Y����J붙��`%�Ĳ�j����j��WY��c ���}J��?��6�J�+��u3~u��`.
�a����x�����=L%v�6����S�e�!���:��]l����� f�A0�/"��T���sg��V�S ��f�Zf�p�L]K|�{{t=�7��aט�;�`wOR��t�7C76�6�������������jg���o���ԥ/��lsiޕvf��k��E����Ͻ�Y�������Yv�����c�#7�Km��.\��]�E\j�����T�SN�.��~��&�眻f�|�}�<��ͷb^�r�~�h�,������.�s�Yw\��pX���,,�\R�]�f��N)Ю�cHLY�O�S��Qy+��������e΁8��A��O�4V�=5T8ҫ9n��NC� ̳.֯���S6��m��m�mm����~Դ�h/y�a�\������f��X
��5���Ţ��Ld���-��2���d�p�㴹��JQ����XO�b�T������7��F��ZK���z}9}���]��:����Ws�x_������}�hu,�3q�:�.o1{�2Aa�WtaW;K��kIFI��ܜ�� ���������2�uM��]G6%{�-/ouA�2�d!��\�S�Ʈ�خ����K�1	P��
��T�S��Ƥ��^�y0Z��^u�n��\߼�&��t��^�gZc����E��t���L��u�W��d��v6��P�3�Av�1�?f�{zԶ��k�����*75\l�K�'Ր��]*���k����\5����|������*�MoC-�hpz;*G�2ya?Z^ũҖ�N[�:ͽ��V�;*�4��|cXsma~��[��k|n�)����4�%��l��Zy�?�?Z��]&�nO�?Z�u~���]���]���թY�wz�7���HT�mY�o8��Q���3A��-wyl
IqW�W�l��㩫��\���55۾�㋵���ɫSTp`������\�Я]2�>��6��\=:�(.������V�"R��4�Az�D<\^|�|,00�����[��^w�����Te��0Oc�/��r@�w��s�z��qρt6��àIB��̼hS�����\�v58V"��h�ңȼu;I|��_��]0ß�������B�&/+����N�J�+�+��N\
��x����+c�S�K�Vj{��Xd3�i�)+���*��K�N�olk��r��v��	��(dk��1���/b�C��^����؇������\��a���i�U��b�.z��M�K��A�����b0nUC8\5����y��A�Kڽ|�եW�ҭT!������\��	�0��w	t�/FZã�U���(�%��	ze1E|��T�5	��lXg�Q��S�ͽ���8]�E��������Ռ��ٞ��SvW8Prp%�����_`��1k^�?TŅX_c��~�#�-�/}��Zc`A��)�h��*�?_d�U>�����KC�:Z���.��b�;��.�s;�Iaѣ��%ȝph�G�+��Ǆ�t��s���H�NŨwV��j&�}�����F����\E��/5ƹ�Ү�������*�,��F��"��tj.)xE$�K�]`1.o��2�I(=0�ie�-�M۪|��hWC0��������ǆ�BwR�Y([���.V"�j�a��\�
��s�UN��.]�q��0C�2��@/U���e�/[j^mOQ��2���H�z<@5��+�9z��e��Oa��ӎ"��nd/��h�<
^��]�ʵ�,��^��/饲%�:��ĩܜ�8޹j�L���8�򇬋�+N�\Q���e�6R],1��;ˆ�=R4w���g��������.��Y���kU���ޯ���-E�0P����(�����_yu*��4׆��,����o18^���ix��S1�ru�����x|$��z�p��<�n���޽M�J�7�K��O���)mux���\�qq6޵r��K@��늂�'͗!S{��rWe.&-�b_��t��okyS��̦�>Cw����^#��+��'�s���H�S�_	ͩ˹��W�qb[ ��;uϒ�%���8�B��_ظ]�e�I���.'��\	����{���tJo��e�vH�2���c.�.*�"�+�������Ќ9��2+�`���*�䋛�"����P%�?'�D'n��G�0*R��A���z�Iȹ��C�K��Y/(��W�E㗇|2<��=��$c���a3L%���5S!�# mjE��[�Ⱥ]M����;����|}'*�>���2�I����,_5UG�L֮��W�8�\1�_�:�q�sN���&59��S��.2��.=&1�s���n�f㨾�'1^fl�`-��zl���CxJ�Pש�����\UX�Jd���v�J_z]��]91�w��w��ٖ)?yqg��Ńz�%�_�.Ԅ�*���<�������~NH��Y��y���˹?�tk�_�q���F�IG�េt�J?�.�'����˿�w�"�W��i�~E�o�`�=�l��$ݾt�s�r����i�|���n����{��Uh21U�1de���H�.^�̷2�^�L�j�%cl���������.q�m�����?�3D�R����R�J��3vT�r帟���\��<����h�2cM4��f&����zM_�!�MM���V��љ��4I��N�4��<L���h��f�љ�h��5�01_ɣ���;��CRfRk=�h�%"���4�#�f��q��Qr������w��L������Y�C��n�@a ������	e����Z��1׺�A������*��Z�:�*T�0G�O��hB*��]tL�:o�N��r���y���Q#AY@�2�?��W�7A�2�	�sRFu*~�������1.^�݉$��>�	�cB���F^�@0	D��;��[:���������UέT}�J]	 �l�qPAPL�I�Ν�`�2D3�`����+-Z5�1t�����e� 2�Y��\9G8]��f�f%(��!���f'B���}**���8u�pII�"Y�}�ip�y`!Q0IFhle��Hψ<:��U���M��ݝ/	��M�,.����-�U��*]k`�w�?�U�!������-��ŝxȹn��,d��D�8�=Z[7�Z��g��|������À��,��<��e��[���2������oi}y7:�qgl�f���1���c�Վ��5{K�zL�eՔlHt���'�Jת��!�Y�0���@�-w�iU�f���(��nr�?t���3ASQ�2H�,�CT͓̣�ݣ�%�����!�+%����r�8�V���}�.�f��L*��&򃓧o٠Q��i����6HFd��7�ݟ3!�d��y�z�4�&���Vds/ۼ�T�Vl�zy�Ր����o��|����Y�,}�c9��^3'�~������3����g�?���M�)GoQ6a�e���qکC�Ox*cR�4�w�照ff&�eE�@i���H�
FW�E��F�$'~����2��t��\b�\n�A�DkQ��ZEI��uc�뉙�=W�她�|;�1��0��u�#���>6��cȳ��f��o��Ĭ��:LփX xL�+��U�ieV���b8M�OI���G�������d��U=��b�{����>��g^����ͭs0�e�L!R^<ҫ��9R0�(�SX��/ޕH^5����жq(���,i9l<�+��{$(��\&վ��l��{�멜���.�U�<��6	�	�{Φ�0�{L���Fv"���ۥ/X��Y�Wh�hθ�X������f�g{�}��3Y��{���k����c=Fcc�go�fi��3 �}���l��`���_��7P�l��k̳Gna-��;e��w��[mg����j;���7��|�˫L���F[q�����~LBc^������2��x��ψLu�ٜ& g�sc�'�b�:��2�3�8�3��maA��{�~(�@�݅����fU�w�f��2�Qı1��dYg�ɕ�x���6	X�8�������er��O�>���T�12�²�̢��(���TDԂ�C6Y,��ȠU��1����2�Y9��$�*���~��^��~E�T��z9��	��_mٵj׌�?OE��b��}��#,�Y�d&b���0�nc'|ل�Vh|f@����3�v��+,>E��C��Ru��x��,�un��S��v
�0堎�Qɗ��
u��2}o���a2�c5�fް0*�&s������`�Al۲4����~����;�ٳf�aݝ7��g����
��%PBBU)!Z��`
�\�����Un_��P��[���v2I&�:]>���㇓�t�A�ryӧ8s�:vC���x�Ou��C��������СC&�K���l�y!}��8����.rO�w�i�]Q�;q�̝���t�W;,�2����Fu�ɕ�B=�. ��|��}��I�l�}�$D�=9��v�Sc,�3ǟ3�P�,�l��ٻ5�=�#���?��G���#�!���O2�z�a����1O��JS_���'��� %� �	�4�����y�ժ����h �j8�ܻ��Чc����7�^=P�����1�9�_�������v�B
��4�1��]�'k��g}C�N��(�:M�)�M��,ԭ/B���sb>V�4�»>�sbŃ���R����1�+����M�N 6�V�������E����Fd�'*�6D�3'���Ce�9�f��M� ��_�m��@�\-���S6��/g�f�^�səǅ�js���-��󧕔ofh��@�>����g���'H*����nA�h��i}Kq;�M�f��X��i��3���<�.wm��I����6[d̺�f���I������4�dZr��[wB�2'�8B�f�K���sr7��g8e�P����8���`e��-w���)��s�[M�� ㋛6pS�)T8't���3\�sK᧏:�k7b�}�,�V[a�!<<�Z�E�R�t�j�7Y�d;�M*Sv����6F�Q��<	��Z�������7���ó�`f��xA�yy�b��3��q�	L�̴�^��z����\��rr淽��q���.L�9rgl�t���8�ꌖ@�-��\lF�}_�)i�3�o[��g ��$���E#��\��.�{�R���\֢K��7Y����J^~&gO���hZ)��?+����[V�M*r�.'9Y�HqAA��/��&6���w�pA��;�L�Է=����C�sz�F�����i�L������Ǻ�B�!��u�8��g:-Z���Հ�0�r/�M�U[�����E:̢�5j�w5�`�p}�����Ǘ�ɻ���<\����(��N��������i��߃��>���ڣɓ��`�'u��Q�A���r���t9P�,��;���ϖD)�n3��|C�r�y��C��r�7npi.�?��-���K��-n�SK@|`��D���x��u%߇�sP�ѡ����C��O��[�� �5:��(8�W��q*e3�Bu�ZC��
��c�{>W��'�>�c�mUÍ�c@�c�n�o;��9���]Z�����{�Gk�;O���+)����5�2(\ZJ7J.��ޚ!r0�C�G��2/K�m9��s`z�09�N3.�.���cKg����|@�e�V�k��꽼�2�V�<
#�M�K�s��9V�����w�]�P��<���ms�ed���szy���r���J����}��7c��<��3���"'��3��1�����Z��Af��r�w6F�Hg�
�_��t�TػHc�h(s�Aƒ��V�䆨]�+,��㪅v��%}��5�k�l-��N�9hKk��p��uC��5��N�9��<�19�J�o������Ǉ[�m��,��A`;��c;ʚ���4/W���q,\��M�n��:��\��Y�Ɗ�suėm�Ù�������gCB�\ 罭�eaylB�)15���Z�f���,Ui���-l�o�ą�իi��Ij���ۙ� r���U\�O���/�c��\��'y�U�q��wQ�N��&�e�[,��7�|m�pT���������8�a�(a_���V����߱	޹��c;z���`�;l��4���Z�d�$�wM�7�M�vt��?���QD 	 - ����mq~;r��h+����v2I&���:��*�ho����Ӿ�h�O�9�cy��T�ܠ��h�v�/��AT��(ҥK(��("N%�5�X-��*D�yXG�aߜJ�e���U\*h�������}��T�k��{���%�B�/��c%�ܵ]����U���B&��Xm�(r�j�,5�ӌJ	QM�>�7j_ELz[�}r�y����R���U�!������}	���έѺ�����Y��������s*5��9�u��X-�^.E�AԚ�4�T�o��Vo�`�w�UN8�k� �)CU��x�PwOJ
�s��hî�����5�Q�I�b#w(�U*ժ�i�Q��
�ڬ�&ӝ�Đ�0��+�Uv,��[�X̩�P�V�z��ʡ6�U �W������+I�@DV��U�@�J�WN�0��^yCHMR{6l��I�O����i����Q�^]7͏J6h_�GCe:{�.jC<��ḋ�[�Q��9�UvEhtt ?���C_��c�S����#o�ȭ�C]���U�)�!��҂���#��:�@o%��M�Koԇ������U�N���[B�����yY9ѹ��f�x��5�N�
B^([��㚩I�{�%U�U��<\'�M���Q#�7(Oq�s��+���{~H�(P��t���n,p8�9x�‰2��U�?�È[�LPK�T�J��
���uF5�{�D�n�J��	u�W2w�w�O窶�T��?n��h�D�k�0q=�ZR���@G���Sv��l*.Y�9T��õ��>c:�Ԁ��m�"k�I���R`���z��D&�9�<|���o�G����3��j�y�C~e���^�w��&b�!���c��
����_`R
���ׂD�?ַ�5Gy��IC�@	)ms�j��*��$>�i�l+l��՘7;���CUft+%C�0�����H�Yt���5���p�U���=���~��]0���3��U���	�����j��Aǐ�6>���$p��Ta�Pw�d9\+V���,Q�27Տ!x��v�,S8f�q�nb��;T���W�81���yA&Vtq�(��:qR�V���|��ЁL?A5N�3�6j@K?�;S��M@�Q(w褕:+�TK���(�*G�S��n�je�gR����_%gY]t�qm��0u��TՆϡ��=v�ژ��\���W�e��%���+�Vz��r��&�y����۟�Wv�=*������=��)z���%~�ycIw������ex�7{��l�W"�_���aR��W_aX,��/Ԯ�ņ�d0��Vm�e�Wa�OJ�m�ݬ����Ec�CL)J���*�^��]��K��q̭~ee�m�Y*���	C�A�X,���$�V}�W�"B�"��܊�zX���
��k|J�ŁX�m+�Y�����AX��5�E�V�l9fe����V��&���`�Yv��®Ԫ��Ʃ�;Z�{գ���\4�;V�jخR�7�C!��L;*�z����D֒���}�ɂ$�T��Y,���8�t&�*�m��Z�+�Xg��.#T�_ή���m�I1�a��d�ϐQ��ݤ!�����*�
���aq̫r��]���}�-�)��YR���@ܤ&]2�}�jh�V	E_yS><��|���wT�6��+�M�r�a���ю)��oQU��j����ڮ��v5֨�QSeB���ݸnhP"�,m�z�I	IJk�C�s�\�񢭿4��ڔ%%˜:�4�
K���s]b��P��e:�X-��U*��B�XQ�e)vY���c3�4�$$.u��^�@HwU���+�%qg{w$ ��T�.(���L�)U�">���'��1V�������n� `�(VmѤ��3�P��BBq�N��OK����tUA(�#o�U}����W(�;:������>��G��Ϗ����<�:O�@��Tqʬ2�5���V�VYf���H16��K,�Y��b�*�]��B�BO� !��!BM�אt	p��l*H�8AqR�Sf�xB�7q�B(�^��\�RXf�!�B9a�>��u�y6���%��~���ۃh��90�3��8B* ���@�#���n`�Xa�P��R,@�t� ��q�6@@Sb%$����q��!��W��4F��G�~���sT�DH��qB�o���% � ����Q��a�4B����^ŋ�C�˄.��0�'+��n��DA]�n�� ��G�%�&�H��^�v�
 N��CP�xO��/:^B�0}f����C����͂��B��qt֪"�Ddu�����,��A�5�܅R֚�N?:�̻k�_�=�(C��&����N�q`����!~��gL%W��Q^lk���di���$�h;��=]����f>�R��Gd �k�0ia{`y��V5��V�Pt+?PSI��P_Q.�j���ȑ�sa�P��u�s`t/H�u�N�B��!�MV��_[h���YӨ번���M%]�A7FX��i|��Ы��`v����CA�鉆�!z��8@��ݖ&�&+��<��
���Kw�e�@@�妑7\4�����H�]2��F�*8�De�Pߌ"��e�r��"���"+V~�C� <(a��%sW}���!������xm��ͬ`BM�[O@��& n~$���=��gp�ݍjխbK]�ɠBw?Yv��
���3���N��DįM���y�o�G��nN!ݡ��)�?Ό��fʩ��4�,���*k���ͮ�V�}��^�`�L���HP�� �q �x/U�a�0A6����7y�!��BC�X��������������E��}D�j?��x�	��D�)�+����L	ū�5�#߁��'S�<eiO�"k�?#���e��O�@�mߘ���4�Fm��	Cx�g:a��Dq���
���}g�bB^�"�A�){�h�eH��8h[G�T��_���,�E�A��v�B��T�l"�*�|i�F��!!�A��)���p�S}�I$����:��y�R"8㢛Bժ�>�#>n�l7�D4Xz%�����:&0�"R�5"P���31a]5��7�_'�	J@�Ɠ2��j0�	�1��5W3|�T:qoUG�TcQ�="&�+Ī3�< �F��`{�6$�Tc�F���^��>�4cO�x�4�%~��=ψ�����M�A�~�̖�.���*l��sp�n[���T�o�!@���y?�hp�u�|WI6"�x���<���m!�#�:�Pkׯ�G�/�8Hs��F0����-}|�D��~OP�b79�u�8?�!,��P�r�`(�c��(�]>��"*�P �
+|;����m]4ӺM�g�-�l��oǶ�`=V��=�&��ay54�!�N���T�~�=�O�-��!֎���bG,�,����!?�,�rY4����z)�����ydA�@Ă>�z*�#=�\c�6�����xÝ+$"%N��q���kp�bo��I���Xv�d�g>y��J�E耸�rXO,�0��Ujǐ�"|�3��~zI �
��/#-.K�v�d�a;�������Y&�yasνnx&�fk�tY�0�utŁ
�\����_������������������` t��  )�� 낭  )��� �� ׄ�  )���`PUSH START BUTTON  (C) 1992   Thin Chen Enterprise � ��	����� �����d�d����������y �w ���z �x d���  x���"� �#�����A���� Sũ����T���� Sũ ����_���� SŜ��N���F������������� ܁����d���� x����������LX����� �����)�� ��	����� �� ��H�e�� e������h����斥���`�  )�Љ`���)� �� ���ι��`������� 
��݂��ނ�� � ��`������� 
��݂��ނ��
� ��`����q�������d���� x���)�R����A�����A��(����JJ�	� JJ�
 |୶i� Q������


 Q������(�����`_�t�������                �   	
  �    !"  �   #$%&'()*+,-./01  �     23456789:;<    �     =>?@ABCDEFG    �߂�	
�� ��	����� �� ��.���� zũ.�y �w ���z �x d�d�� �"��#���t�����t�	 �ɩ����������	 �ɩ��t������	 �ɩ���t�������	 �ɩ��q�����q�	 �ɩ����������	 �ɩ��q������	 �ɩ���q�������	 �ɩd�������������� )���)�(����!ζ����"�� 
��~������ � �୷)� ������ a� �����斥��	��H�e�� e������h��  )�Ў� ��	������H�e�� e������h� ��`u�w�y�{�������	�
����  I���� ��	����� �d�d������������� zŢ ��0����Lo�_)�_`��斥���` H� K��H�e�� e������h��  )��Lׄ`���Lo� 5� H� K��H��e�� e������h�`�������`�_�����������_)�_��"� �# $�� �"��# �� ���  )@�`�  )@���_��0�_�_`(0YS!B1PSTAGE : �_��0`������� �ʭ������ �ʩ��������� Sũ��� ;��_ |�`�������0���������� �ƭ�`����������� ��ƯƯ�`�3����ddL��               � � �  !"#$%&� ,-./012345&� ;<=>?@ABCD&� J%KLMNOPQ&� WXYZ[\]^&� defghijklm&� stuvwxyz&� ��������&� �������� ���������������               �3�5�7�9�;�=�?�A�C�E�G�I�3�5�7�9������������������������� ��)i� ��)�8�i� ��)
�������L��
��U���V���� ����������L��ZH ;�h ��z�L��`�3��������`���� ������`��������`������������ ;���� ����`�������V�����V����x���JJ�	�JJ�
 |�ƫ�`  In the enormous�galaxy,there are�many stars facing�the crisis of�overpopulation.�for example,the�Alexander Empire�is typical nation.�To resolve this�problem,Alexander�is launching 4�fleets and looking�for the heaven in�the legend-�'the Earth'. �(��i��8������,��i��i��8�����������`��)��
i������iɠ�	��� ���2������������)����������������
��m���n����� ��`� ��	����� ���"� �#����d�d��N����d���  � ������ �攊H�e�� e������h����2��`�
��������	 �ɩ
��d�����d�	 �ɩ
����
��d�	 �ɩ��������d�	 �ɩ��.�����.�	 �ɩ��0�����0�	 �ɩ��	������ Sŭ��$ ���% ���& ���'  �ȩ��� ;��/ �.  v��	��� ;��- �,  v��`Your score: plan number: � �"��#�����a���� Sŭ��$ ���% ���& ���'  �ȩ��
� ;��/ �.  v��
��
� ;��- �,  v�`***************** total score :**--------------**              ***************** � �"��#�����&���� Sŭ��$ ���% ���& ���'  �ȩ��� ;��/ �.  v��
��� ;��- �,  v����� ;��� |�`***************** total score :**--------------**              **--------------** plan number  **--------------**              ***************** ����`�������d��� � ��`
�����L�����   	
    �       �� �S���T����m�����m���� m���� m���`U�    `�_
�����������m�����m���� m���� m���`���������'N u0                   	
      !"     #$%&'()*+,-./01       23456789:;<         =>?@ABCDEFG                                                                                                                                                                                                                                                                                                                ������������    ������������    ����������     ���?��    ����������������������������_�U�\TTTTUUUUUTUTUTUTUTUTU�U�@���5�?�?�?���������������������?�?�?�����?�?�?�?�?�?�?�?���������W��WUWUTUTUPUPUPUPUPUQUQUQUQUQUUUUUUUUUUU ��EUE�E����������������������   ? � ����������W�UPUPUPUOUGUEUEUEUEUEUE�UUUUU����������������������?�?�?�?�?�?�?����������������������������W�U_QUQ��_UUUUUUUUUUUUUPUPUPUPUPUP�P���QUQ�Q�������������������  ������������������������������   ? � ���PUPUPUP�@�@� }  E�������C�=    ���� � � @  �����?���   ��������_�] �S�Q_QUQUAUT   UAUAUU U     UUUUTTP   UUU������� �  ����?��    ����������@   ������       �������� � � �  ����� � @  ���  ?       TUUUUUUT�?��  AQQPPU���_   UPUPUTUT����  U UUAA�?�  @TUTUUPUP����  PUTUTUQUU�W�  TUUU U �U�   AAUAUAU����  @PPQEUE����  PUUUUUP ?��           U�������UUWU\��?�_�_�_�WUU_�p�������}UUUU_��< ��_�_��U5U5U� �������WUWU|��?W�U�U�}}�U�U � <U�U�U�}��U�U W ����U_}����5 ���_�_�W\u\�p���������UUUU_��?   	 	                                                                                              `   �   @                                                                 d   �  �  @  @j � �`                             �  �g @v��t tt �Ԃ�W�*�޷j                                       @   �   d     @ �	 �                  @  �   $   	                                                    P   �  ��  �  �@ ) @P  %                �� ��� ��V Tj}T}Z��Z��]>V�w�} ���pG��-}  �  �            e��YA�jA �j �ZPW���F����?�k���Z� h)
~�
���            & i �@j �� }iY �u��_�u���ݯUo� }�@�x@��  }                                     j   �   j  �  h   �   X                                                                                                    `   �   @                                                                 d   �  �  @  @j � �`                             �  �g @v��t tt �Ԃ�W�*�޷j                                       @   �   d     @ �	 �                  @  �   $   	                                                    P   �  ��  �  �@ ) @P  %                �� ��� ��V Tj}T}Z��Z��]>V�w�} ���pG��-}  �  �            e��YA�jA �j �ZPW���F����?�k���Z� h)
~�
���            & i �@j �� }iY �u��_�u���ݯUo� }�@�x@��  }                                     j   �   j  �  h   �   X                                                                                                                                                                            ����������������                ��U �E�T�	 �@�PgTԇ�U&U�.           u	TdP�% �                                                                                                      �   �  ��  �  �                                           8   �  �   ��  �   �  8                                       .   �� 0>  ����
 0>   ��  .                  ��  {'   �  �*
�����ej��j
	 ��Z ����j	�e������ �*
  �  w' ��                 
           U  �)          
                                      @   P   T   U  PE  T�  d @Y� @Je ��e ��Z hj�  @U  UU VUQPeU�Z�Z  jT�U D
@Pjh��P�U�yP�IjRD�TR�Z�E�U  DY  PB  UU E% XU ��`A���D���ET��A�� @�� -�C|�A�                           U   P    E  e  � � Z� i@
  �k� ꪪ@���������oV��o��U��������Z��{���f��k&��k��k����UzV�jJU@R*�U����EZ���V�f���V����~���J������d��!��!A��	���@A���*Va�&U�V�Y�VEY�ZQ��jf�fVzfneA��%�odA�E A�U�Y T��`AB �B fA*�" �	�	zRP*@
(�B

zN)$�Ad�q�v a��UR�w�*��������	��gY��U��P�^*Q��*F��IE��f������j �i  Ze  iU  TU ���@�~ �eQ VU PUAE �� �'Q�m� �ZV��� ��Q @B@�V $A P(� @E�jn XY!@TQ@� ���AQ ` `  � @D@P�F @��W]�Z���Z���f*��`֯��o$U�k�+%Q�)e�*�D�
E@v
Z���Q�P� �eU �VP @Z�  ��  T�  E  Pd  @�   �   P                        � j��j Q�jEFiE�R�V ��VZUU EP PPD U PU  TU   PA�Q @�     @ Q@Y �V@�U@iUYAQDPTUUTUUUU UU JD�EDY @%e � �� �� eU UU  Q  E  U                                          	
    !"#$%&'()*+ ,-./012345&6789: ;<=>?@ABCD&EFGHI J%KLMNOPQ&RSTUV WXYZ[\]^&_`abc defghijklm&nopqr stuvwxyz&{|}~ ��������&����� ������� ���� �������������������               �����       � ���  & ���  ���� ���  �������������� ���                                      ��G0QLDQGD�We��UUUUUU���������UUUUUU������  ��DDEDjf��jf  ��DUQUTU������  ��UUUUUU�Z���j�� � E1E4�Y�           ��V`�        �*D�Q��          
 � UW�WeW�W�W�W*W*W*)����������������������������?������������������������������������?�����Q�D�����������������������~���������������������������������������������������������?h�����?�?������f�iժժժըըը�     � � ` ` ` HH���ʥ~��)��7��f�?�?���������Z*1�ԯֿZZ�j�k            W*W*W*W*W*W*W*W*���������������V���_������������������VD_WT[U�����x������E���f�������������������������������������������?�����������������ըըըըըըը�  H  H  H ` `�������������)���G���o�����������g�g��k�jZ        ������������������?�������׿���f��o�����������W���������o���!���Q(��Z�f�������������������������������������������������O� �?����������D������������������ ` � �          ���~���H�`��V ���?�?�����QDĿZ�֨�*1ZU�                 ���������������������������������I������������������������������������������������������������?PG(����FH&	bf�h���� Jb�p�=��������h�h���������������������       P          UU    �����?    UU    ���      UU   @�p      	 
 
 
 
 �������������������������_��Ee��������Q�}�\������������������������������������X�����.z��m��S�m��Z��å���������{�n�{���        �<���<�����TU�������������UU�����s�|<?�UU����
 
 
 
 
 
 
 
 ������������������U���U_AhYR�V��)|U��c���g�YF֖��}]Q��T�e�g�k�Y��Թ�������_������o���{��U�����������������������           @    P �   Tj@�T�            @P    �``e�a�`�           
 * �����������������_��j�_A_�U�~(]����j���|�X�g�k\Y��V���j�Z�G�Vցݡ�e�i�Z��������������������������������������������������?����������?XCi������������������  ��X XU��  �k���]�U�����T�
****

P`��}<�<�����_P�* � � � � � * * ��������������������G��_�����
z_����V��U�W�_e�B����gi�����TC���~��U������������_���1�$_���Uig��G�i���WZ��������]���������  @     < � � ǐ����
  ��||@              �����*  <0�����0
          ��������������W��������������U��������������������������������������?�O�������[�T}yk~��e�WYK�Yj�j��Z��L�_������������������ <                       @@ P          �
�A�<0           �\           �!*W*W*W*W�W�W�WiW���������������)��X������������������������������U����������������������?�?����?h�ըըժժ�j�Y�V�D%�CUCUC@@j@UQ�QmQ�Q�Q�Q�Q�Q�** � � ���T� �      �!#  WaG�QLD0Q�D _ �������UUUUUU��  ������UUUUUU��  �f��jfEDDD��  ������DUUDT�����j�Z�VUUUUUU��I��D41D�                 � U  � ` @      Q�QmQ������
  P* *\ �     @      �1�"  	 @U@@P�P�P�@�@U �
 	 '@'@'@	 
   U)%A�џ��'U)� T   E � � T @� � }� � 
 )����������������f&�f&�f&�  UUUUUUU  DDD  �*�*�*�*�*�*�*  �.�;�.�;�.�;�.  f&�f&�f&�f&  �?�?�?�?�?�?�?    	
                                                                                                                                                                                                                                                                                                                                                                                                  @������� � � �� � �A������ ��������?��    ?���?�?�?? � � ���������������������������      � �  ������� � � � �?��������������������?�?�?�?�?�?�?�?�?�������      �?�?������������ � ����������� �����@�  ��������������  ������      ??????????????  <� � � � � � �  �����������  �       ���  � � � ����� �  ������ � ?    ���������?�   ?��� � � � �  �?      ������  ����������  � ? ? � � ��                                                                  @������� � � �� � �A������ ��������?��    ?���?�?�?? � � ���������������������������      � �  ������� � � � �?��������������������?�?�?�?�?�?�?�?�?�������      �?�?������������ � ����������� �����@�  ��������������  ������      ??:�
�3�A؜^Ρ���R'��X�y��������,'�&7il;�,��`T��8��R��9(������l�)��m1eKIKH���[�vu`՗�1�j�jUKg�����rUe�1��jV�;���T�ڌ@��&-M2ڕ.k��\�4Z���pS��\��6k1OE���9�6�l��"��W秋�`Ƶ䬂����&�p�\���c6#i�,��S�S��9$�fdXP��;#A���&&��h��.�`�ـ�T�-�
��0�f6�h��+��a'7��q$I�.#�)J���_�q$ll��֛e�	��B�%N6�v��r��V��P�����W��Q�h��Q���b>�� Q�s���m�~�x�<��q�ֽ����oo�q��~���on?��\��n8|%��vxK����PH�3��X��m6�n�/��u�E��5��!����&�_���ēx�j�p[ d��K����q����o#�F�C��펧�`:;�t��%�O{�n�#� � ��˲�[\+;<;�����0 C]^��V�wr����]�N�>	S��7�$�RM��<R���ݶQ����O��=�Zn\�t�� �r��˰��dqy�@�"��Gq:�)V>�n���=v��䀊T��	��+�!C����E�z����ӧR�e例j؊$RЄȦ����[�'y�(7��)O0�ɓ��@��Q OX�����f��)M:�)�%U@�&R�Z>�P8� ){����NCT�Q��p��"Pcj)I��(aHs��d��j�Oc��W�M2'p���ڊjRr�e&�ܒJ�xU)�,#�Q#3�q��=�a	���)&�ԩ�aJ}�0�xE&5��@�VTx|�^H��۽��7&"�>��YVR���{����سfͫJ�Su]ʙ7*�jd��XSmxt��)�Xx����Z����Y3�IM�]�GpI���Un\������mK�N�L
�l�>M�)D�%s�#��A %?�{eE��)(F`�)�֜���5M�~ؕ:�%=P������;�EȷlJS���`�����ji��������]�T��)ۜ���ͽ���]�)�*�_�=��0o�Q��YG#�{4(Q�mb=iJ{5�kkQ{�Sk
�k��УC)N�X9M�~R�-cG��=��������)l�ٳ<2�B�:;;k��˺R���ń%�Ok=r�)7�x�{�"��0�n��B���0��a��f�z
g?<"�֘2�?�)Δ!���A�{Of)����v��.Z`9�$Wbr�����|���M�g�E]�YJ\
��{�K(���%ʁ����s��-��-Ҟ�r��1Mg�J�R��GI����Ѣ��e*x�W��X�9�C��r�L�F2���]�%!M��K����N�:T�)�6�IʘA�H�ѝ�t�TiJE���2Kir�%��HiL����pT�\�[2�H�CrH���v�4��BȰ}j�V�;)�?�R�9Y�wk�SU�U�${�	m��ȏQ:3��)��N�p{W���m��nE�)0VA�)՚��Q(r��ZR����x/����H��(�
fS�h>͔��k��{�Y��Q�����\1Ǥ�T�]Z�Jk4��"g_�Z�C^��$Ts�}-��o��N�U{�8�F<��JI�REdP��E�w+���ƨ;J_fP"�B��:<K8V0)J�)C
@�7��ϕ�iK��E�XSbͧ؏K�D�A��Js�X%ݝV}5���v��F�Ȕp)B�S��m�.LR𓄦�B��
���R|of)�ǳ~N�CQؕ_G�R�����v�Ţ�����x
l�J�����7�r�����>r��e5��d�g���K
<��Fd{�	�h�R�(��7=����Q�6��V��7J�s�8��E*���pל�6+��e.�.��G�'�lP��%9H����1J������S%1�T
g`+�qe��xJzʀ���ħ��Q�Hͱ�OV<�㓀���u�TK����@V����E���*.;r�E���k����B|;�[�'�~����&�����)X�u��'-.6�|;��2�G��T�$H�'
��Q6�f�C��4m�"��^B�*�t��N�+*v^\ƨ�\�	�j/�vM��0ȎZ�7n�����z��@��;��Y0b?��~�;��[�l�gO��(�x���^o4l^���'��Eow|R%�{����hd��2����y��gl���aI��)(��[K�y�*l*�k�� ���'��P�z��!�9�ͱs�T4��9EHp�R�[��1h"��T��%#9Ɛ��NAnlJU��x"�"�&"*��nK7���*�i$�
l���Ȝh=�E����Q/��z��F�CW:Z���p»���)"�B�ڈX�˸]t�f��;�eL��(X%�AR�JSL%b�x7�`�s�١ɍ]a�D��+�S$a�0���P̞�)DW�LZc�x�憉yV�0D��\y�xD�٤vc��0�釄*��.s?ܤ#S�)��e>X6j�*��Lda{��
Bϊ��{���l���F%%0��l���R�����mml�{�B5���a�&E?c��!��[q/m��~���7%�Q�e2D$���c������r�<�n?��5C��9T:�'�P%a�S��o�L¸٬/W `�(�k�Ѵ���c�,�m�q����NOþ_����$`�c� ���m�Z%n_��9׷[Sq��|/��ѐ�'�э��"��48"�(� �& Q�
�!l��!�"�9�	��G}��ɵ-{�:�r`,VK-��T��A�N�f���I���n�V[�6�sD��yfR�܆��P�;�<~@i$��2�8vN�ŔGߕv�i���'���!m��㎓��� 4\�������C� f��i<��n��1��0i�E噖�>���'�3@��<~(k����Ű�h1r�y:�T�vR���4�u���~���<��*NV~����\��3> �T������#$�9��g�*�C��V�8�yx��Xo�s��4���QC{�ynB~�/Xf6t�w�C
l��`���>�k�?s����A����L:2�PUهߊ��A���Gc�`0O�����ā�JzA���� �+� ��UE�R>�7kkW P� m��5��ۋX1c�c{[O״cp�!�݌on�������'�fYA�ίY��6�w1�3�z���K�����u�3�&�o������_f���Hk$��3%��,����uUʐ��=�-q�x���l+��YUG���
�5�^P49�ސi:�P6��d4��a�̀�p�`!$5/�P"�Z��~�n���q�5�_��YUC$� �lr�H���`�,Τ-��.ԃ�_iRX��u�.��u�5q@�cn: �^�eE��*� mhk�> �m7 ����ꔦ�hVځ�tU;n�$�t�LdM�4����*����;w82a�(A��ܛpAg!H�*�hk�C^�(���R��QRB9Xs�-�(���ZHM�	��	�m�	��	��	��	 4� '����hz�@���+� ��� ������m������� � � � ��`
��
m��� �s����������`L	�{1A:)z��dе��|\𩃘|���wQ( �  �Y��7�@d ��� �� ������ �󩠍  � � � � � � � � � � � �	�& ��"d#� ����/�O�o������멀� �`������_���`� ��@����'� ����0e�� e����`�


 Q��
e�� e�`d
&
&
&
&��
&e��e��@e�`H� |�hHJJJJ ��h)	0�:���H�Z�Z�Z ��z�z�z�h`8� d
&
&
&iN���e�� Z��
 ���� ��� ��0e�� e�z����8��~����`�"�NŅ�#�NŅ	F
�	F	*F	*L�F*F*F
�	F	*F	*L'�F*F*F
�	F	*F	*L:�F*F*F
�	F	*F	*LM�F*F*`        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l���  �U�`LX�� ;�� ��������������� ��L[�`dd� Z��� ��z���Z����� ��z�����`H ;���I���hdi��
&
&
&
&e��e�� �� ��������0����1����`����a�����������������	�����
����������� ����!����P����Q��```�$�%� 8�$H� �%�h`H�$E$�$�I�i�hI�i ��$$� 8�,H� �-�h`H���,
�-hJH��e-�-hf-f,��,�-`�%E)H$%� 8�$�$� �%�%$)� 8�(�(� �)�) ��h� 8�,�,� �-�-� �.�.� �/�/`� �/�.�,���-F%f$��.e(�.�/e)�/f/f.f-f,��`````��8��
��i
�$�



$`�$�%��$�fǥ%�gǐ
�%�$�fǅ$8&,&-���,�-`    
  ( P d � � ���@�E�$ٶǥ%��ǥ&��ǐ�&�$��ǅ$�%��ǅ%8&,&-&.����`        
    (  P  d  �  �   � � � @ '  N @� �8��@� 5```I�8i@�@�!���"

JJ(�I�i )?��5�(�I�i � `�� `����` 	"%(+.0369<?ADGILNQSUXZ\^`bdfhjlmoprsuvwxyz{||}~~`�)�(�JJJJ�)�
)


8�(�$�
)�J8�)�%�)


�&�)�J�'�e$f,8��jE,.�$e&8�(�,�,� �	e%f,8��jE,�%e'8�)�,�,�8``�|�$�'ɥ%�(ɥ&�)ɥ'�*ɐ�'�$�'Ʌ$�%�(Ʌ%�&�)Ʌ&8&,&-&.&/�����`            
      (   P   d   �   �     �  �  �  @  '   N  @�  �8 �� @ �  5 @B ��  	=  z ���  -1 Zb ������� ��8���I�i���8�	��I�i������������LLʰ0�Z� ��� k��e�8�����e��e � z���`Z� ��� k��e � 8�����e��e�z���`Z� ��� k��e � �e�z���`�"���H� Q��)��JJ����1�h=���` U��0����?��� ����� �� ��� ;˥8*�� *��m � �m��d�
&m��m������ �8�� ������������8� �� ��������L��`��� D˥����eɠ�� i�8��ɠ�ׅ i�`� eɠ�� k�8� �ɠ��Lk�`� �H�@�I��H����I�I�`�����[������d��������� �� �̭����������i<���`

�� ��˙ � �����`� �/ ������`������@�]�<��8�� �եHi0�J�Ii �K�������J�H���J�Hi0�J�K�Ii �K�������  _ͭ��a�1�]�-�D �բ���HȑH�� ��� �H�Hi0�H�Ii �I��ߩ��� ���_��a�Ș �˭��a�����`��`�����`���M�]�I��8�� �եHi�H�Ii �I�Hi0�J�Ii �K�������J�H���J�Hi0�J�K�Ii �K������� _ͭ��a�1�]�-�D �բ�ȱH��H��'��� �H�Hi0�H�Ii �I��ߩ�����a�����`��`



}�ͅJ���i �K�J��� �չ��eH�H�Ii �I��J�H��`�͖� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �ɍ& ���  ��� � � � � � �� � �( ����6�F�хG �թ@�KdJ�� �J����K�K�`���� ��� �ԥ)������)�S� ��L�9Ѝ������@И �Ь �GЍ�� ���NИi ��� LU�@@@@@@8  0@P`8@@@@@@p�����Т ��	�8�������p���	�i������������i����ɀ�L��d�ɴ��  ����  ����`

���Н��Н� ѝ�ѝ����i������i��� ����`	
+,)*78'(56%&34#$12!"/0 -.                   P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������)��
�`�
�����0'� ���������Z O�z�����۠ ����������Z 7�z�����ة �`����������� �խJJeH�H�Ii �I��



eF�J�Gi �K�JJJJeK�K�)�	���J���J�	�
..
..���QH�HȭQH�HȭQH�H�Hi0�H�Ii �I�Ji�J�Ki �K��L��`e���`� ����`H)��օHhJJJJ�I
eIi@}%օI` 0`��� P���@p��      Hژ��\
�h�Ph�O`�k�l� �kH
��g֍�	�h֍�	� d���(	`l�	m�{։֢ �k� �����`� �k� �����`� �k�( ��������k`� �N�:	� �N��)�� �	�c	� �	��"�� � � �( ����`dN �֢!�c	�	���(�:	�N��` ץN��`�(tN���!�	��L�֜	�W�X� � �W�O��������\� �Y�(	�	��_�`�a�N`�N�`�_��L?����`��`�`� �_�am	�`�\�
�Y�	�Y�� L/ٽ�٪�O�U�P�V�_� �U0L�����L�����L
����� �\����� �ٱU�am	�` ��Lz���� �ٱU�,	�U8�,	�U�V� �VLz����L�����	�	�	}�٨�	�U�	�V ��Lz����- �ٱUH �ٱUH�	}�٨�U�	�V�	�	�	h�Vh�ULz����' �٤_��٠ �U�.	������Ui�U� eV�V�_Lz���� �ٱUHȱU�Vh�ULz����2��ٹ0	)��0	:�0	� �1	� ��U��hڦ_�YL#� �� ��Lz�����_���)��0	)�0	�0	�0	 �٦_Lz�ɀ�(逼��

��qڙ.	�rڙ/	�sڙ0	�tڙ1	 �٦_Lzפ_�(	���٨��ٝ �ڝ �0	� �1	�  �٠ �U��hڦ_�Y �٥_
��U�O�V�P�_��(	��(	��`�^��[��[�L/٠ �S���� �^LK���� �ٱS�8	�S8�8	�S�T� �TLN�

� �ٱS��hڅ[ �ٽPڍ( �Qڍ) �R�)�* 	�* L/�   �U��V`�S��T`H���,	
�-	hJH��m-	�-	hn-	n,	��-	�,	`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   ��{ۅ���  60  0  0  0  0 # 0 # 0 # 0 # 0  0  0  0  0  0  0  0  0 " 0 " 0 " 0 " 0  0  0  0  0 $ 0 $ 0 $ 0 $ 0  0  0  0  0 ' 0 ' 0 ' 0 ' 0  0  0  0  0 ) 0 ) 0 ) 0 ) 0  0  0  0  ��  #0��������4���  :(  (  0(00   (   0 '  ( 00&00��  5 0�  0�  0�  0�  0�  0�  0�  0� ! 0�  0� 	 0� # 0� #  # 	  0�  0� �;ܻ�����  6000	0000��  # 0�  0�  0�  0� 
 0� 
 0� 	 0�  0� 	 0� 	 0�  0�  0�  0�  0�  0�  0�  0�  0�  0� 	 0� 	 0�  0�  0�  0� 
 0�  0�  0�  0� 
 0� 
 0� 	 0�  0�  0�  0� 
0 0�  0�  0�  0� 
 0�  0�  0�  0� 
 0� 	 0�  0� �����&���  :
((0&���  ' 0�  0�  0�  0� # 0��-��ޤ���  :00()�  )�  0� + �  )�  )� ( � ' � ) 00)�  )�  0�  � ) (�  '�  )�  )�  (()  ) 0 ( 0 ��  &0	 0�  0� $ 0�  0� 	 0�  0� $ 0�  0� $ 0� $ 0�  0�  0� $ 0�  0� " 0�  0  0 $ 0� 	 0� $ 0� $ 0� 	 0�  0� $ 0�  0� # 0� 	 0� " 0� $ 0�  0�  0"0�  0� " 0� $����	m�	��	M�	��	��	��	.�	M�	��	m  M  e`�	���ȑ����� ��i0��i ���L��`��ȱ����	��� ��i0��i ���L��`��Hȱ����	��h��i0��i ���L�`�	����
0�������8�0��� ����LD�
� ���	����`�	����
0�������i0��i ����L|�
�����	����`��	���
�������	`��'�����0e�� e��0e�� e���` PAUSE  `

����	� �
��7����BɎ��d

&$
0%��	���	���	���	����i�f
L�Ȟ�	��	��	��	L1�	��m�	�f
L�``H)���uhJJJJ�v
evi@}��v` 0`��� P���@p��      ```����`��� � �Z��ٝ	���ٞ	���ٟ	���٠	�L��)������	����	����	����	Z A�z��	����	����	����	����	)�	� )�z������Љ`��	��	��	��	��	��	��	��	��	)i��	��	)Ji��	�0�~d��	��	m�	:H���E~�~h d᭜	JJeu�u�vi �v��	�



ey�m�zi �n��	J�jJJJen�n��	)��	��	� ��	,�	p��m��	��0�� �mڪ�3����	��	�!�	.�	.�	.�	.�	�	.�	.�	.�	.�	��߬�	��	Qu�u���ue~�u�ve�v�mm�	�m�ni �nΓ	�L��` @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��� �y �w ���z �x ����P���������� �������o� ����������L��Ń�`����� D� =� ?� �� � �� ��L��� ������� 
�������� � ��`���@��o��`�	�� ��)m�8��� ��)m�8������八 �Ưح�������d� ���`	
��JJJ����������
������������ ��`�  ���`�  )���8��ɠ����  )���m�ɐ����  )���8��ɠ����  )���m�ɀ���`��
��������公������������ ����������
��"��#���� ��ƫ�`���ɠ�����ɓ��o� ���������`���6��`�)�`�������`  �  )�`��
��W��X�l c�����楄�Ƅ`��0��`���������������� ���� LX�`�� �o�`����
������������'��(����q����q����� ������� LX�`�	�����





   �!�����      � � 3�3�9�9�9�9�      ��
��������u��v��� ��q����q����`�����������������      �� � � ��������o����������`��`����)����)��������� � �� �� L� ��`���� �ɀjɀjm�i���� �ɀjɀjɀjm�������8�D��` 	�)������i����ɠ���������ɠ���������)����������
�������� ��`�  )�`�����o�`������������`����0`��iɥ���`�o��`���i
�����������������
��"��#���� ��```�� �����4�2�0�.�6�8��������o�\���Z�[�]`��Y�`�Y �� c� �L��`��0`�\0`�������Z��[�	�"�
���@ vȐ�o�\L��`�^���#��������`�����`������`���
���`�\`���Z ��)i�[)�^)i�]���\`�Z8�]ɠ��Z`�o�\`�\0���Z�Z��[��^
��;��<��?� ��`C�E�G�I�����xآ�� �� �֩��	� ��	����� �� �� ��I�& �'�� �  � ��  I����	�&  3�����d�
�e�f� ��	����� � �� :� i��`�ȍa�b�5�� ׭`��`������0
���� X� z� ��  )��v �֩` Q������� Q� �� �"��#���������� Sŭ  )����H�e�� e������h��  )����  )��� �֩� Q������` Q� ����o�[����I�&  �� ��Lo�I�&  �� "� ���H��e�� e������h��	�& ���������`������L���0w�@�I�& ���� �� Z� � q�� ׮_�� �_ �� ������	�& L��b� ���b�H�e�� e������h�L��_�R��H��P��@�a��a�H�e�� e������h�L�� K� 않H�e�� e������h�L�� ��L�� b�L�� H� ��  )��H�e�� e������h� ��  I�����d�
�e�fL��e�Lo��d��e��fL��b��?� � � � ��� ��	����� �� �� ���"� �#���
��b��� S�` ��)�" ��)�#���
��[��� Sŭ���LX�`DANGER        ���� ע ��	����� �� �� ��_�������  �L�� *�L�� �`��ȝ����������g�{���`� ڎg �� -������`�h�| ��g���|����hH�d	
&	
&	
&	
&	��	�

&
e��
e		@�	hH �hHJJ�h)��)�Q�`0��g��d	
&	
&	���8������	���  ��)�p�)?i ������ ��)i��`�&�'��^������d� �� ��  ) ��&���'�'���` ��)i� ��)?i�	�2����01������u�	� �ߝ� ��):�� �ߝ� ��)::�c�����`d������ �����` G���}�����}u�uɠ�Z��}7�7�c}��x�C�
}���� }c�c� Q��u)
��~���	�uJJ� l�i/��Q�ȥ	Q�`^�` < � ��������  �L�� *�L�� �`��ȝ����������g�{���`� ڎg �� -������`�h�| ��g���|����hH�d	
&	
&	
&	
&	���i#��zr�L=����(��fR���0Y�*TG�C.���A����4�z�hŤ�F�����ű�����G����-�*�ƌ3i��IO�˒s���1��;�݀�]�ZB����݈�{����)��4�����4z�i��肽�M���}Ɣ��iC�|�A��M!OkԌ�`#@�z����u��i��A�d���k�EviX�-9����0m�k����2�Rk�j�9��4^�B�I�����KK�hQ�v�: C�n{q����o/��4�|7S����oa��F��B�gANֹ�˕lk�Zb�YZzm|�k+�[,M~�p��4)b"�2�� �c�%�מ`-2۷��Fy����Y�<:'��7�5<��KG��@հC͵ߺ5]�ҭNl���	]V 1�90,{�n�h´�U�5(����
�B˗}� K;^��\#�	X̏�i�c��;#^%#�)l����@2akBk؍	L���A��t�
�`oH���ki�I����EqQ\x^S���g�@mt�+�h+?i4�7���_@�����Ӛ�֛t�Wi���W?�)�y�-�Uz֒S�W���I�lW�OqY���Ɗ`�73k��[[�x�.�̴�Ɨ�Fb�#Fk�-,�_��i1�ZO)�/N�V
��1�u��^-�^�d�5�t�m�*"l�,��J�Tki=�m�cD�Ze;It%�p��ڳ�N�J�VG����A�^�z&�R��ٵ�^�h
O)��'��ˀ��)���1=�.Pf�g)�J�a�pc]VcAz0��h-v��^5^s<0�����Դ��1��[.N�BQޗ��5������3�D�^�h�����4�� x
��T��z,4���Rґ1��f�E�]��Ӄ!���j\�l��dO��sBk���iS7k  5��VVf���e4G�Ȧip�D>cYS��C��Ӭ8So����+D���e�����M��C�������y庘ފ����T�Ⱦ0�9=�xSX�:/�Mן�a�2���/%�YT��	���h�Re��Wr�H��p�"�fR�͟�fĴ�i��aV�,�qX�"����ea�o�Hͦ�g�h&�\h\h�4Y����Ϡg��hMRh7.�8��K�F�o*����hCp2ѫ>;��KR4�a�^%��N����l�5j��wv���G��I�i4#E?:K���lv�Zm��֎�0kv�i��$�<�?<���3Jdn���>#A5�p�KF��i���N����!S���6�&cmB3a��4��b�R2c�1�3�d�l�#�5��A�^�.<�~2��<GBYo�b`MU��k�f�Fr3�C����w��_2��:����0����$����i��7�!�ܵ\�@)���M�I�]��<�p#&��C3V~#��L��r��GS'KJU�Q��&X8L�nǢ1�F� e��$8�չ�&H��5R4�r�x'g4?���|���ՙf*�|�\��ͶHU��M�l�0D�X=+*ͭ�aZW¿5`��Ƒ:�34��!��L�_?�rZ�ʉ�i4�g���H��g���a��V��c1�e�P��ɒ[���p,g+���-|��~�4����h���w��+I�h��k^�c��婬�/��1�q��R8�k����?n8��|x��N1z^15#B�#ڵ�|�U��������$��k���K�i���Y�|M8HψV�}�
����;u��?q�-L4�Btyyo���Q������ыH��Y.h��;F�"\��4���h	�pxs*s��.��:��h�5�-͉I��t��OO{�i���M(2����A�O�(7�1�s��s�S;��D҆Ix�0?�PMpM/Q8m��Ԁ���8����Y��6��I�l=<3a�j��/�.Yh)���Qz�f�dF��1N����K��q�C)O!�����Q�uno�\"Ԧ�q�:�2�>���@�Vhk7ay�K���*�Y�����f��J&�M�x��qkVR���r��i~r��`��#�5������O�Ӎ��Bk�j	��->��+E��KPr�f9֎#Y�i�9L�-h���U�M_��YbZg�䞎v�x�2*"{�b�-���"��m��?Y�-\擛AS�0�kO�E�1��QGnZG�~Z�U��<�R����&i��'I��m'���|L1#>p�?��灘��1n�V���AZŭ[��cw�?�4�A,�g�	��&�4���ӎ|����A1���a3��3,}�C25o� `}J${׵���;�G�$o��m&�I�QH�J~~L���<������(��I��rI��%�M$���P6�������vkmj|��l����>'�,_ҡDX��B��
��j���͠�aE�6^�
�}G��p� ��D��Z��`���*~ņ�:'t'��[�/�0V�^�{L;uݣ8���]���7d�����v�u����E���U�Z�j�]Mssi�Z���շ���˟�x@(�sT�Zt6�|D.�孽��v��l���@�gO�{��C���Gb��u���*t��J����f��E	.�}buv>�k�[ug t�@��MDWZ�ve�'i��ݥH�:���EjW�K������Ҥ��n�����,���X�]�k��!6�mR�n�F�7n��}מy�q�9��L���]p�|���mc8�I��C�t��
6���!������G��{���m�
�z��B����r�.�f�u:�M]b;s}%�-�}\�� �SP�u��\F����7��ǇèG!�<8��C0��}n8'"v��M%�>{�x<]5f��~{3��)ӎ,���Ά��Ύ̼��6�\��Ô[M���å2뜶f��� �X�t���>Ӵ1���s�8�a8�=����� �'�tm����\C�Ł��@v�Su�F�i]^&�c��k��óz�Ϥ��_[K�q�-����br���zX"nK�<膞��ٖiM��5�7�3s�
�MgIy���OQ��Q��ZeF� ��
�}gP�[Ԍ��Z�'�j�u�� �����R<��fa:���1[3���T)=^�|�W�5Դ���em�^�W�S[�0Cں�l2O2m���#�B
8(;,�o�gG:ͿT�D�Q���;#�3J�����0b��[ʺ����
�����	�}������L��u<�e'�&_P��Tpf��N�,r��k.Oa��+�a���uy��kk���HӚ���@6e�x���,]���F04+��Θ�n5uz��A��2�:/�}�o��WP:�둅Ҿ����:	szۋ��T����p�J���º�f�|���e�z3�a�8Ά{w�·�:e�����jO���':�:_!�E�j�Rr����tӖ�b+�ۋ�p\�2�;&�Gp��e]F\}}~��_,�,9Vmh��ֺ���N�~���I��f�ŀ:�}l�$�ʙ�:��\
������V3�]GOK�w�3�Y����`�~��u��>���}���Vk��%���q���1ղ�3�p�C���V=����~��T��@�T\o�=a���BK�C�u|��J��4��x�h���Z�PARK    COM            ��U�  CONFIG  SYS           OUHH U  386SPARTPAR&          ]CI	�  0 PM                   ˎ/�0    TSM     CFG           i=S[�   WINGAME              v�B M    �                    PsE�J                                                                                                                                                                                                                                                                                               �K��