                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �
  ���
�
�
����      8     888        �     ���  >>      �     ���  >>      �   �������>>      �   �������?>      �   �������?>      �   � ���  >      �   �� ���* >      �    ��� � >      �    ��� �>      �   ������>      �   ������>      �   ������>      �   � �
��  >      ��* ��
(������
      �   8� ��    8      �#  ����  >  �      �#  � 
�?  >  �    ���꣪�� �����>����    �������� �����?����    ������� �� ���?����                                                                                                                                                                          ����� *������
���
��* 
 
�� �#��8 �#8 �  8�� �#��8 �#8 �*�*8�⨊����( �#8���/��8
�������� �#8����8(� �����"�#8 ���8�� ���� *�#8 �  �8��� ����(�#8�
�  �8�� ����( �#8 8�  �8�
� ����� �#8�:�  �8�+� ������#8�?�  �8��� �����
�#8 ���8��� ����8+�#8 � �*8��� ����8,�*8�*�* 8�� � ��8  8 � 
 :�� � ��8 
 : પ��>�� ����:���>��������� ���?����������> 8��8��8��8��8��8��8��8��8��8��8��8 8��>��   �� �� �� �� �� ��0�� �� �� �� �� �� �� ����, ��������> :�*8��8?�8 �8�+8�8�?��? �?��;�:+ 8��>������> 8��8��8 �8�8��80 8��8�8 �8��8��8 8��>��    |  �  � �5 �5 p p�\s\s�p�=WU5�= p p p p �����: 8��:��� ����: 8��8��8 �8��8��8��8 8��:������> 8��:��� � ����> :��8��8��8��8��8+ :��>�������� ������� � �� �0 �8 , ,  ��������� � ��_U=��5' 6' 6' 6' 6��5\U����5' 6' 6' 6' 6��5_U=���� <��0# 2# 2# 2# 2��2 2��2 �2 �2 �2��2��2��<< ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ����������������������������������������                                      �                                      �                                      �                ��                   �                <                    �                 <                   �                0�                   �               ���                   �    ��        � ��                  �    � �        � W                  �    ? �    ��?��U                  �   �  <   �UU����                  �   �   �  �WUUU����                  �   0   � UUUU����                   �   < �� �UUUUUU��                   �    �� <�UUUUUU5 <                   �    p�0|UUUUUU� ?   �              �    |U�_UUUUUU��   �              �    \U=�UUUUUUUU�    �?              �    \U��WUUUUUUU=    ��              �    TU� WUUUUUUU�    ��              �   < \U�WUUUUUUU�   ��              �   0 |UU_UUUUUUUU   ��              �   0 pUU\UUUUUUUU=   ��              �   � �UU�UUUUUUUU� �+�              �   � �_�\UUUUUUUU�? �U� ��           �   � \� \UUUUUUUU�?|U9�?            �     �? \�UUUU��UU=0_U�?             �        \UUUUU��UU��U              �    <    \UUUUU5�U @UUU              �    �    \VUUUU5�UUU UU����           �    �   \UUUUU5�UUUU        �      �     ?   ��UUUU5�UUUUU�       �      �     �   ZUUUUU%�EUUUU���      �      �     �  ZUeUUU��U  T� �?     �      �      ��VVUUUUUPUUU5  �    �      �       ��gVUUUUUUUUUUU ��   �      �       ��YUUUUUUUU�WUU ��          �    �� ��ffUUUUU��UU ��        �    ���kZU�UUUU��UU ���        �    �� �UZUUUU���U� ��       ��    ��> �Z�UUUU��U�  ���   �   ��   ���: k�fe�U��  pU=  ���  3 �   <�   ���? �jVUUU�    pU=  �*�  � �  ��   �; �YfVUU5    \U ����  �� �  �   ���: �UUUU5    W� ����  � � �� �   ���� ���YVU5    W�  ���?  3 � 0 �   �����jVUUU5�� �U=  ��� 0 < 0�� 0 �    ��� ��jUU50 ?�U  ��:   0�  �    �> lfVUY�0 �pU ���    0�  �     ����Z�eU�� �|� ���  0  0 �  �     �����UUU���W�  ���  �   0 0  �     �� _�ZUU �W=  ���      �    �     �����Yi�U?�U ���:            �      ���?pUeUU��UU ���:            �      ������YVYUUU� ����         �   �      ����eUUVUU?�����   ��   0   �      ������_�eU��������   ���      �       ������_Uտ������:   ���?      �       ����������������   ����  �    �       ����������������   ����  �   �        ����ë���������    ���  �   �        ���?���������>    <<�   ?  �        ���3���������    <��    � �         �: ���������    ��0?    ��         �?  ����j���    ��3�33     ��          <  ��jjZ���    ��3�33  �����          ���������>     � 3      �          <�����j��     � ? 3                 𬪦����      ��� ?                 ?���j��       ���      �          ���j�ڪ�       000��     �            ���j���       �0000�    �          <  ��j����       ��     �          �  �i�����       0 3     �          � �������?      ��0�0    �            l�������      ��<0    �           (�jZ�����     �� ��   �           ���ꯪ�>      0 �     �           � ������:      0? �    �           <2�����      �0 <�0   �           02��      ������   �           0
2�����      �   �      �           �0 ����               �           � 0 ����   �   ��� �      �           �< ����  < �   �UU�?      �              ��  ��    WuU      �            �  ��  �?     W}U      �                ��         ���      �                ��         ��       �                ��         ��       �                ��         0��       �                ��         ���       �               ���>           �       �               ���:                 �               ���:                 �               �:                 �               ���:                 �               ���>                 �               ���                 �               ���           �       �                ��                  �                                    �             ���?  ��� �  ���      �       ���    �  ����  �|U      �  ��� ����? �? � ? ��?  �\U5      �  �� ����?    ��? �?�?  � ��      �  ����� ? �? �?�  ��� �� 7��      �  ����� ?    �?�  � � �<  \     �  �����   �? �?�  � ��<  p     �  �����      �?�   � ��  �     �  �����   �? �?�  � ��  �     �  �����      �?�   � �� 0 �      �  �����   �? ��  � �?� � 0      �  ������      ��   � �?�   �?      �  �  ���   �? � �  � ���           �  �  ?��   ���? �   � ��<           �  � �?�� ? �? � �  � ��<           �  � ���� ?    ��   �  �           �  � ���� ? �? ��  �  �           �  � ��� ?    �?�   �  �           �  � ��� ? �? �?�  �  �           �  � �����?    �?�   �  �           �  � �����? �? �?�  �  �           �  � ����    �?�   �  �           �             �? �?�  �  �           �                �?�  �  �           �             �? �?�  3  �           �                ��? �3  �           �             �? � ? �?  �           �                �  ��� ��<           �             ���?  ���               �                                      �                                      �                        ��� ��?�����        �         �  ��?� � ������                 �  ���� ����� ��       �<         �  ���� ��?�?� ��       � 0         �? �� �� ���?�  �       �0         �� ��? �� ���?�  �       �<         �� ��? �� ���?�  �        �         ���� �� ���?�  �        <          ����� �� ���?� ��        �          ����� �� ���?����       ���        ����� �� ��?  ����       ���         ����� �� ���? � ��       � ?         ����� �� � �� �  �       ��         �?��� �� � ���  �        �        �?��� �� �  ��  �        �?        �?0�� �� �  �?�  �        ��       �? �� ����  �?�  �                   �? ��? ��?��  �?�  �                   �? �? ����?��?� ��                   �? �� ����?��?� ��                   �? ���? ����� ��                   �? ��� ���������                   �? �?�� �� ��������                                      �����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     � <                  �?                  ��?       0          ��?     � <      �  ???     � <     ���  ?�   �<     ���� ��   �<     �� ���  ��<  � ? ��� ���?<  �� ? ���0� ?<  ��?���� < <?? ?�?�� < ?� < <<� ������ <� < ?�� ����?  �� ��� ?��?� <   � ��   ?��0 <      ��   �?�   0 <      �?   �?   0 <            ?                 ?                  �<                   �?        0               �       �       ���     ���   �����?   �����  ����  ������ �?����� �<����?��<����?� 0����?<� � �<�?�3 �� <�|2 �0<���  3��  ������  ���?0  3��� �3����   ���?   ����   ���?   0�����   ��< �  <�3 � �� < ��0�� 0 3    < 3    0 �  �� �0 �0��  �� <     � �   �� <   ��3 �    ��   �  ? 0   � "�  ��� (�  ���" 
 ��� �����3 ��� << ��� 0 ��� �����   < ?    ��     <�     ��      �      �   H�Z �� � �� i� �� p� �� �ޜ] �� ��  �� 2� �� �ĩ"��  UĜi  �Ʈ� ����i  �ʜi  � 
�i  ,� ���i  �Ȝi  J� � ��i ��
� �� �-0�z�h`H ���E ��F �v�B  q���E ��F ���H � ���E �(�F �c�B  q���E � ���E �<�F �d�B  q���E � ���E �d�F � �� � ǭi ��^ ���� �� �� �� �� �� �� �� �U �[ �\ �] �^  ����� �� �� �� �� �� �� ��  ��  f� ئ�i ��L,��i h`H�Z���N � �� ��= ��< ��7 ���� �� �F �7 �E  ��� �r� �Ε ���8 ���� Ε �� �F �7 �E � �� ��< ��=  �Ζ Ζ �� �F �8 �E ��= ��< ���  ��� �D� �LU� � 譕 �F ��< �7 �E � �� ��=  C��7 i�7 �E  ��8 �E ��= ���  C��8 8��8 �E  ��8 �� �L�� T� ��	 ��z�hX`xH�Z�� 
��S��� �S��� �< �I �= �H  g�z�hX`H� �N  ����N h`W�������? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                                 ��    ��  ���  ?���  ��_ <�? < |�  ��  ��   ��  �� ���
  ��  ��?   �?   ��* � �"   p?    �*   0*�    (�    �    �    �  �    ��   ���    ��    �  "  �  ��"�� �� �(����"�� 
 ��!  � �*       ��  �(�  ��
�  � �� ��  � ��  � ��  � ��  � ��  � ��  � ��     �   �
              ���         ��    ��  ���  ?���  �� <�?? < <�  ��  ��   ��  �� ���
  ��  ��?   �?   ��* � �"   p?    �*   0*�    (�    �    �    �  �    ��   ���    ��    �  "  �  �� �� ��(�(�� �"��""
 ���  � �*    
    �
    �    �    �    ��*   ��    ��    ���   ���    �  ��    �  �
     �    *  ���    ��   ��  ���  ���? ���� ?<��0<0��   ?0   � ���� � �(  0   0  02��?<�0 ���������?�??       ,  �   �    �*�  �   ���  � �  �
   ���   (�    ��  (
��  � �  � � �����  
`*  
    �   �    �     �     �   ���   ���   ���   ���    �    �   � �   (� 
 ��    ��   �
� ��U�� ��    ��  ���  ���?  ����  ?<�� 0<0�� ?�   � ��*��  ���  �/� � ���?�����<�����  ����?�?? �   (    �*   �    �      �*   �   ���  � �  ��   ����   ��   (�  (���   ((� � � �����  
 (  
    �   �    �     �     �   ���   ���   ���   ���    �    �   � �   (� 
 ��    ��   �
� ��U��    � ���?  ����0���� �����@��( @�? O �?0�| �?�| �?�| �? �?    �    �   �  � �  �  �       
   *�   ���   ��    ��  �   ��
  �   ��* �  (   ��*  �  (  ���* ��� ���� "������������(� �� � 0   � �   �     �<  �0�  0�  �< � � < �
  �" (�� 0*��� �*��� ��jP� �� T ��   �j    P           � ���?  ����0���� ����� ��O   �? O �?0�| �?�| �?�| �? �?    �    �   0  � �  �         
   *�   ���   ��   ��  ��   (��
  (  ���
  �  "�
 �   ���
  �/ 
  �    ��� �� ( ���   ���  �>*, � 0�
 �    �    (    
   �
     � * ( �� �� � �
  �
  �*  �"�� ���"	���"
����
��BUUTU   �?     ���� �����  ���?�����  ���  � ��  =� =�� =���� ���   ��   � �  �? �*    
     �   � �    �    �   �
  ��*  � $*  ��
      �  ����  ( �  ���  (   ���  "�� @��� ������0���?�0���?�0������?�?� �             (    �  � �  �  �(� ���� �� 
� �� �� �� �� �� �� �������"������ �����`PUU��*   @U�?     ���� �����  ���?�����  ���  � ��  =� =�� =���� ���   ��   � �  �? �*    
     �   ��    �    �   �
  ��*  � $*  ��
      �  ����    �  ���       ���   ��� ���� ���?� �����  ��?�  ��?   ? ?    ?       �   � �   � �    
   �   ;         �(    �*   (�*  ���*  ���  ���
  ��V  @U              U��UUUU��WUU���_UU?���UU��_WU=�U= |�U	 ��U	 ��U% ��W% ��W%���W
  ��_	  ��%  X�%  X�_�* X�WU�bUUUu?`UUU��jUUU5 �UUU	 �UUU	 �UUU	�UUU	`UUU�(�UUU���UUU��UUU	
hUUU�UU�� �VU%��AUU
*`UiU� XeUdXTeU� F�jUU�EjUUU��aUUU%�UUU%
�UUU%( VUU%� VUU�� �UU��BVU��� XU���`U��U	�U��U%�UU�U%�UU�U	`UUV	XU� V	X� VV� �VV��ZU�UUUUUUU ��    ��  ���  ?���  ��_ <�? < |�  ��  ��   ��  �� ���
  ��  ��?   �?   ��* � �"   0?    �*   0 �    �    �   �       �(�   ���   ��   
(   �  �� �   �  
* (( � ��" d�  � "�* 
� *   ��     �    
�    (    �   �� �  �� ���  ���  �� � ��  �  �  �  �     � � � ���
 �        ��  W�
 �U�
 �U� �U� �U�   W�
� �
  �**  �*�* ���* ���
 ���  � ��  �*  �?  �
  0��  ��
   �   �*   ��  W� �U�
 �U� �U� �U�   W�
� �
� �**  �*�* ���* ���
<��� � �  À*  3�
 0�? 0�
 0��
 ��
   �    �      � ���?  ����0���� ����� ��   �? O �?0�| �?�| �?�| �? �?    �     �    0  � �  �         
   *�   ���   ��    ��  �   ��
  �   ��
 �  (   ��*  �  (  ���* � ��  ���  �� ,�� ���	 �� � �� � 0   � �    �        2   ���   � �    �        (    �   ��h   ��j
  ���
  ���
  P��   @U             �?     ���� �����  ���?����� ���  � ��  =� =�� =���� ���   ��   � �  �? �*    
    ( �     �    �    �   �
  ��*  � $*  ��
      �  ����  ( �  ���  (   ���  *��  ��� ������0���?�0 ��?�0 ����0?? ?�   ?       �0  � 0�  � <� 0 � 0�� �3 <� 0< �� 00 ���(0 ����  j��
 ���* ���* jP�*   �    T          ��    ��  ���  ?���  ��_ <�? < |�  ��  ��   ��  �� ���
  ��  ��?   �?   ��* � �"   p?    �*   0 �    �     �    �         (�   ���   ��   �
(    �   � �  ��   "  ( � �
"  ��  � �*  � *   ��!    �    
�    (    �   �� �  ��B ���  ���  �� � ��  �  �  �  �     � � � ���
 �       H��m� �� �� i �� �� i )�� � ��h`H�)�E � �F �%H�)�E ��F �H�(�E ��F �H�*�E ��F  ��h`H�@�� �(�� �%H�B�� �h�� �H�@�� �+�� �H�B�� �k�� ��W � ���� i0�� �� i �� �W ��h`H�Z�8� � �
��.���^̠ �=�̠ �A��̠ �L�=̠ �.�̠ �7��̠ �8�3Ș8� � ����& ���! ��� ��� ��� ʚ� ך� 䚀 �z�h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<3<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                        �?�?      ��_�W�W�����?����?���?����? 0 ��? �<        �?����<<�? ?������
�� < �?�����
�:�2<  �?ܷ��
��< ? 7��ޠ���
00 < ���(��
���ʀ:� ���(��
���ʃ:�? �
�(�����0? �
�(������������������������?�?����>�*�*�� <?�?����>�*�*��< =�?������.�
<� ?�?����˸��< � � ׀����*�*��
 � ׀����*���0<� � ��è�*��
� � ��è�*�<         �? ��� ������������P�_�U� �U�  T  ?   �                  ��  �����������@��@� WU WU P  ��  �                   �? ��� ���p�_pUUP]]P]]�U� ���  T  ?   �                  ��  ��������UU@uu@uu WU WW P  �� �                   ��  �������� U� ]� ]��UU UU �U  <� ?��?              �? ��� ��� ���@��@��@W�pUU@UU ��  �  �  �              �? ��� ��������U ��u �u PUU@UU  U� �< �� � �             ��  �� �������W����_��UU UU �W �  �  �?     ?   �   ?   �         <   0   0   �   �         <   0          <   0   0   �   �   �         <   �   �   �        ?   �   �                      � < � �� �?             �Z �� ��� �E ��F ��C��� �C��� ��H �m�I  g� �� �� � =�z�`H�Z�E ��F � �C��� �C��� �(�H ��I  g�z�h`��  �� �� �� �� ���  ��`L$�������`ڊ
��G��� �G��� ��E �L�F ��H ��I  g��`     �����������
           �����������                                     � �ꨎ�              ��:�:�         � �਎�              ����8�         � ��8�              ����8          � ����              �〃�:�         � �88�              �〃�          � �����              �����8�         � �����              ��:��8�         �                                     �                                     �      �����������
           ����������� ���� ����  ��8   ���  ���8   ����  ���                         �������*                                                                                                                          8��88   ��8�8   ��8�8   ��8�:   8�88:   8�888   8��88               �#                                                                                                                                  �:��:   � ��:   � �    �:��     8�    �:��:   �:��:               �#                �������*                                                                                                                                                                                                ��:��� ��:��� ��   ��:�  �� �  ���?  ���:                          �������
                                                                      પ����
xH�Z�B �a��$L;��b��%L;��c��&L;��e��(L;��f��)L;��d��'L;��g��*L;��h��+L;��i��,L;��j��-L;��k��.L;��l��/L;��m��0L;��n��1�F�o��2�>�p��3�6�q��4�.�r��5� �s��6��t��7��u��8��v��9��w��:��@��> ����? ��G �F ����@ ����A �E �>-N �@�> Ȳ>-N �@�> ��G ��z�hX`���N �#�E �z�F �v )�B  q�`H�Z���N ��E ��F �� )�B  q��E �E ��  &ꭘ  &� K�z�h`���N ��E �d�F �� )�B  q��E �E ��  &��  &��E �n�F �� )�B  q��E �E ��  &��  &��E �x�F �� )�B  q��E �E ��  &��  &�`���N ��E ��F �� )�B  q��E �E ��  &꭛  &�`���N ��E �d�F � ���E �n�F � ���E �x�F � ��`H�  ���� �h`H�O �  ����O �0�h`H�Z�� � �Lw��E �P�F �  �� x� Э��L��F � �b�B  ���G��E  �� �� q� �ƭ  ������� �� �� {������ �� � {������i  {��7��� ��� ���� ����� ������  ����В {�����  ����z�h`Z�
��O��� ȹO��� ���B i7��z ��`H�Z�
��O��� ȹO��� �����b�8�7�B z�h`H�Z8�7�I �B �a�
�I �B ��A8�7�B ��a�B h`H�A8�7�I �B �a�
�I ��B ��Z8�7�B ��a�B h`H�Z�� �� 0N��� �� 0D��� �� 0:�� �� 0P��� �� 0F��� �� 0<�� �� 0J��� �� 0@��� �� 06��I �� ް ���b� �� ������� �- $��b� �� ������� � �� ��b� �� ������� z�h`�� �� �� �� �� �� � �� �� ����`�� �� �� �� �� �� � �� �� ����`�� �� �� �� �� �� `�� �� �� �� �� �� `�� �� �� �� �� �� `�� � �M�� �P=�@0�0#� �	�@�I �P�2� �I �(�)��I �� ��I ����I ����I ��� �I `H�Z �� ����E ��F � ���E �1�F �	 ��	�E �� )�B  q���E ��  &�L�F �
�E � �� 7�H�H ��E �I  &��E �H  &� �ƭ� ��L�F �
�E �
 �� ϴh�H � �� �� |� � ��H �� �� �� �z�h`��W �� ��  �� h��W �� �� h� ������`ک�H ��I ���N �0 �� �� �� �é. �� �� �Ɯ* �  ���`H�Z�i  �� ��.�K  � #��  ��L�� ���0��	�2�K  �� �� ���i ��L�� �����W � �� ϳ ���W ��i ��L��� �	�<�K  =��i ��L�����.�K  �� #��* �  �� ����� ���	��<�K  =������W  ϳ ���W ����B�K  �� �� �Ƣ�2�K  �� �� �� �� `� �� ��z�h�i `��H �8�I  �� ��`��H �8�I  �ĭK  ��` ��� ���K �K �K �80�2�K `H�Z�K H��	�8�K  �� �� �Ʃ:�K  �� �� ��h�K z�h`��H ��I  �� ��`��H ��I �K  �� ��` ��� ��K �K �K �20�.�K ` ϳ ��� ���K �K �K �B0�<�K ���`� �B�K  �� �� ����� ���K �K �K �H0�B�K ��`H�Z�K Hi�K ��� ��h�K z�h`��H�K  �� ������K �K �K �N0�H�K ��`�� �.�K �0� #��0/ �ƭK H�Z�	���� �����K i�K  �� �� ��z�h�K ��z�h`H��E ��F � ���E �A�F � ���E �n�F � ���E �(�F � ���E �U�F � ���E ���F � ��  ���h`��?< �� ���������?< �� ������� < <    � �?��? < <    � �<��< < <    � ����� < <    � ����� < <    � ����� < ���� � ����� < <    ���� ��� < <    � � ��� < <    � � ��� < <    � � ��� < <    � � ��< < <    � � ��? < < �� ���� ��� < < �� ���� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �* ���ة��  ��� � �S � � �T � �ߍ& ��" � t ����> ��? �� � �>����? ��� ��XL �H�O �e �f �g �h �a �Q � ��Q  ��(h@H�' )��O �a �e �f �g �h �R �# �$ �% hX@                                                                                                                                                                                                                                                                                                                                                                  O���N  � � l���� k�  f� ئ�i  �� �� +��i  �Ʃ  k� �� �� � �ɭ� �� �� �i �� �� i� �ޜa �� �� �U �[ �\ �] �^  p� �� �ޮ� ��  �� 2� �� �ĩ"��  Uĩ��i  �� � 
� �� ,� �� �� �� �� J� � �� � �� ,� �� Jɀ�H�  ����i h`H�Z������ �����  â � ���C���-N ����H �� �íG �H ��I ��z�h`�H �G �@�� � �� �F � ��� i0�� �� i �� �� ���E m� �� �� i �� �(�C �@�D `H�Z â � ��-N ����H �� �íG �H ��I �� 1�z�h`�� i0�� �� i �� �� mH �� �� i �� �C i0�C �D i �D `H�Z�F �H �G �@�� � �� � ��� i0�� �� i �� �� ���E m� �� �� i �� �(�C �@�D � � �C����H ���� i0�� �� i �� �C i0�C �D i �D �G �H ��I ��z�h`H�Z��H ��I ��  ��z�h`H�Z��H ��I  ��z�h`H�Z�
i�ʎE �


i��F z�h`�i � K��J �J �
�-�J �I ��H  �Ʃ�E �(�F ���N  gé �N  g��J �̭� �%�+ �Ʃ�E �� i(�F �
�I ���N  gé �N  g�� �Ω	�J �J � �/ �Ʃ�E �(m� �F �J �I ���N  gé �N  g��J � �ʩ�J �J �
�/ �Ʃ�E �(m� �F �J �I ���N  gé �N  g��J Ά �ʭ� � �& �Ʃ�E �� 8i(�F ���N  gé �N  g�Ά �ө(�F ��E ��H �/�I �
��U��� �U�	�)��� �I �J �F ���mE �� ���i �� � ������H 0� ���� mH �� �� i �� �J �ǭ� � �
��
�L"Ǝ� �� �� � �2i
������ ���	�)��� �d�F ��E ��H ��I ���N  gí� i
������ ���	�)��� �d�F ��E ��H ��I ���N  géߍ& `H�Z�
������ ���	�)��� �� � ��� i�� �� i �� ʀ�z�h`H�Z � � �z�h`H�Z��7  ��7 �� ��z�h`H�Z� �ƭ  �����z�h`H�Z�x ��u ��i �� �� ��l �m  ��[ ��R �������[ �D�x �w  {�����} �|  ��| �} ��} ��  ܭ� �} �w �x �j �l �k �m  �� >� �� ��z�h ��`H�Z�V ���t �u  ��L%����t �u  /�L%����t �u  �ЀJ���t �u  �р;���t �u  È,���t �u  ��L%����t �u  Ѐ��	�t �u  d� ��z�h`H�Z�y ��x�i �� �� �� �� ��n �o  ��\ ��R �������\ �D�y �w  ������~ �|  ��| �~ ��~ ��  ܭ� �~ �w �y �j �n �k �o  �� {� �� ��z�h ��`H�Z�z ��x�i �� �� �� �� ��p �q  ��] ��R �������] �D�z �w  ������ �|  ��| � �� ��  ܭ� � �w �z �j �p �k �q  �� �� �� ��z�h ��`H�Z�{ ��x�i �� �� �� �� ��r �s  ��^ ��R �������^ �D�{ �w  ������� �|  ��| �� ��� ��  ܭ� �� �w �{ �j �r �k �s  �� �� �� ��z�h ��`Hڭ� �0��� ��� ��� ��� �F�
0��� ��� ��� �� �.�0��� ��� ��� ��� ���� ��� �!�� ��� �h`�� mG 

�08���͟ �i�� mG 

�08���͠ �i�� ��`�Z�e �=0�` �e �` ͋ 0���� z�`�Z�f �=0�b �f �b ͋ 0���� z�`�Z�g �=0�c �g �c ͋ 0���� z�`�Z�h �=0�d �h �d ͋ 0���� z�`H�Z ��; � ��: �: �� �ட �� �c�B �i 	���� ��L�˭i 	���� ��L�˭i 	���� W�L�˭i 	���� W�L�˭i 	���� ��L�˭i 	���� ��L�˭i 	���� �L�˭i 	���� рG�i �� �� ����z�hL�	���� �֭i 	���� ׭i 	���� �֭i 	���� ]� �Ʃc�B �V ���t �u  E�L#����t �u  ��L#����t �u  �L#���	�t �u  d� n� ����i z�h`H�Z��� � 2� q����z�h`H�Z��� � 2� q����z�h`H�Z� ��e�B  2� ǩa�B  2� ,ȩ ��e�B  2� �ȩa�B  2� Jɩo�B  2�z�h`H�Z� ��e�B  H̩��i  ǩa�B  H̩��i  ,ȩ ��e�B  H̜i  �ȩa�B  H̜i  Jɩo�B  H�z�h`H�Z��,� ����5��� nՀ.� ������ nՀȩ�U  È��Y ��U �  `̀ ��z�h`H�Z� �� v���� ��L�ͩc�B ��]� ����U� S���� =Ո '� 8٩d�B Ȉ��V  2� q��t �u  ��� �� 2� �ۭU ��"� �� �� lĩ��  UĜU �� �V �t �u z�h`H�Z vҮt �u ��^� ����V��� �����g�B  2� q���V ȩc�B � S���� =Ո '� 8٩d�B Ȉ 2� q��t �u  ��� �� 2� �ۀ�* �  �� �_ �V �t �u z�h`H�Z��,� ����8��� �Հ1� ������ �Հ"���U  �΀�Y ����U �� `̀ ]�z�h`H�Z� �� ���� /�L+ϩc�B ��]� ����U� S���� =�� '� 8٩d�B �ȩ�V  2� q��t �u  �� 2� �� ��U ��"� �� �ĩ"��  l� UĜU �� �V �t �u z�h`H�Z Ӯt �u ��^� ����V��� �����g�B  2� q���V ��c�B � S���� =�� '� 8٩d�B �� 2� q��t �u  �� 2� �� ���* �  �� �_ �V �t �u z�h`H�Z��,� ����7��� �Հ0� ������ �Հ!��U  Ѐ�Y ����U �  �̀ ��z�h`H�Z� �� ����� ��L�Щc�B ��]� ����U� S���� =�� '� 8٩d�B �ʩ�V  2� q��t �u  ��� �� 2� �ۭU ��"� �� �ĩ&��  l� UĜU �� �V �t �u z�h`H�Z �Ӯt �u ��^� ����V��� ������V �g�B  2� q��c�B � S���� =�� '� 8٩d�B �� 2� q��t �u  ��� �� 2� �ۀ�* �  �� �_ �V �t �u z�h`H�Z��,� ����8��� ր1� ������ ր"ʩ�U  dр�Y ����U �� �̀ �z�h`H�Z� �� M���� ��L�ѩc�B ��]� ����U� S���� =�� '� 8٩d�B ���V  2� q��t �u  ��� �� 2� �ۭU ��"� �� �ĩ*��  l� UĜU �� �V �t �u z�h`H�Z MԮt �u ��^� ����V��� �����g�B  2� q���V ʩc�B � S���� =�� '� 8٩d�B �� 2� q��t �u  ��� �� 2� �ۀ�* �  �� �_ �V �t �u z�h`�Z��J �t �u �l ��m ���x ���l �m  �ԩ�V ���n ��o ���y ���n �o  �ԩ�V ���p ��q ���z ���p �q  �ԩ�V ���r ��s ���{ �V ���r �s  �ԩ�����J �L��z�`�Z��J �t �u �l ��m ���x ���l �m  �ԩ�V ���n ��o ���y ���n �o  �ԩ�V ���p ��q ���z ���p �q  �ԩ�V ���r ��s ���{ ���r �s  �ԩ�V ����J �L �z�`�Z��J �t �u �l ��m ���x ���l �m  �ԩ�V ���n ��o ���y ���n �o  �ԩ�V ���p ��q ���z ���p �q  �ԩ�V ���r ��s ���{ ���r �s  �ԩ�V ����J �L��z�`�Z��J �t �u �l ��m ���x ���l �m  �ԩ�V ���n ��o ���y ���n �o  �ԩ�V ���p ��q ���z ���p �q  �ԩ�V ���r ��s ���{ ���r �s  �ԩ�V ����J �LZ�z�`H�Z�_ � �
�_ � |�%��
�_ � |���
�_ �( |�	���< |�z�h`H�Z P�H �� I �� z�h`H�Z ��H �� -I �� z�h`�Z ��H �� -I � ����� z�`H�Z��%� S����'� �� p���  2� �� ��� �� �׀
��U �  `�z�h`H�Z��%� S����(� �� p���  2� �� �� �� �׀��U �� `�z�h`H�Z��%� S����'� �� p���  2� �� ��� �� �׀
��U �  ��z�h`H�Z��*�g�B � S����(� �� p���  2� �� ��� �� ؀��U �� ��z�h`H�Z�� �� ��� ������  2� �� ��� �׀� �� lĩ"��  �� U� ��z�h`HZڮ� �� ��� ������  2� �� ��� �׀� �� lĩ��  �� U� ���zh`H�Z�� �� ��� ������  2� �� ��� �׀� �� lĩ&��  �� U� ��z�h`�ZH�� �� ��� ������  2� �� ��� ؀� �� lĩ*��  �� U� ��hz�`H�Z �� l� �� U�z�h`�Z�J �mJ J����� z�`H�Z��W  p�����$��"��  �� l��F �F  U� ��W ��z�h`H�Z��W  p������� ��  �� l��F �F  U� ��W ��z�h`H�Z��W  p�����&��(��  �� l��E  U� � ��W ��z�h`H�Z��W  p�����*��,��  �� l��E  U� � ��W ��z�h`H�Z 2� ���W  p�����B  ���F �F  q� ��W ��z�h`H�Z 2� ���W  p�����B  ���F �F  q� ��W ��z�h`H�Z 2� ���W  p�����B  ���E  q� ��W ��z�h`H�Z 2� ���W  p�����B  ���E  q� ��W ��z�h`H�r�B  R�h`H�p�B  ��h`H�t�B  ��h`H�v�B  ��h`H�Z�� ��e� �W �� � S�����W �0�W ��9� �W ���� �ۜW �� � S�����W �0�W ���W ���� �ݩ |��� �� z�h`H�Z� L��� ��� �" �����j �k � "٩�w L���̠ � ��̠ 0Lr���� �����j �k � ٩�w L�ۈ��� �����j �k � -٩�w L��ʈ� �LM� ����LMڎj �k � ٩�w L����� �L�� ����L�ێj �k ��w � "�L�ۈ� � �����j �k � ٩�w L������ �����j �k � -٩�w L������L�� ����L�ێj �k � ٩�w L����� �����j �k � -٩�w L���̠ L]ۈ� � �����j �k � ٩�w L����� � �����j �k � "٩�w L������L�� ����L�ێj �k � ٩�w L����� �����j �k � ٩�w L�ۈ�� � �����j �k � "٩�w L���� � �����j �k � ٩�w z�h`H�B H�a�B  q�h�B h`�Z�U ����������������� ����O �P z�`H�Z�i �� �� ��w ��L_܎j �k �w � � ��Lbܭw �� ��Lbܭw �� 3�Lbܭw �� {�Lbܭw �� �� �� ��z�h`xH�Z�� �9 ͌ �L9��8�9 � ��ح� � �L9ݩ �� =�� �x �� A��G �l �m �x �` �[ �} ΅ �� � �t�y �� A��G �n �o �y �b �\ �~ ΅ �� � �K�z �� A��G �p �q �z �c �] � ΅ �� � �"�{ �� A��G �r �s �{ �d �� �^ ΅ z�hX`H�Z�l �m �x ���w �[  ލ[ �w �x ����l �m z�h` >� {� �� ��`H�Z�n �o �y ���w �\  ލ\ �w �y ����n �o z�h`H�Z�p �q �z ���w �]  ލ] �w �z ����p �q z�h`H�Z�r �s �{ ���w �^  ލ^ �w �{ ����r �s z�h`�Z�Z ��0� �̠ �� ���w � |��f�B  2� q� J�����Z �Z z�`�Z�O �=0�P �O �P �0���� z�`Hڭ� 
��ʽ���� ����� �h`H�Z� ���� ����� ���� ���8��z�h`H�Z�c�B � Ȣ � ����	 2� q� �������z�h`H�Z� Ȣ � S���� ��������z�h`H�Z�� �4 ����-�j �k � و� �� �0 � 0��� ������w ��� � �w z�h`H�Z��5� ����-�j �k � ��� �� �0 � ��� ������w ��� � �w z�h`H�Z��5� ����-�j �k � "��� �� �0 ̠ ��� ������w �� �w �� z�h`H�Z��5� ����-�j �k � -��� �� �0 ̠ 0��� ������w �� �w �� z�h` �� lĩ �� C� �� ��v � � ��ʎv  ��x ����l �m �[ �y ����n ��o �\ �z ����q ��p �] �{ ����r ��s �^ ��� ��� Lf�H��x ��y ��z ��{ ���; �Y h`H �� �� � �� ��� �� ��LZ�h �� k��  � ̮ ���E ��F �	�H �7�I � ����� �����  g������ ����� �
�E �i�F ��H ��I  g� ����G  ǭ  ���G �� �� �� � �霂 �� �  k�L8� �魞 �� ��  �ĭ� �� �: �; �Y �U h � ��L;�`H�Z�� �� �l ��m ��[ ��1�n ��o ��\ �� �p ��q ��] ���r ��s ��^ �L�z�h`H�Z �© k�
�E �2�F ��H �I �� ����  gÜ�  � ̮��E �d�F � �� �­i ��	�  ������ �� �  k�L8�z�h`xH�Z� �  r����� r���Ȁ� r�� �ʀ� r�� ����z�hX`�Z 2� �� �o�B  q�z�`H�Z�ލ&  ]� d��E ���F ���N � ��  ��� �����i ��E ���F � �� ���ߍ&  T� ��z�h`H�Z�d�B  2� q�z�h`H�Z�l �m �x ��@�n ��o �	����y �p ��q ��z ��	����z �r ��s �	����{ �n �o �y ��&�p ��q �	����z �r ��s �	����{ �p �q �z ���r ��s �	����{ z�h`H�Z�g�B �w �� (�z�� ��q�� ��h�� T�_̠ �5̠ 0�� �Ȁ( S����Ȁ� (�=����� S������� ��%� 0� S����耻� ��� S����ʀ�� T�  z�h`H�Z��P� S����G�j �k  2� �� ��ȩg�B  �؈��w �| �| ͍ 0(�| � ��w �������w �
Ȝw �j �k z�h`H�Z��P� S����G�j �k  2� �� �舩i�B  R�ȩ�w �| �| ͍ 0(�| � ��w �������w �
��w �j �k z�h`H�Z��P� S����G�k �j  2� �� ���k�B  ��ʩ�w �| �| ͍ 0(�| ̠ ��w �������w �
�w �j �k z�h`H�Z��H� S����?�j �k  2� �� ��ʩm�B  ����w �| �| ͍ 0 �| ̠ ��w ���w �
ʜw �j �k z�h`H�Z�a �<0$� �a �� )�
��� )�i�� �`�� �� �"�E �#�F �� )�B  q��"�E �>�F ��  &� i�z�h`H�Z�U �� ��*��x �y �z �{  E殟 ��  �ĩ"��  Uĩ�; �Y z�h`H�Z�a�B � Ȣ � �� � 2� q�������z�h`��� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� � �b�� �� �� ����$�� �� �� `H�� �� �� �� �� �� �� ��� ��v �[ �\ �] �^ �7 �8 �9 �; �Y �: h`�P �a �` �b �e �c �d �f �g �h �w �x �y �z �{ �| �} �~ � �� �t �u �V �X �_ ��l �m �o �p ��n �r ��q �s ��� ��� `�G � �%��Pm� �� �� i �� �� i )�� ��G �� ��`H�Z�� ͝ 0&��� ͜ 0��� ͛ 0�� �� �� �� �� �� �� ͝ 0&��� ͜ 0��� ͛ 0�� �� �� �� �� �� z�h ��`H�Z�0���������  ��z�hL� ��z�h`H�Z����������  ��z�hL�z�h`ʈ��0��I �JJJ�G �
mG �H ��I � �	� 
��I ���I `H�Z P�H �� I �� z�h`ʈ��0��I �JJJ�G �
mG �H ��I � �	� 
��I ���I I��I `H�Z ��H �� -I �� z�h`ʈ��0��I �JJJ�G �
mG �H ��I � �	� 
��I ���I `�Z ��H �� -I � ����� z�`H�Z�
i�E �


i�F z�h`Hڪ�a�




�I ��)I �& �h`H�Z K�
��U��� �U��� � �� �@�� � � ������(���� i0�� �� i �� �� i(�� �� i �� ���Ωߍ& z�h`H�Z�> �@�? � � � �>����? ���z�h`H�Z
����L ���M � �L�$�&H�H ��� ��h�a��b�8�7�B  q��E �E Ȁ�z�h`H�Z�)�JJJJ�B  q��E �E �)�B  q��E �E z�h`� � �  ]� d� � � � � � � � �5 �6 �ߍ& �* `H�Z� ���Q� ���.� � ]� � � �  T� � d� � � �  ��� � �	 � �� � � � �� ���.�( � ]� d�! �" � � � �  ��( �( �# � ��(z�h`� �� ȱ� ȱ�	 ȱ�
 ȱ� )
��?�� �?�� Ȍ � � �	 � �'� �-� ȱ-� � �� � �� ��Ȍ � ��`� ��! ȱ�" ȱ�# ȱ�$ ȱ�% )
��?��& �?��' Ȍ �( �) �# � �#� �  ]� d� � � � � � � � `� �� ȱ� ȱ� ȱ� ȱ� )
��?�� �?�� Ȍ � � � � �'� �/� ȱ/� � �� � �� ��Ȍ � ��`H�Z�
 )?	@�+ �
 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �5 �� �5 z�h`H�Z� )?	@�+ � 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �6 �� �6 z�h`H�Z�$ )?	@�+ �$ 4��-+ �+ �) �&��% )@��J��+ �+ Ȍ) �&����) �% �) �+ � � �5 �6 z�h`� �5 `� �6 `H�Z

�����- ȹ���. ȹ���/ ȹ���0 � �-� �/� ȱ-� �/� � � �� �  � �� T� ���� z�h`H�Z
��)�� �)��  � ��*  �� ��� z�h` �� �� �� ��� �� �� ��� �� �� �� ��    ��� �� �� � � �� �� �� q� �� �� �� �� � � ��    ��� �� �� ��� � �� � �� q � � q� � q� �� �� �� �� � �    � �� � �� �� �� ��� � � � q� q� � q� q� q� d� q� �� � � � �� �� � �� �� ��    �� ��� � � � ��� �� ��� �� � ��� �� q� �    q� _� _� q� �� �� _� q� _� q� �� � � � �� �� ��    � �� �� �� _�  d�  q�  w�  �� _� �� �� �� �� �� ��.� �� � �    �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� q$�    q$� q$� q$� $� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� w$�    �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$� �$�\$��$��v�    �� ��    �� ��    K� %� _�    � �� �� �� �� ��.� ���T�h� ��    �� �� �� �� ��� �� �� ��� �� �� �� ��    �� q� Y� �� �� �� �� �� �� �� �� �� �� �� w� C� ?�    T� q� d� _� K� T� _� �� �� �� �� �� �    d� T� _� q� d� � q� �� ?� T� K� T� K� O� T� d�   ������������.�������\�������.����h���T���@���.�   .����h���T���@���.���\���:����������\�:�    � � � � � � � � � � � � � � � �   �� �� �� �� �� �� �� ��     �� �� �� �	� �� �� �	� �� ��    ��  _�  ��  G�  8�  /�  %�  �  �� �� �    _�  d�  ��  ��  ��  �� � .�  ��  ��  �� ��  ��  ��    �� w� d� K�    � �� �� �� �� �� �� �� �� �� �� ��    ��� �� T�     �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��    �� /2�    �
	�

		�
	 �


�
	 �





	�

		���������#���3����r����  n�n�n�n�n�{�{�  ����  ��  ����"�z��  ��  ��K�v�����)�@����9�  F�I�T�g�o�|�������  aaaENTERaYOURaNAME$PAUSE$aaaaa$abaMOUSE$abaWOODENaBLOCK$abaIRONaaaBLOCK$PRESSaSTARTaKEY$TIME$aaaaMINaaaaSEC$BONUS$aaaaNOaaBONUSa$MUSICaBY$XIAOaLIWEI$PICTUREaBY$BANaYONG$PROGRAMaBY$ZHANGaXIAOMIN$]�p�v�|���������������� � � ����������
dnx� � �  � � � @ @   ��� ��� ���
�
�
 �                         
� ������
�
�
� �   �                       �
�
� ���* � �
�
��"                           
�(���(��
�
�
 ��                          �
�� ���* � �
�
���                          �(�
�


���

�
�
�
��             � �           � �� �( �� �� ��
�
�
                            �� �(�
��* �� ��
�            �             ��� ���
�
����
��

                         ��
�
�
��
���
�"��                          �� �� �(
�
�
�

�
 
�
                         �(
�
��
�
�� �"
�

�
�
                         � �����
���

���
 
                  �       ���*�
 ��
�"� �                           � � �
(� �* �� �
�                          ���
�
�
�"�
(�"��                          �
"
�"
�
�
���
�
                           � �
*
� ������ ���
                     �      �(�
�
�
�� � 
���
 
                �             �*�
"
�
�
�
�( �� �

             �             d������D�|�����$�\������<�t������T��� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p�������� ������������������������������������������������������������������������������������������������������������������      h$�$�$
%@%v%�%�%&N&N&N&���0�p����0�p������ԉ �$�t�č���d�З��ԉ��T�)�	����0�                                                                                                                                                                             R� �v�