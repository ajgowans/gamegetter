  �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��?������  �?  �?  �  �  �          �  �  �  ��  ������� �  �?  �� ����������?�o�>�o�>�o�>���?���?���>,��8,�>8�>0�0  < � ��<    < ��ۀ� << � � �<      �<�� � � <      <�� � <  < � ��Ӏ<��?���������?���:+����l9���:��;�;���:���        �����(� �(�(���*(�((�(��(�����  ��  ������������� �� ���������������(���(�`UU	�VZUU���ZUU��(`UU	( ��� �?  ��   �             �  ���?  �������������������
"�����������"""
    << �  ? ���������������/���������?������������������������������������?�����������������������������?��  >  8�         < <   ���� �?����� ������� ��몪��? ������> ������ �ꮾ�� �믯��� ����?� �����<  ���   �������0�����  ?  �?       �        �                                    �         �      0 �     < �? � ������?�������������������? �  ��?�     ��      ��      ��      ��      ��       ��       ��    � ��  0����?<�����  �   ��  �(>  �� ��A��� Fl`	9^�Uj�����껻�������L      0 00   � 0   �  80  0�  ��  �}  |�=  �}  ��   �    <  �� ��� ��� ���   �?   �   �   �               03333���������������?�������?�������� ���? ��� ��� ��� ���? ���� �������  <��뫪�j9�j8�V8 8 9 p9 �9  ;  , �  �  �  +9 �*� �Z��ZA�jU:���?<  ������lP5����� �: � � �  8   � ����<�<�<�[��[���<�<�<���� � � �? �? �� � �        � � �? �? �� ��� pU  4 )lU�������� ��  ;   ? � � �  �  � � � � �? �? ���������?\}5����<��<��<�<������,<8���� � �                      � �? �   ?  ? �� ����?���� ����������}��}��}��}�����������������������W��������������������������������������W�������������������U��U���UU��_���UU��_�����_���_���UU��_���UU��_����_�_�_��UU��_���UU��_���UU��_�������[nyut mm@����@{     �������|<W �����U���� �_ �����?��ꫪ������Ѓ��� ˃�������? �  ,� ��Hp8����	,� 2�,Έ#b"�Ȍ؈#"�!��16�1K	 ����	 ,�  �   0   ���    !  ��   0 �� ��  !� 0�b @$� 0"��@��0"�H  � # ��#B �0B  #4    �  00   �   0   0 � � 0�0 ?�?�� 믳 뚯 �V� �^E� �j����� �E� oU:  �Z� ���� ����>��� � 0 � �   0  �0�>; ����F� ��? � �f� �^������ 0        ��      ��      �j�      oU�     �U�    �ZU��  �Z���>  ������   ���Z�     �V� ��?�kUU ����kUU:𫪕�ZUU��VUU՚Z��UUU�ji��oUU��V�e�kUU��UUZ�kUU��UUj�[UUo�UUi�[U�[�UUe�[U�VoUUe�kU�UoUUU�U�UoUUU�U�UoUU���V�UoUU���k�UmUU�>���U��U�? ��V���� _�Zտ�� _�_U��  U�Z��  �U���5  �UU��5  �WU�p  �U� �   ��     �     V	 ��  V%�oU X	�VU ��UU9 ���UU9 �jiUU9 �U�UU� [U�VU��WU��U��VUY�V�UU[UU�kUU[UU�kUUkUU>kUU���[UU���[�WU�� ��WU�? ��_�� ����   ���   �Z9    ��     �    �?   ��   |��  ����_iU?�UZU�_UVU�WUUU�WUUU�[UUU��U]�?�V}�>��� o��  �V?  ��  ��V��U�[U�WU�WU�oU=�[ �  �?  �� �����|l�9\�~5`�_	��� �?  W� �UUpP\@5|UU?������������lQ\@k@:[@9kQ:��:lf��pU��������`Y�� �� �� �� �� pj��pU��       ��3s53��w����W �WU5\U��kU:��?��  pw |w ww�wwsww�GD� � W � W@5 \U �� kU: ��? �?  ��  �� �� �U �� �������_? ��? p�? ��? �� ��  �   �  �� �� ��? p�? ��?��_?������� �V �� �� ��  �?   �0 ��;������������@UU������:�����������3��� ��  �� ���@UU������:�����������3��� ��  ��  �  ?�??�?�>����������V��[�  �:  �?  �  �   0<� �?<   �   �  �  �> ��� ��� ��� �V��[��:?�???�? �      < ��    �  ��  �; ��. �? ��? ��?��������� �? � ��    �?  ��  �� �� ��? ��� ����^ �� �� ��? ����� ���<�<0����  �> �z� ��0�9��� ��� ��� ��  9 ��� ����� ��<��<.��������?��3ln����������?< �  �/  �� ��������?�������?���������:���:뺺����3�  �  �/  �� ���������?�������?���������?���;�������� ��?�� ��,8000080������  <  �  �  �  �  �  �  � ���08,088,0������  ??  �  �  ,    8  0  ??  �?  �  �  � ��� ���������?���?����������_�������  ??  �?  �  �  �  �; ��� ������������������_������� ?�� � �  �  �  �       � � � �� �? � � � �          �  ��0��? ��?  �?  �?  �?  �?  �  �  �          �  ��  �?  �?  �  �  �          �  ��  ��?������ �3  3  3    ?  � �������� �? � � �  ?  ?  ?      ��� �� � � � �    ?  �  � � �������������� �?      ?  ?  ?  ?  � �?0������������? � � �  �  � � � � � �3 ��������  �?  �  �  �      ������� �����������?  �  �  �   �   �  �  �  �  �  ������ ������������ ��?  �  �  �  �  �  �  �  �  �    �       ��?     ���  � ���� � ��� �� ����? �� ���� �c�o��V���c�Z��V�ɣ�Z��Z�_ʌ�Z�몥_2�֪�����2�֪�����2��� ���2�ֿ�����p������Wp��UUU�_�UUUUU� l�ZU��9  lUiUiU9  l��Z�9  ��UUU�;  lU�U�9  lU��VU9  �U��~U:  ������:  �jUUU�:  �jVU��  �j�Uj�   k��Z9    ���V?    ��     WU�      ��>      ��   @ PP\|�������������<�?33�/8��  ��
�
�
�)�)�)h�n�o�o�o����?��    ��    ��    �>�    p:k1���?L�[���������W�?���WUU���ܯVii��7� Xj�% ?�����
��������?�����:\�?�*�Z5������?������?ܟ�����7\�V����5p�V�_�����꫖V���UU���Ze]uY��Ze}}Y� k���Z�  l���W9  ��UU�?  �V����  ������  ������  :�[�?�  
���  ���    [�      l9      �   �������������������������������������������������������������      ?�    �7������6������6\�:���5L����1L��ðo1���o00}*��}0]�ڧVu�_U�VU��ZUUUU��Z  T��j��T��j��
R�𪅠
R�𪊪�������������ꫪ�����k�����z������_������W�����ץZ����W�j�� �W�j��  �W�j�:  �����:  �����  �����   ���                   � 

(���(����d���d $� ��  d�  �   �X   �X  %`U @	�UU ZE�  ��       
    &   $(  �� ���X��Eb��aAb� FAb�@b�
@I�
Z@e��V@U�VU U�V P�V P	X P`U@� �VQ*  ��  HHHHHHHHHHHHHHHHHEFFFGHHHIZ++JHHHI+ZZJHHHI+Z,JHHHIZ0,JHHHI,ZZJHHHIZZ*JHHHKMMMLHHHHHHHHHHHHEFFFGHHHIZZZJHHHI--,JHHHI/-,JHHHI---JHHHI-.-JHHHI,-ZJHHHKMMMLHHHHHHHHHHEFFFFGHHI+,,+JHHIZ++ZJHHIZ,,ZJHHI+Z)+JHHI,0Z,JHHI+,,+JHHKMZZMLHHHHIJHHHHEFZ,FGHHI,ZZ+JHHIZ-Z+JHHI-.-ZJHHIZ-.-JHHIZZ-ZJHHI*ZZ,JHHKM,,MLHHHHIJHHHFFFZZFFFZ,,ZZ,,Z+ZZ++ZZ+ZZ,ZZ,Z+++,ZZZZZZZ,ZZ+0,Z)ZZZ,ZZ0Z+,ZZ/ZZ,+ZZ+Z,MMMZ+MMMHHHIJHHHHHE+ZGHHHHIZ,JHHHHI,ZJHHHHI//JHHHHKMMLHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHHH�TTTTTTTTTTTTTTTTFFFFNTTTZZ7ZOTTTZ3ZZJTTT7Z43JTTTZZZZJTTTZZ6ZJTTT34ZZJTTT3Z77JTTTMMMMSTTTTTTTTTTTTTTQFFFFTTTP3ZZZTTTI791ZTTTIZZ77TTTI3ZZZTTTIZ8Z5TTTI3ZZZTTTIZ732TTTRMMMMTTTTTTTTFFNTTQFFZ7OTTPZZZZJTTIZ7Z9JTTI3Z7ZJTTIZ4Z5JTTI6ZZ3JTTIZ4Z7JTTI7Z3ZSTTRZ3ZJTTTTI33JTTTTIZZ7FNTTRMZ7ZOTTTT4Z3ZFNTTZZ37ZOTT37ZZ6JTTZZZ8ZJTTZ2ZZ4JTTRMZ77JTTTTRZZSTTTTTIJTTTTTTIJTTTTQFZZFNTTPZ37ZOTTIZZ3ZZFTI34ZZ6ZTI3Z6Z81TIZ4Z5ZZTI7Z7Z3ZTRZ3Z2ZMTTRZZZSTTTTKMLTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTTT�YYYYYYYYYYYYYYYYYYYVFFUYYYYPZ<OYYYYI<CJYYYYIZDJYYYYIAAJYYYYWMMXYYYYYYYYYYVFFUYYYYPZZOYYYYI==JYYYYIBBJYYYYI>?JYYYYWMMXYYYYYYYYYYYYYVFFUYYYYPZ@OYYYYICZJYYYYI;AJYYYYIZ;JYYYYW@CXYYYYYWJYYYYYYVZFUYYYYPZBOYYYYIBZJYYYYICDJYYYYIDZJYYYYW<<XYYYYYIXYYYYVFZUYYYYPZ@OYYYYIACJYYYYIC:JYYYYI@AJYYYYW@ZXYYYYYIJYYYYVFZZFUYYPBZZBOYYIZ==ZJYYIZ>?ZJYYI<ZZ<JYYI<ZAZJYYIZ@Z:JYYWMZ@MXYYYYIJYYYYYE<ZGYYYYIZ<JYYYYI<ZJYYYYKMMLYYYYYYYYYYYVUYYVUYYPOYYPOYYIZFFZJYFZZZZ@ZFZZ@ZZZZZZZZ>?ZZZZZBZZBZZZB=ZZ=BZZ<>?>?<ZAZZZCZZAZZ<ZZ<ZZMXW<<XWMYYYWXYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYYY�	
##''++,,11 !
"d��������������	!%++,,//666  '## R������������ &&))016677889999:?? " (
#(((^����������������      )*(+-4(0*0'0#.*F&($2$&$,(&(+)+'P

		


          $(&*$+$-&'$'%"&C(&''+&'+%)$)$+*P




				

         "&%"""!"Q








                                                                                                                                                    �������������������������kjjjj����������                                                            �������������������������jjjjj����������    �    �    �    �    �    �    �    �    �    �    �    ����������ꪪ��ꦦ��檪���jjjj�����������PUUU     UUU@ PP Q@AEEU@QPTU UUA AUUA AUU UPTEU@QQ@AEP  PUUU@     PUUU                                                                                    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    ������                                                                            �����    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    ������                                                                                                  ��  ��>  ��  ��  �� �j~@ ��P ��T ��T��~T��_ P��P k� TA�> UA� UA�P@� U U_P S      �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �   ��   ��   ��                                                            ;    �    �   �   �:   o�   ��  ��  ��:   ��  �� � �k: �� A��@��@ԫ: �� ��  �� �� U�@U�PP �P  �U  �UT1@T PU P� @5     T �  A5  @  @  �   4         �    0            W   \T0@T�PU SU LU@ 0  P �T T  WT  \T  p P  �P    WA   \A   pA   �@            0    �U   UT@T PU PU@U@   P T TUTAUT@U P@P  TA UA  UA P@ U @UPP P     ��  ��>  ��  ��W  ��T �j~ ��_  ��W ��U��~ @��  ��C k�PQ �>P@�_ A�W P�UPUP T P    o�   ��  �  ��:  @��  P�� P�� �k:  ��   ��T�U��:P��DP�� P �� T ��@U�TPU�  T �    �    � @ 0 T  EP@U� P 0 P  P  �    4  T  U  �   D0           �    4                @  0T �EPU WPT  P 0 T  �T  U  \ @  0    �    S    L   p   �        \    p    �      @   T  EPU@UPTP PP T PT U  T @T   U@ PQ DP@ P A T P@UTPUP  T P                                                   ?   �U�  \UU |U����; ���� �������� ��� ��         0   ��  ��>  ��: ���:���;�k�;�;����;����:����:���������꼪��������ګ��j���������뗾�?��?                           �    �   [  �[�  �n� �j� �f� ���  ���  �:   s   p  �  ��  ���                       �    �   �  �j  ��
  �k/  (�*  ���  �n
  �k
  ��+  *l�   l   �o   ��  �                          �*@ @��B  �j
 �& ��* ��)  ��� ��         �  HP                                               �   ��  ��
  ��*  ��  p�  |U  |}  �}  ��   �?                                       3  ��  pU:  �>  ��  ��  ��  �{  ��  �{  ��  ��  PU                       0  ��?  ��� �������/��������
8������U� ��������U���UU=��WU���_Uu���Wu������  ��?                                         �?   �5   �?   �?   ��   �� ��  ��� ��� � ��� ��� �?    �   ��  ���  ��� ����������-�Z�5��Z�6��j�:�zj����j�ڬꪭ�ꫵ�������������V���������������+  
�   (*  ��� ���
 ���* ���+ ���. ��( :��  �   �
   �   �
   �   �
   �   �
  "� ����
 ���                 @
   @
   �*   ��   ��  ��
 @��* ���* PUU%  ��  ��  �  � �� ��� ��  ��                 z
  �~
  ��*  ���  駪@���
�~��*T���*�ZUU%�ꧯ�j��j��j��j��_�����_U�?   �<   ��  �� ���? ���> ���: 쯯� � 믪� ���� ���: ��� ���  �  �_  �_  �_ ��_ ��} ��?  ( �  � (  �
.  �*+* 諫
 ������
����
���*+����,����   ��   �   �   �   �  �  �  �
  �(              (    �   ��  ��
 P��* ���. ��� ��:���:������ � 0. ��
 ���
���� �*�           �            �    �
   ��  ��j �i�	 jj�*��j�����������? ��?3 ��   �   �  ��  ��  ��  �?                       �   |��  WU�  �_�  ���  ���  ��.  ��.  ��>  ��>  ��: ���? ��� ��  �                                      ?   ��   �  ��  ��: ���� ������������:���������*������
 ��+         @   �=   ��   p�   ��   ��   ��   �  {u  �~. ���: ��� ���  ��  �>  �       �� ���                  �    �  ���  ��� ��W �zu �j�	 ��U ��w ��^ ���   �>  ��  ��  �?                                ���� WUUU ���� WUU� ���� ���� ���� �U�� |U�� |U�鰻���������@AAA� � @AA��    �   �   l   ���� �{U� ���� V�U� V�� V�� ���� ��� ���% ��ک ��ڻ����.�����PP �� ��P    �   p  0� �p; �p; �p; l�= l�z9 �k� ��  �   p   p   p   p <�  �p � ��   �                                       ( �  � (  �
.  �*+* 諫
 �������
����
��?+��,�CUE  TAP                �   �7   �V   �� ��u ��W �z] ��U �ju ��� ��W  �U ��   �^  ��> �� ��  �?                 �  �   (    ,  �                  �   �/    /   �/   �
   ,         (                                ��<  |U� |�� ��< ��� ��� ��� �j� ��p ��p���p����  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��?������  �?  �?  �  �  �          �  �  �  ��  ������� �  �?  �� ����������?�o�>�o�>�o�>���?���?���>,��8,�>8�>0�0  < � ��<    < ��ۀ� << � � �<      �<�� � � <      <�� � <  < � ��Ӏ<��?���������?���:+����l9���:��;�;���:���        �����(� �(�(���*(�((�(��(�����  ��  ������������� �� ���������������(���(�`UU	�VZUU���ZUU��(`UU	( ��� �?  ��   �             �  ���?  �������������������
"�����������"""
    << �  ? ���������������/���������?������������������������������������?�����������������������������?��  >  8�         < <   ���� �?����� ������� ��몪��? ������> ������ �ꮾ�� �믯��� ����?� �����<  ���   �������0�����  ?  �?       �        �                                    �         �      0 �     < �? � ������?�������������������? �  ��?�     ��      ��      ��      ��      ��       ��       ��    � ��  0����?<�����  �   ��  �(>  �� ��A��� Fl`	9^�Uj�����껻�������L      0 00   � 0   �  80  0�  ��  �}  |�=  �}  ��   �    <  �� ��� ��� ���   �?   �   �   �               03333���������������?�������?�������� ���? ��� ��� ��� ���? ���� �������  <��뫪�j9�j8�V8 8 9 p9 �9  ;  , �  �  �  +9 �*� �Z��ZA�jU:���?<  ������lP5����� �: � � �  8   � ����<�<�<�[��[���<�<�<���� � � �? �? �� � �        � � �? �? �� ��� pU  4 )lU�������� ��  ;   ? � � �  �  � � � � �? �? ���������?\}5����<��<��<�<������,<8���� � �                      � �? �   ?  ? �� ����?���� ����������}��}��}��}�����������������������W��������������������������������������W�������������������U��U���UU��_���UU��_�����_���_���UU��_���UU��_����_�_�_��UU��_���UU��_���UU��_�������[nyut mm@����@{     �������|<W �����U���� �_ �����?��ꫪ������Ѓ��� ˃�������? �  ,� ��Hp8����	,� 2�,Έ#b"�Ȍ؈#"�!��16�1K	 ����	 ,�  �   0   ���    !  ��   0 �� ��  !� 0�b @$� 0"��@��0"�H  � # ��#B �0B  #4    �  00   �   0   0 � � 0�0 ?�?�� 믳 뚯 �V� �^E� �j����� �E� oU:  �Z� ���� ����>��� � 0 � �   0  �0�>; ����F� ��? � �f� �^������ 0        ��      ��      �j�      oU�     �U�    �ZU��  �Z���>  ������   ���Z�     �V� ��?�kUU ����kUU:𫪕�ZUU��VUU՚Z��UUU�ji��oUU��V�e�kUU��UUZ�kUU��UUj�[UUo�UUi�[U�[�UUe�[U�VoUUe�kU�UoUUU�U�UoUUU�U�UoUU���V�UoUU���k�UmUU�>���U��U�? ��V���� _�Zտ�� _�_U��  U�Z��  �U���5  �UU��5  �WU�p  �U� �   ��     �     V	 ��  V%�oU X	�VU ��UU9 ���UU9 �jiUU9 �U�UU� [U�VU��WU��U��VUY�V�UU[UU�kUU[UU�kUUkUU>kUU���[UU���[�WU�� ��WU�? ��_�� ����   ���   �Z9    ��     �    �?   ��   |��  ����_iU?�UZU�_UVU�WUUU�WUUU�[UUU��U]�?�V}�>��� o��  �V?  ��  ��V��U�[U�WU�WU�oU=�[ �  �   �  ,  8 �j� �Z��jU���: �   �   �   �   �   �   �   0  � ���,l��	�2�6�:�8�0� � 0 ��?���[U� ��U�WU�W}�WU�WU�������\U5pU����?���[U� ����WU�W}�wU����� ����\U5pU�� 0  �  ��#�">�!9�!�l �l!�e��f>����     � < � < � � l� ,�/����\�� |�� ��= �� �  ���+ :�  �  �� ���UU:lUU9[��[�7�l�C9lUU9��Z��W�V� [�  l9  �  � ���:����������UU:lUU9[��[���l�C9lUU9����_�֗ [�  l9  �  �  ��  ��  ��    ;  ����?�U�=o��U>����������  ��  ��  ��  ��  ��   ��    ?    ?      ������  ; ��U?��5��:��:������������ ��  ?  ?    �  �� �j��V���[:l}y9k��[W��[W��k��l}}9��[:�V��j� ��  �  < ����U>l=9_��ۢ�ۆ�ۆ�ۚ�o��=9�V>��� <    �   �   �  �?  �� � �? |� o� ��  �� �[ ��? ��  �  �  ?   �   �   �  �   ?  �� ��? �?�  O> �� �� |� �> �         ??? ���� �!?�����  /?>  ��  ��: ���� ���,��*���9����8,B ��՛�3�  ��   0    <?��,?��0?��.��8��2��:��:��8��8o>�� 3 �� 0  �   � �� �� �<? p<����?���������������?�_U ��  00 �?0   0�  �  ?  ��  �� �� �<��<���?���������������?�U� �    �?  �   �  �  [9 ��� �V� ��� �V� 0�?0[9�z�  �> ��� 0��<��<��  ? �� ����lU��lU��3��3������.��<��<�� ������_}�_}�_��_��_�����������_��_��_��_}�_}���������������_�W�_�_�_�����������_���_�_�_�W����������������������?���  �  �  �  �          �  �  �  �?  ��  ������� ��? �����                  ?   � �� �� �� ��? �� �? ���� �  �  �  �  � � � � � �? �����  �?  �  �  �  �                  �  �  �?  ��  ����? � � � �                   � � �����������?��0    ? ��� �� ����?������?��? �� �? � � ����������?   �   �?   ��  ��� ���  ��?   �   �   �    �    �   �   ������� � � � �  �  �  �  �  �  �  �  � ���� �? �? � �               ?  ����? � � � ?                 ����� �?  ?  ?  ?      ?  ���? � � � � � �  �  � ������� � � � � � � � � � � � � ���������  �  �  �  �  �  �  �  �   �     ��?   ��  �  ��  �� ��_�����_����zUUUU��V�����h)��*���*����*�� ��*��  ������  ������   � �  _U�_U�  �Y�_e�  _f�_��  �Y��e�  l���V9  l���V9  �����:  ��曦>  ��曪>  ���[�?  ��[�  ��_�  ��_�  ���߯  �����  �����   ����    ���?    ���     �:      �?      �   U}}}}}}}}}}}}}}}}UU}}}}}}}}}}}}}}}}U    <    �?  �  ��� �A W>�UpA����Zp��� [����  [������ �[�������[������|[������=��������kW��U����k��zU����k�UzU�Uk��UzU�U�:��UzU�U�? �UnU�U�  ��kU��  ��U��  �
U��   U��    �U�?    �U�    �U�    �U��   ��^U��  ��ު��  ��� ��   �>ü�    �?���    �?U��   ��{��  ����  �:����  ���    ��      �U   0<0333333????���    * �� �� �� �� �� �� �� �� ����/?>?<<< <? ? 0    <        <        �       ��      ��     ��A�    ��A�>    ��U��   �j��~� <�V���:<<lU��U9<�oկ��W���j���
����_�������V � �����V�P�����U�PU�?���/ �_�?��}u ]}�?��wA�� �=w��|:  �����:  �U��ZU:  �U) hU:  �V����>  �V����  ������  ������   �����    ��(��    �[U�    �+��     ���      ��>      ��   UUUU���������UUUU       ������������������������������������������������                                                                                 	    	     
                    	    	
	
   
          
   	                  	
                	 	
 
         
    	     	             	  	   	                                                                  �                
   !   !!   !   !  !     !  !	!  !!
  !  !   !   !      	 ! !
!              !	        
   ! !  !   	  !	
!  
!      ! ! 	 !                         ! ! !	!  !!   	 !! 	 ! 	 	


 !! 	 !	 !! 
!    !      !	!	 		  	                                                                  �          
  
''   '      ' '    % '
 %&$ '  '   ''''  %$  (((((((( %    %%##"##"##''    %'' '  %&' $    ' ''   '% '	 '  '%	'$ 	 	
       
% $  ' '	 '$ '    '   ''   '        '   %&'  %%%     	 ''     '$ '     (((   % %% '#"#"##"#'    '      '' %     %'    '%     '  $     $  '  ''  ''  ' '    '%  '	'  '   %%   ' '$'	    	                                                                      �""#'**+000 
#"

#0���������������""#%(,225 '
$
$
_����������$$**++..23 



`L������������������       452<43637345463F534635345365363P



				



        030204130803142A14.128041403192P





				



        +2,1.1/01/80+12J+-.1+006.0-02.,P




				
                                                                                                     T)  @T9   T9  @T�   P�  Q�   P�  Q� @P�  P�  A� @�  D�  @� @P�  P�  P�  U�   U9   U>   T=  U9   T9  @T�   T�  @P�   Q�   P�   Q�   T-  P=   T9  @T9   T�   T�  @T�   T9  @T9   T9   T9    l   l  l   [  [E   [ �Z  �VE  �V  �VA �V  �VA �Z   [E   [   [  [   lU  l   l   |   l  l   �U  �U   lU  o   k  o  lU   �U  �U   �U  l  l  �   �U  lU   l  l  T9  @T9   @9  T�   Q�  A�  UU�  UU�  U�?  ��  ��
  �                                                       D@  UUUUUUUUUUUUUUU�Vi�V������Ͽ� ��                                          �U  h   [ �[ �VA  �VU �@U �UTU �UUU �U�� �Z��  ��   �                                    U>  @�  P�  T�  @�   U�   U>   �   �   �    ?                                                                                                  �    �   �>   U�   U�  D�  A�  U  U>  U>    l  l  l  �U   �V  �ZE  �oU   �U   �V   ��    �                                                                                              �    �   �[   �V   oU   [U  �[  �V  �U  l  lU                          @ P   DT   @T  @@U @ A�  P�   U> D@U> @�? T� T�  @�?  P� U�  T9                        A U   U UU   �U@ �Z  �k   oE  �  �@  �V@ �V �[   o  l   l   | �oE  �[  �[ �V �� �k  �VA �UE  jU   U  U  U   UD                         T9  @T9  T�   U�  T��  AU�  T� T�?  U>  DT�   Q�   AU  DU    U    P                                                                  ?�����믾���j�UUUUUUUUUUUUPQEP@@  @ E                            �    ,  �  �  �?  ���  �
�  �J�   3<   <   0  �?#  �?  �                       �    �   �   �.  �+-  �:3  �2�  ���  ���  ��   +4   �<  �* T?   0  �3  �?#  ��S  �                                           �   W�  �j=@�_� �yu� �zj� �z�= ������ P@UU  P                �� �WU �UU5 ���? �  ��� �� �� �� ��� �*P     UU     T  P                                           �   |1   _�  �� �� ��0 �:8 �8 ���  ��0  �� ��                   �   �+   �    K    K    K    K   �K �{K �_K< ���5 ��� ��5��@5�WUU=�_���������� ��        ��?   � ���7 �70 7���7���70 P7 �S7<�_70 P7< Q�0 P<� 0@P< P0 P�<33  ��� 033         �    �    �4�:������/lA�9k �1���1l��,l��l�_o�  ��   �                             ;   �2   ��   �  �
  �
  �
  �

 �
�" �*����* ��*(���* <�������� |���� ��?                          ��  WU ���;  �0 ��� ���                                                                        �    �  � 0  �;  ��5  �U5  �e�  ���  ��� �����������:����:����������?�                       �  �g�  �b � �f@ �� �j ��� �ǳ ��  �    �0 ����       PU                   �    p   �   �?  ��@  �@ \@ �? ��   �   \   �?  ��   �  �� ��@ ��                                   �  ��9  _�  �   03   03   p7   ��  ���  ��  ��                                                �   �   �   �   �   l�   l�   l�  ���  ���  ��+                      0   ���  ���3 ��� �u�  �U�  ���  ��� (  
 � (`	
 �
 (  
    833���?�833�833�                          �    �   l   k9   k1  �Z�  ��  �Z� �V� �Z�   �;   �  �  ��  �                                     0 �  ���  ઺  �f� ��� � �;��?���U��{�U��U�U�P ��� frU՘���?�                                                                 ������������UUUUUT P ����������                               p�� �i�9 ���? pww7 pww7 ���. �   ��� �� ��� ���       �
   �                      �   p   �5  ��  �u   w  0�=  ��7 W5�  �0  �5   ��   �?�   �  Q�                                 �  �U=  ��7  ��  p]�  q��  �u�  �w���w� p�w� ��� �����    E�   HU        ?   ��   ��  �&  �( ���� �o  {� ��� ���:  |�  ��* ����  3<  �3  ��; ��? ��                                                                  
0 ��/������W��W�U{UUUU}UUUAUUUU UTU P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                ��33030�3�  �� ��� �� �       ���          �?�?      STAGE$CLEARED$BONUS$ENTER$GAMEaaOVER$SCORE$CONTINUE$PUSHaSTARTaBUTTON$CREDIT$RECORDaBOARD$ENTERaNAME$��������������Ăւ݂EKQ�!�,�5�<�E�K�W�e�PROGRAMMER$HUANGaYI$DRAWER$ZHANGaLI$MUSIC$XIAOaLIaWEI$bBONaTREASURE$COPYRIGHT$!#PdxEKQY�Z�\���^	_@_<��^_X_S���^._o_i���_`�`���_&`�`� �_F`�`?�? �_f`�`_�_ ��� � � � � � � � � � �( �) �* `� � � �  � �� � � � � � � � �* �G �O � ���H �S `�����`��������������������`���`�N ���������������
�i�k��l��m�	�������
���c�5� �:�?�d�4�6��9�;��>�@�e�7��<�	�A�f�8��=��B�p�q��x��y�z��{�|� �}�����������1� ����,�������2�� �����������
�������������
��������ʊ
��}��h ����j ����l ����n ����p ����r �Ń�t �у�v �}� P�i ��� P�k ��� P�m ��� P�o ��� P�q ��� P�s �Ń P�u �у P�w ��D�C`H �� �ĩ�X �F�Y � ����X �Z�Y �  ����X �Z�Y ��f  �� �� �� �� �� ��h`H��X �2�Y �  ��� �X �2�Y ��f  ���X �A�Y � ����X �Z�Y � �� ȩ�X �Z�Y �D�f  ��C ��  ��C��D�3�D���C�
�8�C��C�i��i �ة�M  {� �Ā� �� �� �� ��h`H� �ǩ�X �P�Y � ����X �d�Y � ����X �� �������M  {��( ����� �� ���h`H�Z� �  � ���_0P���^0F�
��]0<�:��\0P���[0F���Z0<��Y0J���X0@���W06��L 
� *� J��^� �E������`�- p��^� �Q������`� 
� ]��^� �K������` ��z�h`�Z�]�[�^�\�_� �K�Q����`�W�Z�X�[�Y�\� �E�K����`��W��X��Y`��Z��[��\`��]��^��_`H�Z�`� �Lɉ�(�Y ��X �	 �����Y ��X � �� ͉ ����t��Y � �'�f  �ĭf H�a�f �o��X  ��h�f ��a�  ���' ��a��o��X  ���a�  ���
 ��a�������M  {��f �'� ��Ld��
�f Ld������M  {��f �'� ��Ld��#�f Ld���"��M  {� �� P��e P��o��X  �� �L���$��M  {� {��o��X  ��� ��� {� ��L���L {���M  {��o��X  ������� {� ��Lz�h`��X �P�Y �
 ����X �d�Y � ����X �x�Y � ��`��X �P�Y �Y ��X ��W ���X �d�Y �\ ��[ ��Z ���X �x�Y �_ ��^ ��] ��`Z�
��w��T ȹw��U ���f �'�i7��^�Tz �� �`Z�`��
��w��T ȹw��U ���T�^�8�7��'�f z`H�Z8�7�\ �f �\ ��f ��'�f h`H�A8�7�\ �f �\ ��f ��'�f h`HڜW�X�Y�Z�[�\�]�^�_� �^�E�K�Q����$�E�K�Q�h`�Z�P��������z�`�Z �ǩ�X �P�Y � ����X ���Y � ���	�f � �X �P�Y  ���  )�� �����ީ �P����X ���Y � ���'�X ���f  ���M  {���'�X ���Y �J����f ��a�f  �� ����ܩ� �� ��z�`H�Z� �d�$��a��b��c��d�8�7�f  ��Ȁ�z�h`H�
�����d ����e  ϋ�h`H�Z���c  �� �� �f��h��g��b���c�c�Y �b�X  ��c�|� ���c��t�d���e�c�c�Y �b�X � �f��g ��e�e�e�Y �d�X ��g��f ��e�N� ��L`� �� ���c�Y ��g�b�X � �f ���bi�b�X  ��d�X ��f ���d8��d�X  ��d�d� ��L�� |� �򩀍M  {��d ���� ��z�h`H�Z�f
��ɍ�T �ɍ�U ��8�Y �g��g�Z �h�[ �Y �\ �Y �D�V ���W �X JJ��T-c �V�T i�T �U i �U �[ �[ � �Ȁ��Z �Z � ��\ �h�[ �LQ�z�h`H� �c  ����c h`H�Z�/���� ���� ��z�h`͍�� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              H���T ���U �	�Z �] ��[ ��X �
�Y  �h`H��X �
�Y � �f �(�Z ��[  a�h`�         �?�������<<��� ��<<�� �?�?����� <<�� � <<��� ��?<�����H�Z �� �ǩ �` ��X �[�Y �  � ��X ���Y � ����X ���Y � ���"�X ���Y � � ���a ���b ��X �Y � �Z �7�[ � �f  a� ��X �a .�[ ma �[ � 8�a �i�  �mT �T �U i �U � �Y ��Y  �a ��a � �$�X �b .�[ mb �[ � 8�b �i� �mT �T �U i �U � �Y ��Y  �b �7�b �b �` � � ��L����X ���Y ���f ��Z �[  a��X �` � � �ĭX ��֩��Y ���f ��Z �[  a�` � � �ĭY 8��Y ��ة�X ��Y ���f ��Z �[  a��X �` � � �ĭX �)�֩�Y ��f ��Z �[  a�` � � �ĭY ɍ�ީ(�X ���Y ���f ��Z �[  a��X �` � � �ĭX ��֩�a ��X �-�Y � �a �Z  ��a �] ��a �` �� � �ĀЩ�a ��X �E�Y � �a �Z  ��a �] ��a �` �� � �Ā� �� �ĩ ���P�  �� ��������� �� ��z�h`�  �����` `HZ��$��Z �] �*��[ �
����T ȹ� P�U zh`0���򙖛&��" 1    ��*                               ���                              ���
                              �������                          ��������                         ��������
                         ��������
                         ��ꫪ����            ��           ���������           �       UU�������ꪪZUUUUUUUUUUU��VUUUUUUUUU��
�������ZUUUUUUUUUUU��VUUUUUUUUU��
�*�����ZUUUUUUUUUUU��VUUUUUUUUU��
�
���
�ZUUUUUU��jUU��VUUUUUUUUU��
 ����ZUUUUUU���VUU@UUUUUUUUUU���  ��  �ZU��UU����jUUUUUUUUUUUUUU�� �� ��V���ZU�����VUUUUUUUUUUUUU�� ����V���jU�����VUUUUUUUUUUUUU�� ���jU����V�����ZUUUUUUUUUUUUU�� ���j�����������jUUUUUUUUUUUUUU� UU�V�����������jUUUUUUUUUUUUUU� UUPU������������UUUUUUUUUUUUUUU TUPU������������VUUUUUUUUUUUUUU TUUUU������������VUUUUUUUUUUUUUU  TUUUU������������VUUUUUUUUUUUUUUUUUUUUU������������VUUUUUUUUUUUUUUUUUUUUU������������VUUUUUUUUUUUUUUUUUUUUU���
��*��
��VUUUUUUUUUUUUUUUUUUUUU����* �
��VUUUUUUUUUUUUUUUUUUUUU�� ��* ���VUUUUUUUUUUUUUUUUUUUUU�  ��* ���VUUUUUUUUUUUUUUUUUUUUU�  ��* � ��UUUUUUUUUUUUUUUUUUUUUU�
  ���  ��UUUUUUUUUUUUUUUUUUUUUU�* ����  ��UUUUUUUUUUUUUUUUUUUUUU�* ����*  �jUUUUUUUUUUUUUUUUUUUUUU�* ����*  �jUUUUUUUUUUUUUUUUUUUUUUU) ����*  �UUUUUUUUUUUUUUUUUUUUUUUU% ��UU  UUUUUUUUUUUUUUUUUUUUUUUUU @UUU  UUUUUUUUUUUUUUUUUUUUUUUUU @UUU  UUUUUUUUUUUUUUUUUUUUUUUUU @UUU  UUUUUUUUUUUUUUUUUUUUUUUUU @UUU  UUUUUUUUUUUUUUUUUUUUUUUUU @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU <����?0<0<< <?<?  �������� � � � < �  �  ���� � � ��?  � ������:��oU���: ��[k�l9���nU��9 �� [[Ul9��í��l:l9 �����VUl9�����?l9l9 l9��ÖZ[9��p�  l9[9 l9����o[���p:  ��[ [��p�oW�p9l���� [�o�p>l�V�l9�V��� �_n9llÖ�o9�V���� ��[9l\Ö[[۪� {9 ���[��Öo[���  _ �9 [���WÖ   [ �9���������   �� p�� ��9p9����   ��  l�� [jl=����? �9  ��9 [�l��[U9 p9  ��9 [� l�6�[U: p  � � �> ��:��� �  < � � � ���� �     ���  ���? ���  �z� ���:𯪪C  [����VU9�nU�� �Z�[��VU>lmU�  �V[�֪�l���  ��[����l��?  ��[��  k9    �����  [>    �寖��   [    ��Z���  ��    l�V� l�������?  l�V�loU���VU:  k�j�k[U鰶U�  [��U[�������  [>�U[��?���� �Z���Z  ��    �V��Ö  l�    ����Ö  l9    ��|���  [:    ��_9����?���� ���>����:۫�� l����UU�ZU�  l�U� �nU��VU�  ��� �����>  ���   ��� ���     �������                      ��oUUUUU�>  ��������?           �UUUUUUUU� �_UUUUUUU�    ���  �_UUUUUUUU� _UUUUUUUU�� ����� �ZUUUUUU����WUUUUUUUUU�?��UUU�> �ZUUUUUU��oUUUUUUUUUUU�?WUUUUU�������VU�jUUUUUUUUUUU��UUUUUUU ��������ZUUUUUUUUUUUU��UUUUUU�> ��������VUUUUUUUUUUUU��UUUUU��?      ���VUUUUUUUUUUUU���������        �����jUUUUUUUU���������        ��������jUUU���� ������     ������������������   ��?     ��ZUU���������������          𿪪��U� ������������           𪪪����                        �������?                  ��?                            �_U�                       �����_U��                       pUUUUUU��                       ��������?                       �������� �� ��hU
XU	ZU)VU%VU%��*  ��  *    9 @� �Z     H�Z������� �	�������(�
�������?�� ������i�����i���!�b �` ��a  �Ǣ �� 塽��X �	�Y ��8�Y �[ ��[  ����a ���b �b ����a �b �(�<�!�7� 塭��X ��Y  a�!�������(��!��������!�b ɂ���a �b ɖ�~�` ���X �i�Y � ����X �v�Y � ���b ���T�b �` �` �
�G�n���X �i�Y � ����X �v�Y � ���` �x���X �i�Y � ����X �v�Y � ���` ���B�	�	ɩ�
� �	����
�
ɩ�
� �
� ����ɩ�
� ���� ��Lx� �� �� �� R� ��z�h`HZ����Z �] ���[ �
����T ȹ� P�U zh`!���j���ҧ!	 ��� �? � ���?   ���? � ����?  ����� �: ����   ���� �: �����𪪪�� �� ����  ����ê� �:��������>����ê��� �����ê��:��j�:��j�ꬩ������� �����ê��9k�V�:��V�ꬩg���eU�  ��eU����g9[�UYꫥ��֬�g�s�e�?  p�e�?��e�e5[f]Y֫UUU�lY�UUs�U   p�U �eUUe5WVsU�WUUU�\UUUUsUU�  pUU��UUUU5WU�U�WUUU�\UUUUsUUU  pUUU�UUUU5WU�U�\UUU5\UUUUsUUU  pUUU�UUUU5WU�U��_U�\UUUUsUUU  pUUU�UUUU5WU�U� pU5 \UUUUsUU�  pUU��UUUU5WU}U� pU5 \U�UUsUU   pUU �U�UU5\UUU� \U5 \UWUsUU�?  pUU�?�U5WU5\UUU5 \U5 \UWUsUUU� pUUU��U5WU5\UUU pU5 \UWU�UUUU �UUUU�U5\U5\UU� pU5 \U\U�UUUU �UUUU�UpU5\UU5  �W pUp� _UUU  _UUUW�U\U�   � ���? ����  �����  ���             ��              ��VY�      ���
  �UUUUU	      jUe�
 `UUUUU%     �UUUU��ZUUUUU�     `UUUUUUUUUUUU�     XUUUUUUUUUUUUU    VUUUUUUUUUUUUU�  �UUUUUUUUUUUUUU�e �UUUUUUUUUUUUUU  VUUUUUUUUUUUUUU� �UUUUUUUUUUUUUUUD"�UUUUUUUUUUUUUUUUP�UUUUUUUUUUUUUUUh��`UUUUUUUUUUUUUU�  ZUUUUUUUUUUUUUU�   VUUUUUUUUUUUUUU%   TUUUUUUUU��UUUU)   XUUUYUUUU% VUUU
   �e���UUUU
 hVU�    �
 �ZUU� ���
         ��U
                ��               �     D�V     �XU�JD�VUUUeQ  aUUU�   �*UU     �Z�      �           �               �Z���            �VUUUV� �
     ��jUUUUUU�f�
   �e�VUUUUUUUYUU   jUUUUUUUUUUUUU%   VUUUUUUUUUUUUU�  (iUUUUUUUUUUUUU�  �UUUUUUUUUUUUUUUPEUUUUUUUUUUUUUU� %UUUUUUUUUUUUUUe �VUUjUUUUUYeUZZR   ����UUUU������        VUU�             he�              ��*         ���������������������� � � �?@�����������G����� �
�� /d��     �

		�
	� ���� ���� ���� ���� ���� ���� ���� ���� ���� �8��� ���� ���� ���� ���� ���� ���� ���� ���� ���� �8���     ����������������������}8����������������������}8�     � C�� _�� 8�� *�� �� #��     � _	�� Y	�� T	��     � C��     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ���ة��  ��� �� �
� �ύ& ��"  ݃� t ����T ��U �� � �T����U ��� ��XL �@H�Z�s�S ��� �� ��' )�� � ��2� ��������# �$ �% (z�hX@                                                                                                                 ���c  � K��n���#  � �� �� ފ� �J  H� E� N���� �� �Ā� P� � x� Ŝx �2� ��0������&  	��0������&  � �� M� 4խl��l����������� Z���� k� �� s� �� �� }� �� V� I� �� �� G� � ,ƭ����n �ŭ����4���,�  ���%�)�� �ĭ  )���ύ& L� ��La��)��� i�Lq��ύ& � � � �  � R���� +����� �J  H�L:�L��ύ&  Y���� ����L=����� ��n��L��)�
���&����)�
�������)���ɖ�i���)����5�8����l�q�) �l�k�g������������l �í�����������������j�������$��������i�j��8��k��M  {��)����L�é�������/ �à ������i��������M  {��H���؀A�� �à ��-ȹ�(��i���8�����8��ș��M  {�������`�������������i�`Hڭ��n��8��o� ����O��ɪ�H��D�o��o��o8����/���n��n��n8�������n��i����o���Х�h`H�Z� �� �� $� � �� �� �� 9��� �ɭ�8��0
�� q� z� ��z�h`Hڢ(�  �� ������h`H�  ����h`Hڢ�  ��� ������h`�Z�à���������z�`�Z�(��������z�`Hx�΍& � �  K� � �� �� �ĭ  ��� �� �Xh`Hڢ�������
����������
�����������������������x ���h`H���%��� �x ��
�M  {��x ��8����d���h`Hڭ��n�� zʪ���Z �] �
�[ ���X ��m��Y ��8�Y �[ ��[ �.��X ����� ��� ��������8��������������h`Hڭ��0�������&�������� Ŝ�������������h`H�Z����8��0L�Ʃ���� � � � �  �� � q� �ɽ4� zʹ��Z �] �
�[ �9m��X �>m��Y  ����S ��H  � �� ����б �� � q� �� �ĭ���
��������8�n��	������0��8�������i�����zh`H�Z���u�Z ���[ ���X ���Y ��8�Y �[ ��[ �Y ����D�V ���W �Z �X �V)U�V�����Y �[ ��z�h`H������h`H���$�����������������s)i��h`H�����M  {����i��ɨ���h`HZ���F��8��0=��9��J�3�� zʨ���Z �] �
�[ ���X ���Y ��8�Y �[ ��[  �zh`H�Z�T �@�U � � � �T����U ���z�h`Hک�X �
�Y � ���f  �������X �
�Y �� �����)�X ��f  �������M  {��
��h`H�Z���d� zʭ�8��X ���Y ��Z �] ��[ ��8�Y �[ ��[  � zʭ�i�X ���Y ��Z �] ��[ ��8�Y �[ ��[  �� zʭ��Z �] ���[ ���X ���Y ��8�Y �[ ��[  a�� zʭ��X ���Y ���Z �] ���[ ��8�Y �[ ��[  ����;��� zʬ���X ��i�Y ɪ�^���Z �] �
�[ ��8�Y �[ ��[  ����9��� zʭ�i�X ��i�Y ���Z �] �
�[ ��8�Y �[ ��[  ��z�h`HZ���@����� zʨ���Z �] �
�[ ��8��X ��8��Y ��8�Y �[ ��[  ��zh`H�Z�k�a8��0)��%�i� zʹ��Z �] �
�[ �j�X �k�Y  �o8��0)��%�o�Y �n�X �m� zʹ��Z �] �
�[  ��z�h`HZ
����T ȹ�� P�U zh`Hڭk�s8��o� ˜k�c�k8�o��i��j +�i��oi�k�n�j�9�j�j�n�	�n8�j�8�n�i +�i�����j��j�k8��k�h`Hڢ ���@����9�o8����.���n�&�������+��-��,�������M  {���ж�h`H�Z� ��V ����O�� zʭ��Z �] ���[ ���X ��Y ��'8�
�[ ��8�[ �\ m\ mT �T �U i �U ��Y  ���Рz�h`H�Z�



����[ ��Y ���X �Y �D�V ���W �X �V�	��V�	��Y �[ ��z�h`H�Z� ��O����F p� �̽�;����0���8���"����,����8���	�8����Чz�h`H�Z��Y ���X ���[ �



��Y �D�V ���W �	�X �V�Ƚ	�V�Y ��[ ��z�h`H�Z���k��m��o��q� �v�/�p�*�ri�l�t�2��n��p��r ���� >�L����Ǡ �}�t�$�p�� "� ����b ��L����  "� ����L w�L� "� ����< ��L��!��  "� ����& ��L� "� ���� ��L� "� ���� r�L���Ђ� ����L���2�EZ����p�
�rz���l���n ����#��i��i �ة0����M  {�L���Ш���0����u�p���r���l���n ��������M  {����z�h`Z����p�
�rz���l���n`H�Z���v� �}�!�l���n�	���������)i�}�����z�h`H�Z��������i�
�
��}���&�������	�����ރ�����M  {�z�h`H�Z��������
��}���z�h`H�#�} ��h`H��} ��h`Hڹ�8������} �Ӏf� �}�� ���R�8�


i3����P���������s)������I�i��s)i�4�l� �� �ۀ��Ф�h`H�!�} ��h`H�Z���Lgҭ��l���n���p��8��r� �}�L_��$������o�
�q���k���m ����ٽ}��A��5�[�!�"�*��i��i �ة*�}�����S����}�I�����}�>��i��i �ة)�}�������i��i �ة(�}�������M  {����L�Ϣ ���Lѽ��+������o�
�q���k���m ����ֽ��,�"�0��� ���2��0����M  {�����W���M  {����G��)�Z �$mZ ����i���Z �Z ���Z ��mZ ��i �ة
�����M  {����LiЭ��1����8��o�
�q��8��k���m ��������������LgҢ ���2�O����o�
�q���k���m ����/�0�����Ν� ����������.�����	�M  {�Lg���Х���.����u�o���q���k���m �������ΝLgҭ��t� ���h��u�o���q���k�	�m ����H�����Ν�;�����
������)����������������.�����	�M  {����Ўz�h`H�Z� �p�:�|�b�x�]����p�	�t�z)��2�x�:�r�z)��B�v�z�-�t��i�i�tɪ��p��{��p���p��p��Џ�{���{�{z�h`H�Z� �p�L�ӹt8��0����r�X �t�Y �0,�pi z�Z����Z �] �
�[ z��8�Y �[ ��[  a�p z�Z����Z �] �
�[ �` z�r�X �t�Y ��*8��[ �` 8�[ �i�Z  �mT �T �U i �U ��Y ��8�Y �[ ��[  �����L��z�h`H�Z� �}�L�Թ�8��0�����X ���Y �0;�}����0�#�,�}i z�Z����Z �] �
�[ z��8�Y �[ ��[  a�}�$���i����� �}�m�} z�Z����Z �] �
�[ �` z���X ���Y ��1m[ 8��[ �705�` 8�[ �i�Z  �mT �T �U i �U ��Y ��8�Y �[ ��[  �����L��z�h`H�Z� �}�^��M��D���������}���}���}������0
��}�����0��i����������ɪ��}��И������Λ�z�h`Hڢ �j�x����q���g�8�
���l���n���sJ��
ms)i��������j i�j �k i �k �l i�l �m i �m �n i�n �o i �o ����Џ�h`H�Z� ���Lg�8��0����Z���'���Z �] ���[ �` �
����T ȹ�� P�U � zʹ��Z �] �
�[ �` z���X ���Y ��2m[ 8��[ �705�` 8�[ �i�Z  �mT �T �U i �U ��Y ��8�Y �[ ��[  �����L��z�h`Hڢ ���)ɩ���� �����(����� �� ������������h`�����J�ޞ���`H�Z�����7�


}�ɛ���� �,�������Z ���,�[  
׀����z�h`H� �\ �] ��@��T�Z ��������\ ��8�Z �Z �h�[ ��������] ��8�[ �[ �|�T�Z �,�i�Z �@�j +�i��
JJJ�h���T��h�|�(�j�Z �i +�i�|��h�T���|���h�h���|���\ ��@I�i�@�] ��TI�i�Th`Hڢ �,�K @ؽ,�Cސ��}@��h��ޤ��,}T�,�|���,ɪ�������,��,��Ы�h`HZ������L�ح��l���n���p���r����o�
�q��k�,�m ����F�,���Ν�9����
������'����������������.�����	�M  {�zh`H�Z� �,�?8��09��5�Z� zʹ��Z �] �
�[ z��X �,�Y ��8�Y �[ ��[  ���зz�h`H�Z������8��0	�����L��2�M����F�Y ���X ��8�3ZH
��q�T ȹq� P�U h����Z �] ��[ z��8�Y �[ ��[  a��Z� zʹ��Z �] �
�[ �` z���X ���Y ��1m[ 8��[ �705�` 8�[ �i�Z  �mT �T �U i �U ��Y ��8�Y �[ ��[  ��� �L)�z�h`H�Z���L��ξ���L�ۭ8�


i3�Z ���)��t��j� ���[�pmZ ���v�P�)�[ �s)m[ i������s)������I�i��s)i�4�l���� ��L����ЛL�ۍ[ �������\ ���] ���Lv���] ��8���)�` �s)m` i�] �_ �a ��b �v���s)i�] ��a �b �pmZ ���] ��ma �] ����_ 8�b �_ �l�s)������I�i��s)i�4�v�P�� ����[ Т�ʭ�����m] ��\ �L�ڱr���z�h`�P��F��7�	�F�
�W��S��O��L?������LK������L����L��L�ܽ��������L�ܭ��
��� ���4L�ܽ����s)i�����s)i#������4�P���J��
�sJ�������h������4����
����4�������������&������,�����������'�����4������� `H�Z�s)i�������� ��L�ݜ��� �� ���L}��2��������J�������l0m�P��6��2��3��/�	�0�
�1��-��)�� ����������� �݀ �݀ �݀
 .ހ cހ ��0�,�����ɪ����l�P�������� �����L�ܭ�����z�h`H��}����}4��h`H�l��Ji�4 �ݽl���l�I�i�h`H����� �݀K�4���?���: �ހ5���4�P�	�$���4�P�����)��������� �݀^4h`H�����4�P��� �݀�
8�l�4 �ݽl���l��h`H������4�P������� ��h`Hڽ��9�2�5�P����*�����"�4�P������� �ݽ�0�-�����н�h`H���#����������ޤ������(� ��h`HZ� �,�����Z ���,�[  
�ވ��������zh`H��1�1����� ��L��� �������8�

�����C��h������L�ߩH�������2�z������������2�d�s)i�� ���s)i������������3��2�2�������������3�(�2�������������2�3�h`�	�Z ���[ � ���\ �Z��[ ���\ �Oi�\ ����[ 8��[ �Z ��`HZ����3�L�������8�����ؐ����u�Z �] ���[ �` �
��E�T ȹE� P�U ���X ���Y ����.m[ 8��[ �` 8�[ �i�Z  �mT �T �U i �U ��Y ��8�Y �[ ��[  �����8���� ��zh`H���8���1����������� W� �� �� �� .� c�h`H��0��	i��L���2�2�
��~��z�[��2��[ ��i�\ ��i �] �^  ���[ ���\ ��i�] ��^  ���i�\ ��i�] ���^  ��L���m������"���I�i��h`H��m��������#������3I�i�3���m3��� ����{����3�2�K��2��[ ��i�\ ��i#�]  ���[ ���\ ��i�]  ���i�\ ��i�]  ��h`H��m��������$�������m3������Ʌ����3�2�P��2��[ ��i�\ ��i#�]  ���[ ���\ ��i�]  ���[ ��i�\ ��i�]  ��h`H��m3���3�0��Ʉ����3�
���H��3�}�2��(�2��3�l��m��������"������2����F��[ ��i�\ ��i#�]  ���[ ���\ ��i�]  ���i�\ ��i�]  ��h`H�3��3�3�
�������LF��m����
�����������i��ɩ���3�`�2�[��2��[ ��i�\ ��i!�] �^  H�
�[ ��8��\ ��i�] ���^  H��i	�\ ��i�] ��^  H�h`�] ��ɦ� ��`H�2�2�&��2��[ ��i�\ ��i�] ��^  ��1����)� �,���i��Z ��i�,�[  
׀����h`Hڢ ����[ ���\ ���] �	�^ �������h`HZ� ���R�	8��0I��E��Z��u�Z �] ���[ �
��E�T ȹE� P�U z���X �	�Y ��8�Y �[ ��[  ����Фzh`Hڢ ���L������7��D�	i�	�]���	i��	i	�	�	�P�A��}���5��}����&���	i�	�������J����������,��	ɪ������LK��h`Hڢ ����2��1�����������h`�	�Z �����[ � ���\ �h��[ ���\ �Oi�\ �h i�h �i i �i ���ԭ[ 8��[ �Z п`H�Z�h����|������ɨ� '߀j� ����H���o� ��ɪ��R��������O�O���H���\ �h���8����\ �Oi�\ �h i�h �i i �i ��H����z�h`H�Z _ˢ ��8�� ������ CĠ� ����8�������0� � _� CĀ� CĽ��0� ����@�� Cĩ�` ��i�\ �Y�8�\ �] �m] ����] �\ �[ �O�X ��Y �
����T ȹ�� P�U �T m] �T �U i �U  ����` п C� �z�h`Z�[ �O�X ���Y �
����T ȹ�� P�U  ��z`H�Z�_ �Y �D�V ���W �X �^ ��_ �T�^ �V�^ �_ ����Y �[ ��z�h`H�Z�Z �\ �Y �D�V ���W �X �^ �_ �_ �T�^ �V�^ �_ �\ ���T m] �T �U i �U �Y �[ гz�h`H�Z�Z �\ �Y �D�V ���W �X �^ �_ �_ �T�^ 1V�V�^ �_ �\ ���T m] �T �U i �U �Y �[ бz�h`H�Z�Z �\ �Y �D�V ���W �X �^ �_ �_ �T�^ V�V�^ �_ �\ ���T m] �T �U i �U �Y �[ бz�h`�ni�m�mr8��m�
�(�m�q� �l�k�mp�k����k�o����� `ڪ)�����	�)����`H�Z�Z �\ �Y �D�V ���W �X �f �V��\ ���Y �[ ��z�h`Hڪ)�JJJJ�f  ��)�f  ���h`H�Z�f �a��$��b��%��c��&��d��(����T ���U ��Z �Y �D�V ���W �X �T�V�T ȲT�V�T ��Z ���X �X z�h`ڪ��i�	��mi��� �`ک �i*�j��j�i����` 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p������������������������������������������aja�a2b�b�b^c�c&d�d�dRe�ef~f�fFg�ghrh�h:i�ijfj�j.k�k�kZl�l"m�m�mNn�nozo�oBp�p){)�)C*�*+o+�+7,�,�,c-�-+.�.�.W/�/0�0�0K1�12w2�2?3�3� G!�!"s"�";#�#$g$�$/%�%�%[&�&#'�'�'O(�( �L�LMBMlM�M���Fp1��ABTB`BlBvB�B�B�B�B�B�BC"C@CdC�C�C�C,D�DE�EF�F�F�F�F�FG4G[G�G�G�G�GHH3HKHeHH�H�H�HIKI�I!J�B�MN[N�N�O=PcO�O�MN[N�NsP�P�N3O�MN[N�N�P;QkQ�Q� ���� \� ��� @� ��t�\�aJ�KML�L 
	
		 		
$	�Q�QRNR SkS�R�R�Q�QRNR�S�S{R�R�Q�QRNR�S�STIT��`�����`��C��`�g���




	 ( 	  qT1�U�U�U1�W2WkW1�X�XZ1����0A1�9� 	 	 	  % % # # #  (2<FPZ� ���%�+ � ��$ � �% �  F��+ �+ �& � �� ���%�8 � ��1 � �2 �  ���8 �8 �3 � U� ���X� ���� � �� � �	 �  |� ���� � �� � � �  ��� � �
 � j�� � � � �� � ��`� �� ȱ�	 ȱ�
 ȱ� ȱ� )
��x�� �x�� � )0� ȱ����H �S Ȍ � � �
 � �LT�  @�� �� � �� ��Ȍ � ���! �"�$ ȱ"�% ȱ"�& ȱ"�' ȱ"�( )
��x��) �x��* �( )0�- ȱ"����H �S Ȍ! �+ �, �& � �� � � �M )����� �.  U�`�. �/�1 ȱ/�2 ȱ/�3 ȱ/�4 ȱ/�5 )
��x��6 �x��7 �5 )0�: ȱ/����H �S Ȍ. �8 �9 �3 � Ш� � � �M )��@З��� �!  ����� �� ȱ� ȱ� ȱ� ȱ� )
��x�� �x�� � )0�  ȱ����H �S Ȍ � � � � Ч�  ^�� �� � �� ��Ȍ � ���J 
����K ���L �K� ȱK� `�J 
�� ��K � ��L �K� ȱK� `H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; � �8�� �� )0� Ȍ ����� � � �; � z�h`H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; �  �8��  �� )0�  Ȍ ����� � � �; � z�h`H�Z�' )?	@�; �' I��-; �; �, �)��( )@��J��; �; �- �8��- ��( )0�- Ȍ, �)����, �( �, �; � z�h`H�Z�4 )?	@�; �4 I��-; �; �9 �6��5 )@��J��; �; �: �8��: ��5 )0�: Ȍ9 �6����9 �5 �9 �; � z�h`� `� `H�Z�H ���%�I ���H �O �I )?
����Q ���R �P  U�z�h`�O �* �G `�P �Q�C ȱQ�= ȱQ�> ȱQ�D )
��x��@ �x��A �D )0�E ȌP �? �B �C � K��S `H�Z�O ���LD��= �F �C I�F )��F �B �@��D )@��J��F �F �E �8��E ��D )0�E ȌB �@����B �D �B �C )�; �I )����
�@����; �; �F �( �; �G ��* �G �? �? �> � U�z�h`H�Z�  @�  ^� � �� �  j� �� |� �� ���� z�h`H�Z� � �
� � ��N �M )?�N �Q�� �K�N 
��4��" �V��/ �4��# �V��0 �! �. � � � �M )�����  U�M ���  �� �z�h` ��F� ��B� ��B� ��F� ��F� ��F� ��F� ��F� ��F� ��F� ��B� ��B� ��F� ��F� ��F� ��F� ��F� ��F� ��F� ��B� ��B� ��F��F� ��F� ��B� ��B� ��F��F� ��F� ��B� ��B� ��F� ��F� �T�T�  F� j�F� w�B� ��B� ���D� ��F�     � ��F� ��F� ��F� ��F� ��F� ��F� ��F� ��F� w�F� ��F� ��F� ��F� j�F� ��F� �F� T��t� _�B� j�B� q�B� �B� �8�D� �8�D� �8�D� 8�D� q��t� _�B� j�B� q�B� �B� �8�D� jp�T� ��F� ��F� ���t� ��F� ��F� j8�D�@8�D� �8�D�8�D�     � �8�D� �p�T� ��F� ��F� �p�D� �8�D� ��F� ��F� ��T�     �R�FBR�FR�F�R�FR�FBR�FR�F�R�FR�FBR�FR�F�R�FR�FBR�FR�F�R�Ff�FBf�Ff�F�f�Ff�FBf�Ff�F�f�FR�FBR�FR�F�R�Ff�FBf�Ff�F�f�FR�FBR�FR�F�R�Ff�FBf�Ff�F�f�F     �R�FBR�FR�F�R�F��FB��F��F���F��FB��F��F���FR�FBR�FR�F�R�F��FB��F��F���F��FB��F��F���F��FB��F��F���F��FB��F��F���F��FB��F��F���F��FB��F��F���F     �R�FBR�FR�F�R�F��FB��F��F���F��FB��F��F���FR�FBR�FR�F�R�Ff�FBf�F��F���F��FB��Ff�F�f�FR�FBR�F��F���F��FB��F��F���FR�FBR�FR�F�R�F��FB��F��F���F     �R�FB��Ff�F�,�F��FBR�FR�F�R�F     �     � ��� T�� %�� #��     � ���@��}�����     � �� q�� d�� _	�� ?�� 8�� 2�� /��     ��� f��@��f��     � /� �� �� 	�� /�� �� �� �� /�� �� �� ��     � �
�� ���     � _�� K�� ?�� /��     � _?� ??� %?� ?� /?� %?�     � ��� ��� ��� ��� ��� �������.��     � _
�� Y
�� T
�� O
�� K
�� G
�� C
�� ?
��     � _� � ?� �     � �� d�� T�� C�� ;�� 2��     �&�+�L�m�z����8   q/ p� p� p� q� q� q�    q/ p� p� q� q� q� q�  �( �  �    � �� � �_ �O �o ��  �$ 
�
	�
	 �
�



	�
	

			�
	
	 �"�*�������  �����  �.�.�.�.�.�.�.�.�.�.�Ϩ.�.�.�.�.��4�R�p������$�B�l���Q���M�w������������������ �F�                                                                                                                                                                                                                                                                                                                                                                                L� �M�