xآ���ɍ& ���  ��� ����� � � � �H�H�H� H� �� ������������� ��h� h�h�h���"���! � 0ĩ(�������� )��b� ���� � � ����� i� �i ���� J�� ���.�/���B w��)��0��0�.)�S�/��L�	��-���,��� }��/���-� �,���i }��/L%�@@@@@@8  0@P`8@@@@@@p�����Т �c�	�e8��e�����p��c�	�ei�e����������.i�.�.ɀ�L��d�ɴ�
�	���	��L�

��ˁ�c�́�g�́�k�΁�o�-�b�fi�j�n�,�e�mi�i�q���d�h�l�p`	
+,)*78'(56%&34#$12!"/0 -.� ���+��+��'�$����������(�� � %����� ���2d��3�1��W��X�i �� @ȥ/� ���	������ ���L��Lꂭi�2�� �LD��)��1�=�1� ���2m3�20�
��3I��3L����D�2���
�W�`�X�ւL�`PRESSSTART
��+�8�:��$�'��L�� ��� �W��X�$�� j��� ���� ��L�THIN CHEN ENTERPRISE
      PRESENTS


@1989:
     PENGUIN & SEAL

@1992:
     PENGUIN HIDEOUT


Design by:
     L.C. Tchacvosky
Artist by:
     Shyh-Dwo Maa
Music by:
     L.C. Tchacvosky  뽜$�%�&�������������������)�*�+��2� ������������������� )��+� ز n� ���ˢ� �� � 温��B������� ����� x��+����� �� ޴ �� ,� O� �����" ��� ��
���L�����������L��ӄ�
�
��ۄ��܄� ЄL��l     

������(�Z�[��������`��������`���敏��`���䩀��`��)�;��)�4Ls���)�*��)�#�����J���� w��� ��� �L&�`` �� n���W���X���� j��4�)��5��5�)�� � 䅭�6��6� �#��7�э7� �)Lu�CONTINUE     DIE �  䅭4I�4��5Lu��4���� ��LJ�H�4����W���XhL�� � �@�� �� � �������` )�� O��+��*�L�L�� ��b���`�
�W�@�X���� j��� ����$�!�-�� ������ ���/��)��1��1)� ��L`� ��L`�L����������Ŀ
�GAME OVER�
����������� ��W�@�X�䢆 j��+���� ���� �����2�� � ��L��< ��L�������������Ŀ
�!! FINISH !!�
�������������� �+�`���)�:�	�: H�LF��8�a�JJJJ�9�a�)�:�8 H�8`�9 P��
��ۄ��܄�l6@!@ !#! 1! @3@/?/?e���`�  �  ���  ����`@Hm��Hm��Hm�m � ���
��
���  I���
>���	��+����xL� .� ��h�h�h@�;�� �<� �����<m@�<�A��;`
�
e�� �9��<������;`�,
��� 8� � 
�@@ 
��<� TRADE MARK "SACHEN"�C��D���W�G�X�H� ���
���*�	�-��, � ��L��`�G�W�Xiɪ�骍XL��� �W��L�� ���H)�DhJJJJ�CL��HJJJJ �h)	0�:�iL����`�L�M�N ����O	0 ���`�E�FH


i�
��i �hJJJJJe��X ��mW���I� �
�JH�D��CJj.J.K
.J.Kh���J�ȭK� i��i0��i ��Iн ���E�F`�LH�MH�NH�� �O�����L8����L�M�����M�N������N�O��L�����Ly���LȭMy���M���о�L�Oh�Nh�Mh�L`���@B��' � d  
                                                                                                                                   08<80                                                                                                                                  <<  cc"     66666 ?T>~ac3c 6;nf; 00`     000   66   ~    0    ~           0` >cgksc> ? >c0c >cc> 6f `~c> 0`~cc> c >cc>cc> >cc?<       0 0`0   ~  ~  00 >cc  |�����| 6ccc ~33>33~ 3```3 |63336| 14<41 14<40x 3`oc3 cccccc << f< s36<63s x00001 cwkccc cs{ogc 6ccc6 ~33>00x >ccko> ~33>63s >c`c> ~Z< cccccc> ����f< �����ff �f<<f� �f<< C1 <00000< `p8 << 6c                  <>f; p0<633n   >c`c> 6ff;   >c`> 20|00x   ;ff><p06;33s    f<p036<6s    v{kkk   n3333   >ccc>   n33>0x  ;ff>  n300x   0> ~   ffff;   cc6   ckwc   c66c   33<  ~0~ p   pp ;n       6cc  ?_/W(T �����
(T(W/_?

����� �����     �����(T(T(T(T



 ��� �� ���     ?��     ���     ��� 4  b  � �� � ?�  � ���������!�����	���������q�pa� � � �  �@@@` ��,.((�h  `�  �        ������������������������  U�U�  ((((��������癙~~�����������$B��$$<<$$�B$(O��O(��                                                        ��ժ������U�U�����W�]����������������������������������ժ����U�U�����]�W�            �   �       �    �   �                                                                                                                                                        �        			`�������
�l`   �ff<8    �����`�` `����  >>6~`&<��~nz�>6   X� ������p	~d|a ؠ�`���?�?                                                                                                                                          �
��b����� �
������
i�
�i ��i��i ���ةb����X�W� � ������Xɨ��`�Z��WJ��XJJ���e���i ��H� �hz��\�]�



e�
�i ��JJJJe��X ��mW��� �
�ȱ
��
i�
� e��i0��i ���� ���]�\`�X�W���0�� iɪ�骍X�W`H)��/��hJJJJ�
ei@}?��` 0`��� P���@p��      �)��~�`�~���d�B����;� �B��� �L��WJJJ�
ȱ�X
mXe
��W)��B=
��1�B
��B�X
���mW�
��i �WXXX� �
 ���i��i �Lt�bz�����
":Rj������*�@ �B���� �c�C�eJJJ� ��������bJJJ���������i��i ��H� q�h�����в� ���`��[�b ��eJJe��i ��c�



He�
�i ��JJJJHe�he�he��i ��e)�\���Z��
�Y��
�\�8*.Y.Z8*.Y.Z���1�ȭY1�ȭZ1��Z���Y���\�
.Y.Z
.Y.Z���Q�ȭYQ�ȭZQ����i0��i ��
i�
�i ��i��i ��[�LŔ`�
��`���`�)��~�`�~���d�B0'� �D��_�C�^�E�`�F�aZ ��z�����۠ �b�C�c�D�d�E�e�F�c�Z �z�����ة �B`�b�^�c�_�d�`�e�a��[�^ ��aJJe��i ��_�



e�
�i ��JJJJe��a)�\�Z��
�Y��
�\�
.Y.Z
.Y.Z���Q�ȭYQ�ȭZQ��i0��i ��
i�
�i ��[�L>�`569:78;<-.12/034!"'(+, %&)*?@O ABPQCDRSEFTU	
#$GHVWIJXYKLZ[MN\]^_`a                 �@ePQTDDPEDV� � �f��?�9�>������DQU�ڪ֪��� �@��     P &��`E��`    U `F5�:�5 � W ��t���!`Ud@      * � �   � � � � � ���> � ������* � ������갪����       � �FZV�e��຀� �  �?�>����    UU @��������D�Q��ժժ֪����m � � ` �      ��� 4       ( ( h����B�Z�
��+���:�;��j� ����������*��_ �.�.�����/������������
��
�
�*�*��z��� �     � � � � � �  ? O p ��� �    � � �À� � V        ? �   � � 0   � k�k? � � ?H
U	 �  ��_  � ��A  2 <�? @B�A� � < ���� �� � � ��$   �ꪊ�*�*�~��  ( ()
�
�
�*�j � � 0 � � � ��   �u  5 �  �  4@ ] � \ G    ? � � ���_��������  � � � � � 7 < �      � � < �������?O     � \ ��O�?�_�       � �    � u � }�5�_�A     � ������p�����C  @@@?� � 0 ? � p�|  � �  � ?�?��P� ���      � � ���������   ? ? ? � � �   � � � � � ���   ? ? ����?���?��0���?   ��?���� ������?����0 �?�?�?���     @ @    P  �?���?                 � �                          � � �                     � � � � �                � � � � � ���          � �
�*��������@�@�         * ��
 � �����@�@�`U`U   
 
(
(*�����         � ������
�*���:���*jj   ��(�(�*�
���* � ":VVU	U	 �               � �                            � � � �                       � � � � � �                @�h����j�j�� � ��*��������T��*�*`U`U`U�U*UP    �����*�*�
���
�����j�Z�V��
��j�)�*�
�
�* 
 �j�j�����������*U	U	U	U*U��              @ A�V�?���?    �U % � �j���� �@
�*�������*
    �����������������?          �� � � � � � � �                �              ������ ?    ���� � � � � � ��� � ? ?    ������������ � ����?�?���� ? �� � � � � � � ��� ? ?     ������������ � �       ? ��� � � � � � �����                              �? � ���?������ � � �����������      � � �          ?���      � 0 �� � � � � � ��?       �� � � � �    �?�����?�?�?��� ���� � � � � � ����� �  ? � � �������������� ����?�?����  �� � � � � � � �� � � ?  ����? � � � � � �����? ? ? 3   ?�? � � � � �������           �?� � � � � � ��?�?����� � ? ������ � ����� ����? � ��� ���������� � � �? ? ? ?   ?�� � � � � ����� �� � � � � ����  � � � � � �0��������?    ������������ � ����� � � ? ? ? �������� � � � �   ?   ?<�� � � � � ����� �    ? ? � ��?� � � � � � ���������?    ���������� � � �������� � ? �������� � � � �    ? ?����� � �   � ����    ? ? ?���?� � � � � ������������������������� �   ��������������������?����������������������������?�������������������������?�?��������������������������������� ���      ? ? ������������ � ��� ? ? ? ?   �����������   ���������?�?  ��   �   � � ����?�����   �� � � � � � � ��?����������������?�������������������������������?�?������������������������� ����?�?��������������������?     ? �� �         � �    � �����     � � � � ��          ��  � � � � � �����       ? ? � � � � � �?��������������?�<�0 ��?�?�������0�         � ?� �      0�������                                                                                                       	
                                  	
        !"#$%&                                                                                                                                                                                                                            ����������������� ���?�?�?�?�?��   ����? 0 0 0�?  ��� �����?�?���?\5\5\5\5\5\5\5 <�?�?�?�?�?�?�?� ���?�?�?�?  �?�?�?�?�?�?�?�?�WWWWWWW�?0000000��������������           ���   ����  �? 0 0 0�?����������������\5\5\5\5\5\5\5�?�?�?�?�?�?�?�? <  �?W5W5W5W5W5�?�?�?�?�?�?�?�? ?WWWWWW�? 0000000�?�?�?�?�?�?�?�����?�?�?�?�?�?�?�?���MT��OT��OT��O � �U�U5�?U5 � �������������? ���:�?���������������� � � �TUTUTUTUTUT T T �����?�?�?�?�?�?�?�?�?�?�?�?�?�?T��OT��OT��OT����?U5�?U�U�  ������������ � ��������:�?��?  � � � � � � � �T T T T T T T T                    P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������<�Z�x�����ҫ��,�J�h�����¬����:�X�v�����Э��*�H�f�������ޮ���8�V�t�����ί�
�(�F�d�������ܰ��UUPUUPU�P^ePYYPgvPZ�@UUPUUPUUPU@UUPW�PVePYY�gvPYY�VePU�PUUPU@UUPVVPVVPVvPV�PVvPVVPVVPUUPUUPV�PU�PUePUePUePUePZ�PV�PUUPUUPUUPZ�PY^PY�PY�P[VPZZPUUPUUPUUPV�PV�PVYPV�PV�PVYPV�PViPUUPUUPZ�PUnPUYPUfPY�PV�P[�PZ�PUUPUUPZ�PYUP[UPz�P[UPYUPYUPZ�PUUPUUPUUPe�Pf�Pf�PnnPeVPj�PUUPUUPUUPU�PZ�PU�PZ�PU�PZ�PU�PZ�PUUPUUPUUPUVPi�Pf�P[�PV�PY�PeiP�UPUUPUUPV�PV�PVfP^VPZZP]UPZ�PUUPUUPUUPYePYePYePY�PZ�PU�PUePUUPUUPUUPVYPVYPY�P[�PVYPVYPUUPUUPUUPV�PYYPYYPYYPY�PYiPYyPV�PUUPUUPUUPU�PVfPV�PZfPY�PZfPV�PUUPUU�j��eU�fn�f{�fU�f��eU�j��UU�UUPUUPZ�PY�PZ�P[UPZ�PYyPZ�PUUPUUPUUPVZ`Y��m�Pj�PkePY�PVVPUUPUUPUUPUUPZ�PY�P[�PY�PZ�PUUPUUPUUPUUPV�PVvPVfPV�PU�PV�PUUPUUPUUPZ�PYBPY�PYfPXPZ�P[^PZjPUUPUUPUUPUUPUUPe�P���^�PUUPUUPUUPUUPUUPUUPZ�Pgw����YVPYVPUUPUUPUUPU�PVYPYmPVYPW�PVYPUmPU�PUUPUUPYe�e�P^YPY�e�PVYPYe�e�PUUPUUPVePU�PV�PW�PU��e�P[�PV�PU�PUUPUUPV�P[nPVyPU�PU�PVYPYVPUUPUUPUUPV��[[Pj�PUUPUUPj��UUPUUPUUPUUP���ffPYYPUUPYYPf�P���UUPUUPUUPZ�PZ�PY�P[YPY�PZ�PZ�PUUPUUPUUP]�PYVPY�PY�PYUP^�PUUPUUPUUPYe�VfPU�PU�PZ��U�PU�PVfPYe�UUPUUPU�PU�PZ	PYmP[�PZ�PUUPUUPUUPUUPUVPUY�V�`Y�PefP���VU`UUPUUPUUPeU�iV�f[�e��nY�iV�eU�UUPU�PV�PY�Pi�PZjPZ�PZ�PZYPV�PUUPVYP^[PjZ�eU�eՐeU�eU�jZ�^[PVYPUUPU�PZ�P^[P��YVPZ�PUUPU�PUUPUUPUZPVnPV�PV�PV+PU�PU�PV�PUUPUUPV�PZ�PYYPj�Pg�PjjPeVPeVPUUPUUPUUPUZ�W��Z��V�PV�PV9PU�PUUPUUPUUPVYPV�PZ�P^iPVyPVYPV�PUUPUUPU�PZePY�P[�PY�PZ�PVYPZ�PUUPUUPUUP���ff`jj`UUP���ff`UUPUUPUUPUUPf�Pi�P[�Pi�Pe�PnUPj�PUUPUUPUUPUUPVfPU�PV�PU�PVVPUUPUUPUUPUUPZ�PY�PYiPZ�P[�PYYPV�PUUPUUPUUPUiPU�PV�PZ�PV�PU�PUiPUUPUUPUUPUUP^�PY�Pb�Pi�PVPh�PZ�PeUPeUPeUPjuPU�PU�PU��U��UU�UU� T��p����� �J���)`)H T���=P����p��h� �
������`?�����
m�����JJm����)�`  ���

������
�WH���ı


�X�ѱ m��ұ m��Xi�Xh�W�ӱ m��ԱLm� 
 
====� ���������t��� t�� �����������d��` 										                   										�c�������t����  z�� ������`��� ��2
����� ����!� � ������`���L;�� �2L;�� ��L;�� �
L;�m$�$�m%�%��$�!�����`�$�!�%�"�&�#` z� �� �L���W�(�X���� j��!�L�"�M�#�N ����O	0 ���`HISCORE- �
�W�8�X�ݢ� j��$�L�%�M�&�NL��SCORE- �
�W�H�X���� j��iL��STAGE- ��W�X�X��� j��*L��PENGUIN- �W��X�I�� j���W��X ����WLȳHI-        SC-
      STAGE-









   [PRESS START]



   @1989 & @1992

THIN CHEN ENTERPRISE ��W�@�X�Ӣ� j���W�P�XL��HI-SCORE  `�����L���������)@� %���	@��)H���� �h� L���)���}P�����}T����
����JJJJ) ����)���`  ��    ��  ���
��v���w��l����ʵ����`�\� ����c����g����k����o����bJJJJ���eJJJJ��� -������L��)���5���� �b�f�j�n�L���L����+��w�� ���P ��hh`�)������JJJJJN�(.�� x�Lθ����`��� ����L������X�ye�e�m�X�yi�i�q�\�yb�b�f�\�yj�j�n��b)�|�e)�u�eJJJJ���bJJJJ��������Z �zΞ�5hhL��Z �z� ��e�b�� ��/�	���
����� -� t����� ����c�����������L9�`��JJJJ�	�JJJJ�
��o�0�	�'�s�0�
��P�m	���T�m
�� �� �`�����	�	�	�
����8`�� 	 	��� ��]ɀ�Y������M���	���
 #��>ɀ������-L޷����L޷����	���
���  -� t�8``�	���
���  -� t�� �������`�P�c�	�i���`����������������8�

�����c����g����k����o�




�b�fi�j�n�	



�e�mi�i�q�8`� ��i

�����c����g����k����o���b�fi�j�n���e�mi�i�q��d�h�l�p`�)����)��>�_�`�D�^�>�_���a`���#���� ��
��$���%��� !������`l8�L�L�L�L�L�L�L�n���`����c���������)����f� ���` ��  �����>����� e�) ������
���JJJJL������ w��L����J��P�}����T�}���)�ý�)м��L���)����JJJJJ^�(>���i�L�`� ���b��c�g�k�o`�

���H��H�b������c����g����k����oh�b�fi�j�nh�e�mi�i�q�` 0@�mmmm `��4� ����c�g�k�o��bJJJJ���eJJJJ��� -�Lt���J���� ����`� �����



�b�fi�j�n��



�e�mi�i�q�����c����g����k����o���I�� x��  -�Lt�H��� ��b��������e���Ȍh`��1���P�}e�e�mi�i�q�T�}b�b�fi�j�n`���`� ��L�����`���'���(��%�&�)�*��-�.� ����e�+�b�,� ������`���ߢ �������+���,� ������`����`� ����	� ������`���'���(� ���%�e�+�b�,� ������ -�� ����`����`� ����L㼹b�(�e�'���u�����b�(��e�'�芨������(��Z�zھ��bJJJJ���eJJJJ���� -�zLͼ��� �c�g�k�o������ �c�g�k�o�������LT�`�'e%f$8�+�jE$.�%e)8�.�$�$� �(e&f$8�,�jE$�&e*8�-�$�$�8``Hژ��=
�h�1h�0`�L�M� �LH
��a����b���� ^���0`l�g�u���� �L� �����`� �L� �����`� �L�( ��������L`� �/�B� �/��)�� ��k� ���"�� � � �( ����`d/ ���!�k����(�B�/��` ���/��`�(t/���!���L����8�9� � �8�0��������=� �:�0���@�A�B�/`�/�`�@��L9����A��A�`� �@�Bm�A�=�
�:�	�:�� L)������0�6�1�7�@� �60L����L����L����� �=����� ���6�Bm�A ��Lt���� ���6�4�68�4�6�7� �7Lt����L�������}�����6��7 ��Lt����- ���6H ���6H�}����6��7���h�7h�6Lt����' ���@���� �6�6������6i�6� e7�7�@Lt���� ���6Hȱ6�7h�6Lt����2����8)��8:�8� �9� ��6��b��@�:L� �� ��Lt�����@���)��8)�8�8�8 ���@Lt�ɀ�(逼��

��k��6�l��7�m��8�n��9 ���@Lt��@�0��������� ��� �8� �9�  ��� �6��b��@�: ���@
��6�0�7�1�@��0��0��`�?��<��<�L)�� �4���� �?LE���� ���4�@�48�@�4�5� �5LH�

� ���4��b��< ���J��( �K��) �L�)�* 	�* L)�   �6��7`�4��5`H���4
�5hJH��m5�5hn5n4��5�4`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   ����m��  ,����  &                                          �� �}¥����  ,��  
� 	 	�  � ! ���  &�  �  �  � & ���������  &(����  <(0 � ������������H�o��  ����  *		

�  �����*���  /	���  4(		��� ��@���������`�����[������d���͏���� �� Yŭ����魓����i<���`

�� ��ę � �����`� �/ ����ΐ`������@�]�<��8� ��i0�
�i ��������
����
�i0�
��i ���㭒���  	ƭ��a�1�]�-�D �����ȑ�� ��� ��i0��i ���ߩ��� ���_��a�Ș �ĭ��a�����`�`���Α`���M�]�I��8� ��i��i ��i0�
�i ��������
����
�i0�
��i ���㭓��� 	ƭ��a�1�]�-�D ���ȱ����'��� ��i0��i ���ߩ�����a�����`�`



}:ƅ
�;�i ��J��� ��>�e��i ���
���`@�@� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �  ͕�I�  �������=������2���	�- � �����W�8�X� ���Ii�b��<��b� j�L�Ȝ�`IIIIIIA*@XPP[cc=! 'I*!,'I,'=,;9; :,ccIIIIII9;,:,'=:i��������� ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� �  H  ������������?�� ���������?��?�� �?������� ?��           ]!D!JVUE  ���+�:|G�E�;�(����;�A�C�B�@�7�0���7�:�9�4�"�������  ^&.&.K5L?K^G_'^&  A,=.ICOCQ8A,  �I�N�O~O�U�U�h�r�wv���z҇�����x�v�o�e�[�V�N�I  �U�U�`�n�p�`�V�U  ��z�{����g�`�/���N�N�,�2�6�:�֏ԍ�Z�Z�}����������������ѮǸ�ǻֻշë�����������ڢ������������  � ����-x-w!s!p8fIbRkRsGv2�2�A�D�G�8�3�/�%�-�-�����  .'((9	8>D>6`$z	��)�)�)�3�6�6tG�O�Y�Z�N|LvYkek`eS]IrGu>s:q<iRCY?Y9O1I3D9594>A>.  �>�G{`iszj�W�M�I�E�>  �A�E�U�o�q�f�[�A  �W�W�r��d�Z�^�x�x��������������ةݥޡԙЛ̠��|����z�fÃҒ�������݋�{�e�a�\�W  ˦���݅���̦  � �
�
��&u&ggbgof�e�`�W�[�g�p�t�tV�V�W�p�������{�{�|��������㍡�����Ԭ���ݡޢ������������������������ܜ���{�{Ą΅с�V�V�Q�I�G�O�Q�Q�A�>�9�4�G�Q�Q�A�>�9�4�G�QuQt+�+�&��&�&�����
  .'((9	8>D>6`$z	��)�)�)�3�6�6uG�O�Y�Z�L{JwXlYkek`eS]GtCv8pRCY?Y9O1I3D9594>A>.  �V�V�u�v�v�V  � -&''9	8>@>2b }�	��(�(�(�2�5�5wG�L�T�U�I|GvRlSk_kZeM]Cs?v7r9jPBT@V:H0@9493=@=-  ��rt��%�/�$�)�3�:nGhHnL�B�:�>�L�N�E�?�5�1����  �Q�W�Y�Y�_�_�l�q�s�i�n�x�~������σҁۅ����|�z�n�f�b�]�Q  �Q�W�Y^Y`_�_�q�uiiin{zy�c�Z�]�v����������{�e�b�]�Q  ������U�O�R�����p�N�S�{ԗ����ݟ�����������������������������ާ����������  � -&''9	8>@>2b }�	��&�&�&�0�3�3tD�J�T�U�FwSk_kZeM]Av7pPBT@V:H0@9493=@=-  ���wtut>sTseg�[�[�e�e�b�!����  ���6�7�7��  �<�<�U�V�V�=�<  �m�w�w�}�}χ������Ȝ��ͷ�ȬЩԾ�Ӽݱ�������ݾ���������������}�w�n�m  �m�w\w^}�}��l�T�Q�_�z������i�K�I�^�ŏ����ݑ�~�r�r������ݠ��}�w�m  � ������  ��� + E`t	|wn&])Q*%�%�R�Y�^�l�p�q�c�v�}�{�t�p�a�\�Z�p�k�_�[�I�G�C�;�B�R�T�;�%�%� �� � ����  �)y/u26299�9�4�)  �>�@|EOF@>@kKiLd{d�g�e�N�J�F�>  {KLKL^M_|_|L{K  do_oG���1�1�/�'����)�6�;���������ܩ�������������މԔ���������w�diztxstdo  ��P�;�9�?���������  ՙ������֚֬ՙ  �>�>�?������  ձ���Í���ֲձ  �>�=�=�>Ā��  � �	�	��*t*tpn1dD^L]QiOq@s/�/�>�A�D�5�0�,�"�*�*�����	  MA	 X YM  P0C99@\@];P0  �A�JyJ|Q�Q�L�A  KU?]]dVdW_KU  �c�n�n{fxgxsx�w�wЃ҄������������w�s�m�d�c  �s�s����Ȗ�t�s  Kw?�V�W�Kw  K�A����������B�C�C�L�O�O�T�W�L�K�  Ǜ������ȿȜǛ  B����C�C�B�  ������c�]�`�������  � zzo(d:p8x)y��1�4�#����{z  L?	 X YL  �(�(�;�FiFlM�M�N�e�et]t����������_�bƣƤǣգ�����������������զ֮���m�i�e�]�_�d�e�M�M�H�@�>�F�H�H�5�3�1�-�(  Q1E99@\@];Q1  KU?]]dVdW_KU  �j�j����փ�k�j  �j�j�������k�j  Kw?�V�W�Kw  Ո������֡։Ո  ��������������  K�A����������B�C�C�L�O�O�T�W�L�K�  B����C�B�  � ���keh � �!�?�?r7r�}�~�ڈے��G�B�>�6�<�?�?� � ��  MA X YM  � � �?�?�!�   S2F;;B_B`=S2  �D�D�d�f�d�N�N�O�b�f�l�o�o�k�E�D�\�o�s�p�\�E~D~��ۃ�E�D  KW?__fVfWaKW  Ky?���V�W�Ky  ��������n�q�������a�[�^���������尺��کе������������  K�A����������B�C�C�L�O�O�T�W�L�K�  B����C�B�  � ����(�AvAh8hxh�g�g�`�R�N�U�e�o�u�uF�F�O�^�i�����Ώ�{��̽�����������������������Ȥ�k�i�a�\ȑƕ���\�F�F�A�9�7�?�A�A����  L?"X"YL  ����/�1�'� �  R2E;;	B^B_=R2  MUA]]dXdY_MU  �X�`y_|f�f�a�X  MuA}}�X�YMu  �~����~~~Ɉǉ��������������~  ��������������  ������� �B�C�C�M�O�O�T�U�K�G�C�"��  B� � �!�C�B�  � ����)_)b0�0�1�QxQmIjJjVj�i�i�v�vV�V�W����ܼ����������������Z�V�P�F�Q�Q�0�0�+��+�+�����  L?!X!YL  R2E;;B^B_=R2  MVA^^eXeY`MV  �^�l����~���������~��������ȡ��䮱ױجͤǢ��������׍؈�~�����m�i�c�^  �_�d�w�~����t�i�_  MvA~~�X�Y�Mv  M�C� ���������D�E�E�N�Q�Q�V�Y�N�M�  D����E�D�  � NBYZN  ���bd���\�R�D�5�/�+|(zDn]_lVrZung~Q�M�N�\�f�h�j�j�c�_�[�`�`�_�A�A�<�2�<�<���)�,�"���  V-I66=b=c8V-  LP@XX_W_XZLP  �r�}}tuqvq�q�p�p�}�}��������߾߲ܲ������������������|�s�r  Lu@}}�W�XLu  Ԃ}�}�~�՜ՃԂ  M�C����������D�E�E�N�Q�Q�V�Y�N�M�  ԡ}�}�~�ջբԡ  D����E�E�  � �
�
��=r=d4dodzc�c�Z�L�H�L�^�j�q�qB�B�Q�T�W�H�C�?�5�=�=�(�(�#���!�#�#�����
  I="T"UI  O5C==DZD[?O5  �J�J�Z�evhxl~o�m�l�����х���{�q�d�d�w�{�}�z�w�j�i�d�d�_�U�^�c�c�X�T�N�J  KU?]]dVdW_KU  Jy>���U�V�Jy  ْј͝����������o�rććˆ������������������������ۿ������ْ  J�F�B������A�B�L�N�N�S�T�J�  A����B�A�  � K?
VWK  ������V�T�L�L�T�R�O� ���  ���xiiYtWuL�L�V�T�Q� ���  ���F�G�G��  �uuFvG�G��  T2G;;B`Ba=T2  KS?[[bVbW]KS  �`�jujoirp�p�k�`  Jx>���U�V�Jx  �߉ފc�]�`���x�s�|�����̰���ܾ��ُݮ���������ٵ��٤Ѧͪ���������  J�@����������A�B�B�K�N�N�S�V�K�J�  A����B�A�  � ��tqrq@pVpg|i}^�^�h�h�e� ���  MAXYM  �}}6~7�7��  U1I99@`@a;U1  �<}<}X~Y�Y�=�<  GS;][bRbS]GS  �o�y�z]zWyZ������ۅ�{�}�����s�q�f�X�K�T�`�r�v��ԝ����������������ޫ���̩֝�������{�o  Gu;}�R�SGu  K�G�C������B�C�M�O�O�T�U�K�  B����C�B�  � ��|qnnn]msm�y�z}�}؆���#���  K?VWK  ���H�I�I� �  �zzH{I�I� �  T2G;;B`Ba=T2  �N�N�w�x�x�O�N  �NzNzw{x�x�O�N  KS?[[bVbW]KS  Jx>���U�V�Jx  ��������������  ���������������������ֿӾ�߷��ݐ�������  L�B����������C�D�D�M�P�P�U�X�M�L�  r�n�l�`�Z�Y�e�m�q�r�  ةԫڴ�����������ة  C����D�C�  � ��o(l,~+�*�)�GeGhNyNzOz{\y_�y�z�z�e�h�������^�a���������宸������ٳـ���{�q�y�{�N�N�I�A�?�G�I�I�&�����  MA
 X YM  V0I99@b@c;V0  �N�N�z�{�{�O�N  �N�N�z�{�{�O�N  KU?]]dVdW_KU  Kw?�V�W�Kw  ˀ������̳́ˀ  ��������������  K�A����������B�C�C�L�O�O�T�W�L�K�  B����C�B�  � ��} ppZpgo�o�g�Y�W�_�m�v�x�x����������覴��������ȴ�������������������������z����}|j�j�q�q�n�F�B�<�2�=~=}$�#�"�!�!� ����  NA"Z"[N  Y4L==DeDf?Y4  �B}B}d~e�e�C�B  OTB]]d[d\_OT  OzB���[�\�Oz  �ȊȮɯ���  ��������������  ��������������  ������� �E�F�P�R�R�W�X�N�J�F�"��  E� � �!�F�E�  � ������8�E�Q�K�J�E�9�-�"���  B6MNB  �r6\KSSkF�.�&�!��  O0B99@[@\;O0  �6�>z>}E�Eyjrw{y�t�e�e�r����������������č�v�j�f�`�Z�`�`�E�E�@�6  HU<_
]dSdT_HU  Gz;���R�S�Gz  ݙӤv�k�h�i�i�U�X������������ޚݙ  J�F�B������A�B�B�L�N�N�S�T�J�  ԩ�������ժԩ  �������䰪��  ��t�t�u�䌪��  A����B�A�  � ���pjm � ��  L? X YL  �/�:�:�2}3~?}P|f|w�y�m�m�v�v�s�C�?�9�0�/  Y2L;;BeBf=Y2  �?�?�g�h�h�@�?  MVA^^eXeY`MV  MxA���X�Y�Mx  �݊{�p�m�m�m�l�l�x�y�����������������  ޏ������ߴߐޏ  ��y�y�z�������  L�B� ���������C�D�D�M�P�P�U�X�M�L�  C����D�D�C�  ޹���ݲ���ߺ޹  ��y�y�zޥޤ�  � ����~~P�N�F�F�N�L�I�!���  OB![!\O  ���@�A�A��  ]3P==<
CiCj>]3  �Q�[�\j\d[gb~bc�f�l�p�t����������������b�b�]�Q  OVBa_f[f\aOV  �b�b����ׁ�c�b  NzA���Z�[�Nz  ֆ������ףׇֆ  Q�G�"�������� �H�I�I�R�U�U�Z�]�R�Q�  ֨���͑���ש֨  H� � �!�I�H�  � ����F|F{$�!�no*n@nTxU{Q{K�K�S�T�P�$�!���*�F�F�����  L?!X!YL  U2H;;BaBb=U2  MVA^^eXeY`MV  �^�h�iei_hbo�o����x�m�j�j�j�i�i�v�v�������ꛔ����������ޔޕ������������������������ݏ���o�o�j�^  MyA���X�Y�My  M�C� ���������D�E�E�N�Q�Q�V�Y�N�M�  D����E�D�  � ��'�'vv�}�t�t�~�|�/�*�&��$�'�'�����  QD]^Q  �,�,�J�K�K�-�,  \0O::9	@h@i;\0  �P�P�n�o�o�Q�P  OTB]]d[d\_OT  OvB��[�\�Ov  ��ԏӐk�e�h�������o�r�������Y�\��������������ӯɻ��������  P�F�!���������G�H�H�Q�T�T�Y�\�Q�P�  G��� �H�G�  � JD9!-51,6*@9B?HBK6D.<(NVVJ  poo!o�n�n�{�{���������|�{������~��|�{\�\�d�b�_�$� ����}p  �����!�!�"�W�V�\�\�g�e�b�$� ��  �!{!{V|W�W�"�!  ]5Y7MK4aqu"p;dBm<z*��!�6�E~IN�H�2���&�;�M�S�R�K�C�)�+�7�:�I�S�]�_�]�RzDaLXaBiBi<]5  9>"N%X+Y.V.K"=9  �q�v�z�z��������Ȯ܉�����������������������t�r�q  ݀����ʻѳܐ݀  � ����F�F�$�!�st*s@sT}U�Q�K�K�S�T�P�$�!���*�F�F�����  JD9!-51,6*@9B?HBK6D.<(NVVJ  ]5Y7MK4aqu"p;dBmCq-���8�D�J�L�N�8���"�<�P�S�R�K�C�)�+�7�:�I�S�]�_�]�RzDaLXaBiBi<]5  9>"N%X+Y.V.K"=9  �^�h�iiichfo�o����}�r�o�o�o�n�n�{�{�������꟔��������Ôߔߕ������������������������ޏ���o�o�j�^  � JD9!-51,7*A:CAHBJ@K5@*?$LVVJ  ��vx��-�@rRZ`Ydcb�P�8�#�<�T�\�X�V�R�D�.� ���  ]5Y7MK4aqu"p;d@eDp0����%�8�F~JO�:�$���'�A�O�S�R�K�C�)�+�7�:�I�S�]�_�]�RxD^UPaBiBi<]5  9>"N%X+Y.V.K"=9  �F�Q�O�V�V�Q�F  �h�szsoklllxl�k�k�x�x����Ñē���x�x�����������x�xx�x�y�ގ�ރ������ݤ|�x�r�i�h  �k�k�~����޶������������x�u�q�k  �w�w����������Ƅ́�|�w  � ��|qnon?mUmfzhz���h�h�e�"���  UK �����L�M�V�Y�Y"^aVU  LDEMEML  �.�7�7�>�>�9�.  LJJqrMrMKLJ  �L�U�U�\�\�W�L  �n�y�y{qxrx~x�w�w����������������~�x�o�n  Lww��M�MxLw  �~�~����֛��~  ՠ������ֽ֡ՠ  (����-�8�6�(�  H�D�T�X�`�b�`�R�I�H�  �߅�����  � �	y	y.0!y!z"z//.5y5z6zB.B0HyHzIzVVU\�\�W�K�W�W�H�H�N�L�I�5�5�0�$�0�0�$� ����������	  �!�!�/�0�0�"�!  �5�5�B�C�C�6�5  �b�c�f�u�~��t�i�b  7b's}�$�.x6i7b  �c�g�s�x�{�o�c  bc]cbqbxh{jykncdbc  �z�|��G�8z8�C�DͿ�������̊ц҂�z  ��D�D�E�������  ��D�D�E�������  ��D�D�E�������  e�D���!�a�d�s�q�e�  �חנ������������  � vvk(c1`8l6r.u��+�3�3�"����wv  TJ �����K�L�U�X�X"]`UT  KDELELK  �&�&�9�AjAmH�H�I�a{apYmZnfm�l�l�x�y�������]�`Ȟȟɞ��������������ìë�Ө԰ݰ��j�f�`�V�a�a�H�H�C�;�9�A�C�C�3�0�+�&  KJJqrLrLKKJ  �f�f����ԁ�g�f  �fyfy�z����g�f  Kww��L�LxKw  ӆ������ԣԇӆ  ��y�y�z�������  &����&�,�6�4�&�  F�B�R�X�Z�X�N�F�  � �	�	�&�'h'k.�.�KpIsP�P�h�o]m`t~tv�]�Y�[�b�}��t�t֎�������ـ�t�t�o�c�o�o�U�P�P�K�C�A�I�K�K�.�.�)�!��'�)�)����	  SI!�����J�K�T�W�W%\!_TS  J!!GHKHK"J!  JMMtuKuKNJM  �P�P�j�o�o�P  Jzz��K�K{Jz  ύˏǔ��}�}������������ӝؙٕύ  ƚ������ǻǛƚ  %����+�5�3�%�  D�@�P�R�Y�[�Y�M�E�D�  ������������  � }vw!w5Z3]:v:w;w_P_P'T#WKA #�����B�C�L�O�Od�d�v��º�Ԛ�����������������������������ϸ����z˩Ɯ�d�d�_�Q�_�_�P�������,�T�_�_�:�:�5�-�+�3�5�5����}  �"�#�&�4�B�B�?�3�%�#�"  B##IJCJC$B#  BOOtuCuCPBO  Bzz��C�C{Bz  ������r�c�c�n�oɕɖԠҢϢ�������  ��o�o�pĖĖ���  ?�;�I�Q�S�Q�I�@�?�  #����&�(�3�1�#�  � E	>	??,*1>1?2?UU\0\1]0�0�)����)�7�=�=\M\M]M�A�2�2�@�E�F�O�X�Z�Z\|\}WlKbWLWK1r1s,h$b"Y*Y,L,KUXUE	  �
�
��G�G�?�@�L�����đ�޸������P�L�F�<�G�G�*�*�%��%�%�����
  �L�L�j�k�k�M�L  �p�p����ߏ�q�p  vv��
���+�*}v  eya{e�q�w�z�y�g|ey  ޔ������߳ߕޔ  ��g�i��ұа̡�  ��������������������  � ;
4
55,*141525WU\(\)](w'�"����%�1�5�5\A\A]A�9�+�+�5�=�>�H�N�N\j\kWZKPWBWA1d1e,Z$T"K*B,AKNK;
  qpp!p�o�o�|�|���������}�|������~��}�|\�\�d�b�_�$� ����~q  �����!�!�"�W�V�\�\�g�e�b�$� ��  �!|!|V}W�W�"�!  �q�v�z�z������Ǳڔ����������������������׿����t�r�q  ss{�
�����~!z#vs  YxUy_�a�i�g�Yx  ܀����ɺηڕ܀  � B<==207<7=8=]
]d<d=e=�4�$�'�0����
��!�&�8�N�h�|���������������`�J�H�H�r�s�c�[�[�I�Hdwdx_hS^_I_H7o7p2`&V2I2HRURB  ������?�J�E�A�5�$� ���  ��=qL}G�7�(�'�!�  �1�:�8�?�?�@�[�[~T~ЈΉ����������c�_�[�S�Z�[�?�?�:�1  �?�?�[�[�@�?  �`�`Ƀ́�l�l�؃وЋ�����a�`�y�������s�a�`����ޠ�a�`  ݥ������޻ݥ  � @
9
::1/696:7:`
^e9e:f:�*�#�%�/�)}���	���� �6�K�]�z��������������[�F�F�s�t�i�c�[�[�G�Feyez`iT_`G`F6n6o1d)^'V/V1G1FPSP@
  ������_�]�W�W�^�\�Y�#���  � � �5�6�6�!�   �;�;�Q�R�R�<�;  �f�pxprouv�v�w������������������z�n�r�Ë������ź���������󿼿�������ҋɕ���v�v�q�f  � �
�
�(p(j'm.�.�KrIuP�P�o`mct�t{�c�_�c�w�z�z������������֝ߘ������ۂ�w�t�t�o�c�o�o�S�P�P�K�C�A�I�K�K�.�.�)�!��'�)�)����
  TJ  CYjl\/\0]0� � �*�-�*z������R�d�b�=�=�`�a�V�P�G�=�=\K\L]LjUjXgX$] `UT  K  VWLWL!K   �P�P�l�o�o�P  �t�t}�����ɕώԎ�t  ɚ������ʻʛɚ  ������������  � YO#BXi k!^6^7_7�!�!�+�.�+z������X�i�h�C�C�g�h�]�W�O�O�D�C^P^QgZg]d]"beY  ���vps � ��  P!!X"YQYQP  �0�;�;�3�4�@�Q�g�x�z�n�n�y�y�v�D�@�:�1�0  �@�@�h�i�i�A�@  �ኁ�v�s�s�s�r�r�~������������������  ⏶��������  ������������  ⹶��ݷ�����  ���݀ުީ�  � ����/�/�������/d-g4�4�5��Y�\�n�n�n�n�x�{�{���������|�{эǙ�����������������������߸ݻû���������ۓѕ�4�4�/�#�+�/�����  TPL#jh \1\2]2���&~z������Q�d�d�>�>�c�d�Y�SK�K�?�>\K\LfVdXaX!]^T  K  V!WLWLK  �4�4�P�Q�Q�5�4  �V�V�s�t�t�W�V  �y�y����ĕ�z�y  ��{�{ʄƐ���  � |
v
ww2_0b7v7v8vqv������v�v�q�e�q�q�7�7�8�N�b�c�_�Y�Y�`�a�]�7�7�2�*�(�0�2�2������2�2������2�2���|
  TPL#jh \0\1]1���%~z������R�b�a�=�=�a�b�S�J�>�>\K\LfVdXaX!]^T  K  V!WLWLK  �7�7�S�T�T�8�7  �~�~����_�b�����y�X�\�Κ����ޥ��ﲫ�������������������������ۜ���������~  � �
�
��*g*j1�1�@|[aq^sax�b�I�=�]�q�r�n�8�S�h�p�p�j�j�f�Z�J�4�1�1�,� �,�,����
  TJ"AWhj \0\1]1���%~z������R�b�a�=�=�a�b�S�J�>�>\K\LfUfXcX"]`UT  K  V!WLWLK  �q�|�|�t�u�����ыӌ�����������؅݁�{�r�q  ˁ������̞̂ˁ  ˣ��������̤ˣ  ������_�Y�\�������  � ���{xyxAwWwh�j�_�_�i�i�f�"���  UQM"jh\1\2]2���&~z��	����Q�c�b�?�?�c�d�Y�S�K�K�?�?\L\MfWdYaY!^_U  ���9�:�:��  LV WMWML  �?�?�Y�Z�Z�@�?  �n�p�{h{bze������ڏ̃���������z�x�m�_�W�`�o�}āƋՠ����������������߮���ԝʩ������|�n  � ����� B~X~i�k�^�^�i�i�f�$� ��  XTP"jh\1\2]2� � �&~z������R�c�`�?�?�b�c�T�K�?�?\O\PfZd\a\!abX  OV WPWPO  � � �:�;�;�!�   �@�@�X�Y�Y�A�@  �j�l�wlwfvi}�}��y�^�X�\�y���������f�h؂ʛ����������Ǔ�w�|�۵�ǰКߚ����������ߩ��������������������}�}�x�j  � ��p%p(�'�'�%�$�?�?x7x{�y�o�o�p��{�p�m�m�m�l�l�y�y������������͖�Ʒ˻������Դơ��Ư������������������������������������Ᏻ��o�o�x�v�s�G�C���`�`



}:ƅ
�;�i ��J��� ��>�e��i ���
���`@�@� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� xة�& L �������