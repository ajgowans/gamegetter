� 
��=��] �=�i��^ ���[ �A�\ � � �]�[��(���[ i0�[ �\ i �\ �] i(�] �^ i �^ �����L��                                                                                  �                                                                            �                                    "�                                     "                                     "�                                    , ��                                    ,��                                    ,���     �������������������  ���?      ���     0                      0     ,���     0                      0     ,���     0                      0     ,���    0                      0     ����    0                      0     ����     0                      0     ����     0                      0     ����     0                      0     ,  �     0                      0     ���     0                      0     �  �     0                      0     ����     0                      0     ����     0                      0     ����     0                      0     �
 �     0                      0     ����     0                      0     �
 �     0                      0     ����     0                      0     ����     0                      0     �"��     0                      0     �"��     0                      0     �"��  �  0                      0     �"��     0                      0     �"��     0                      0     �"��    �0                      0     �"��  �  0                      0     �"��  � �0                    ���?     �"��  ��0                            �"��  ��0                            �"�� ���0                           �"��  ��0                  (         �"�� ���0                  (�
        ���� ���0                  *�        ���� ���0                  "�
   �  ����� ���2                   �
�
 �  ����� ����2                   �
� �  �� � ����2                  , �
�* �������������2                  ,  �*�� �* ���������2                  , �� 
 *�������"2                  ����  
�* �������" 2                  ������*���
�"���  8                  �������*� �"����*��8                  ���"���
��(��"��  ��8                  � ��������(��"�� �*�:                  ����*�����* �"��  " 0                  �(��
�
���*
�"��
��"0                  ����� ���*
�"��
��"0                  ����������* �"��
��"�2                  ����
 ����*��"�� ��"�2                  ����*��������"�� ��"�:                  �������������"��*��:                  �������������"�� ���:                  �������
  ���"�� ���:                  ������    ���"�� ���:                  ���      ���"������:                   �����������"�����"�:                  ��
  
  
 ���"��*��"�:                  �     
 ���"��*��"�:                           ���������"�:                           ���������"�:                           
��������"�:                  ��        ��
�����"�:                           ���������"�:                          ��������"�:                        *  ���������"�:                       �� * �������"�:                      ��*   
" �����"�:                      ��  
  *�����"�:                           
�**�����**0                           �  �����*8                           ���������*�:                           ���������*�:                           ���������*�:                           ���������*�:                           �����������:                           �����������:                           �����������:                  *        �����������:                  �        �����������:                  ��
       �����������2                  ��        ����������
0                  �
        ���������* 0                           ���������  0                           �������� �?                           ��� 3����0                           �� <       0                                  ����?                           �������   0                           ��         0                  ��               ���?                  ����            �   0                  ������?   ��   �   0                   �����������  �   0                     �������
 < ��   0                       ����� � ��   0                           
   ���
   0                  <           ����   0                  �    ����   ����
   0                  �   �      � ��    0                    ��       � ��*   0                   ����       � �
    0                   ���        ��
   0                   ���        ���    0                   ��*       �  �
   0                   ���         �
    0                   ���      �   �
  0                   ��          ��    0                   ���      �* ��   0                   �
�
        �    0                   ���      ����
 ��  0                   ���+         �*    0                  �*   �              0                    �
        ��  (  0                   �
��              ��������������������
   (        ��            �*          ��*             �*      ���   ��*        ���                     ���*              ��                       �*
          (�                            "                                  �          ����                      ������           ��                          ��        �                                                                                *                                                                                                               H�Z����� ��\� �� �0�A iL�E ��B i�D  ���� ��A i8�E �9�B i�D  ��P�A i<�E �9�B i�D ���  ����� ��A ih�E ��B i/�D  ���z�hLK�  �
 ���  ��
�* �
  �
����  ����* �
  �
���� �����* �
 ������ �����
�� ��������*�
�� � �*��*� ���  � �*����+  ���  ����
��*�+�*��*  ����
��*��������*  ����¯�*��������
  �
���+�*  ��* �
 ����
�*  �
�� �������* �
�� � �*����� ���  � ��������  �* ��� ������ �*  �* ��+ ������� �*  �
���
��*����* �
     ��
��   ��
  ���*�   ���  ���*�  ���� ��
�
�*  ���� ���*�*  �*�� � �
�
 ��
�� �+ �
�
 ��� ���¯ �� �� ������ �* �� �����  �
 � �
��  �
 �+����* �� �*����* ��
 �
� �*�
 �� �
� �*�
 ��
�� ���ʯ����*�� ��������*���
 ��������
���     �* �� �
 �*   ���
���*���
 ����
���
���
��
�*��ʯʿ
 �� �
�*���� �
�* �
���
�
   ��
   ��� �   �  ��* �   �   ���
 ���  �*   ��� ���
 �*   ��
   �
 �
 �����
   �
 �* ���*�
� �
 �
 �*�
�
�
�� �*��
�
�+�*�� ����¯�
����  ���*���+���*  ���
� �+���              �?                        ���?                     � ��                     �� �                     ���                     � �                      � �                  ��  �� ���             ��� �� ���            �VU �� |U�            �  = ��   >            /  � ���  �           �  ����  �          �  @lT|   �          �|   =lT   @>          o�  �_T�    �         �[�  PUU    �        �V|           �        �|             P>        o|    ��     P�       �[|    ��w     @�      �V|   |����   @�      �U |   �����    U>      oU �  ����    U�     �[ � �����    T�    �V |  ����� w  P�    �U | ���������� PU>    oU | �����������@U�   �[U | ���w�����@U�  �VU | ��������@U�  �UU | ���������! UU>  oUU@| ��������UU� �[UT�| ��������цU��V�������������AVV��U%%y����}�����mXXU>lUII^ |  ����� ���aaU9kUR�W    ��  �  @Ն�U����ZU�|UU���UU=_U�~�꫺�~���?�����������/�������       ��       ����           ��                      ��                      ��                      ��                      ��                      ��                      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��k �4�H �;�I  �   ����
�����/�� �N  ���N �k �k �0��k �;�I ��N�I  ꀿL��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          H�Z�0���
��K��< �K�i��= ��H ��I �����> ����? �	�<-N �>�< i�< �= i �= ��H �H � �� �̩�H ��I �I � мz�hL(�  ��             ���  ���?             ���  ����             ���  ����           ���� �����            ��� ��?��            ��� �?00�?   �       ��� �?  �?   �       �� �?  �?   �       ��� ����?   �       �_�   ��?            ���   ��?     �     ���   ��?     �     �W�3     �?   �?��?    �?0     �?   �?��� � �0    �  �����  ��?   ��  ������  <    ���  ����0  ���   ���  �?���<  ���   ���?� �3� �   ���  ����?�  ������  ���  ����?  ��?�?�   ���  ����?  ���?�?�   ���  ����?  �����?   ��� �����?  �����  ����������?  �?���  ,���*�����?  �� ��   ����������?           �����          �g ��H �P�I  ���   ���0������� �N  ���N �g � �
�g �P�I ���g �d�I ���g i� L;�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ������� ��A il�E �x�B i�D  ���L+� �                         0 ��0 ���?�?��??����� ?????0 ���� �?<????? 0?????�0 ���� ??? ????? 0? ????�0 ���� ??� ????? 0? �??�3 �����?�??�?�0? ????�? ��<� ??�????? 0?????�? ���� ?? ?????? ��� ????? ���� ????????  0 ��< ����???��??� �                                                                                       ���? �                   �<<����                  �<<����                  �<<�� �                  ��?�� �                   � < �                    �  <�                   �  <��                  �� ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�   % UU%        VUeUUVUe          Ve        UVUeVUeU           	 % � VY	e%�UVVYYee��VVYYee   V Ye�VVYYee��VVYYee��VV � X�UXU        U�UY�UYU         @ T@�TY        �UYUU�UY           � ` X V��`eXYUV��eeYYVV��eeYY @ P T �@ePYTV��eeYYVV��eeYYVV��   0      0      �0      33    �����     �;   �������?< �:<    <    (��(??���?������������������������������UUUT���?�?�?�?�?�?�?�?�?�5�5�5TTPP� ������wwwUUT T <������UUUU???7��?_���_��?����=�=���__�� ��� <�<??      T��T       @   P  P  �  � T�U�~T� �  �  P  P  @           @U   @Y   ��  �� P��_T��_���T��_P��_ ��  ��  @U   @Y                T    U   e  @�  ��  �� P���T���U����YT���UP��� ��  ��  @�   U   e   T                 ��?              �� � �*� � �        �� ��?� � �?    �         �         �         �         �         �         �        �        �
       ���?       �>    ���������� ����0     ��        <<                                        .        .       ��      ����     ��   ��������? �3���    ��                                   ��?     .   ������� ���33    �                    �,?   �  ����� 3��         ����?      �         �         �         �         �         �         �        0      �?��     ��   ��������� �γ��0    ��       �        �                                                        3      �?�     ��   ��������? �3���    ��       ?                                     3    ����    ��   ������? ����    ?     0    0    0    0   �3?   �  ����� 3�3  �   �             �      0                �  0 �0   � 0�        ��     ̯    ��    0�     ��    ���    0�?    �     �      0      �           �     0                      �    0          � �0  00�  ��  ��  ��  ��   ��   �   0        3   �    0                  �    0    �    �  �<   0?   �0   �   �          �   0    �                    0      �            � �   0 0   �0     �     <�     ��     ;�     0     �<    �    ��0     <�            0      �            �      0      �               0    �    0� �  0  3  ��  �  �3   �   �3   ��        0    �        �    0    �        0    �     �  ��   �<   �3   0�   �<   ?    �        �    0    �             � � 3  ��  ,  �  � ��  0  �   0                    0      �             �   3 0   �0    0�     ��     �     ��     �?     ��    �:    ��0     �            3      �      0            0      �               0    �    0� 0    3  ��   ��   ��   ;   �0            3    �    0        0      0  �0 03  �  �  �  �3   �   0   �                  �      0               �   0 �0  � 0    3    ��     �?     ��     ��    ��    ��    0�        �      0           3     �      0                      0           �  �0 0  03  ��   ��   ��   ;   �   0        3   �    0            @ � YT� �
�*�J�����f��"�IZP��U �@�� @�j  ��j	 QTR	 QUV� UV�UV�"UE�T!��%U�VQT(Y��H Z�j ��U D      ��V ����P��V�iVA�e�
X��YE�*��
��Ui��RU ( V@ ��R (e ��� ���Q@����U�je�j*d	�Z��JDVR �VYV�� PU   T     dU    PU�	   P    T�*U �U��VU d����U �Z��VV��iVU��e�
��Y��YU��*���$��Ui���RU ��%V@ �Q�R (e�� ��D�� ��T�U@��T��U�jUe�jjhe��ZV P���JT�fVR Z  �VYV  ���  ��V�  XfUU    AU    TU     �     ��    P��	  @P�   @ �  �VU� �F��
 ��
��* h���  X����� X��T( Z��A` (PB�eV% ��	� @�j
�Z@U"�T @TU
�U  DU)�U D�&�U�HU�UfUHf*hf	DU)P�UUZ	�FV�iZ
 ���Z�
@�f��@J�J @Y�PU*  �V��
   � * ����;  ���? ������ �   �� � ��� ������
��� �   ��  ���� �� ����������*��������  �    ���   ������ ���   ���*  �����? ������ ������������誫����믿�� �
 ��
��ww����* �� w������_���_www_���_���*  ���*  ���  333��*�����33333�����33333����������  �����  ����z  ����_���<��\���������<��<�s�������<��<�s������� ������   �����z   �����^   �����_       \��������ܪ��    ���z��������_       \��������\       \��������_       \��������\       � ��������?  �  ���������� � ��� �>���������  �   ��  ���� �����������������������   �    <�    ��  �����? ����������������������������������                               @                   �   �                      � �                            ���  ���                     �         �@             @   �            �                            �      �      �     �     �     �   � �@   � �   �     �    ��     ��                 �*  ��
                           � �         �    �   �@� �    �@  �     �    �      �     �      �      �           ������������������������������������������������������������������������������������ ��0���������������������������������������?��                        �������������?��                        �������� ��0��                        �������������?��                        �������������?��                        �����������0 ���������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU    @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU UUUUUUUUUU��������������������UUUUUUUUUUUUUUU������������������������������UUUUU����������������������������������������������������������������������������������������������ZUUUUUUUUUU��������������������������������������������������������������������������������Z�����������������������������������������������������������������������������������������������UUUUUUU�UUUU����������뿺~UUUU����������������j������������������~��������_���������������������������~��������_����������UUUU�����?  ���~UUUU����_�������������������   ����������������������������������     ��������������������������������~UUUVUU���������������������������    �      ������������    ����?� 0    �     @���3����0    ��??�����??    ��      @����<�<���?    ��?������??    ��     @��3�<�����?    ��?�� � ??    ��      @��3������0    ��?�����??    �;@UUVU@��3���?���?    ��?������??    �;@    @����<�<���?    ��?���<� ??    �;@   @���3���0    �����������    �@    @�����������    ����������������@ TV @�������������������������������@ @ @�������������������������������@ C @�����������������U��U���UU����ȏ��������������������U��U���UU���@ C @�����������������U��U���UU���@ @ @�������������������������������@ TV @�������������������������������;@    @�������������������������������;@   @�������������������������������;@    @������������������������    ����@UUVU@�����         �������?    ����      @����?         ���������?    ����     @����?         ���������?    ���      @����?    <    ��������?    ���     �����?         ���������?    ���>      ����?         ���������?    ����WUUVUU�����?    <    ��������?    ��﫪�    ������?         ����������    ��뫪�? 𯪪����         ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �m��� ���� �������������������������0������?����� �������������l �m �n �,� �� �-�P�s��#�� �������
������������L�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  ��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                ��<� ��<�<��   �� ��� �� �       ���        ������                ������       ������     ������            �?�?                                                                                                                                                                        <<�������?�  ��:�:�:�:�3 �w=��\=�5  0  <<��W�W�\5��<?��������<����.�;��;��PT�W�_�_�WTP<0���?��?��?�0��?���������?����W�����W����??���?��?���0000��������?�?�����0������0��?�������?0<<?�    ?�<<0����Ƅ��F���؅uvwxyz{|}�lmnopqrstuvwxyz{|}�cdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}�Z[\]^_`abcdefghijklmnopqrstuvwxyz{|}��08@HPX`hp�$,4<DLT\dlt|����  0@P`p���@��������@  0@P`p@�  0@P`@  0@P`p������������������������������������PRESSaSTART$TOaPLAY$LEVELaSELECT$PRIMARY$MIDDLE$ADVANCED$MISSION$C$O$M$P$L$E$T$I$N$A$G$V$R$bbbbbbbbbb$baREWARDab$MISSIONaaCOMPLETE$BONUS$TOTAL$BANK$BEFOREHEADaCOMPLETE$eeeeeeeeeeheeeeeeeee$MUNITIONSafEQUIPMENT$eeeeeeeeeegeeeeeeeee$GUN$MISSILE$FUEL$FUELTANK$ARMOUR$SELF$GENERAL$ADVANCER$SPECIAL$SMALL$MEDIUM$BIG$LIGHT$HEAVY$eeeeeeeeeeieeeeeeeee$eeeeeeeeeeeeeeeeeeee$WIN$RESULT$dddddddd$COMPLETE$HITaFIGHTER$HITaTANK$HITaWARSHIP$APPRAISE$SCORE$ENTERaSIGNATURE$CONTINUE$END$COST$�'�/�<�D�K�T�\�^�`�b�d�f�h�j�^�l�f�^�`�r�n�f�p�t�v���v�������������Ç؇����������^�#�s�(�0�9�A�G�N�R�X���������������ƈψՈ &���
Tf	Qamy(
2222222222222222
22

&
.>JXdt� 
  " *2 :B JR Zb j r zFIRST$SECOND$THIRD$FOURTH$FIFTH$SIXTH$SEVENTH$EIGHTH$NINTH$���������� �(daENEMYaaFIGHTERa$aaENEMYaaaTANKaa$aENEMYaaWARSHIPa$ORDNANCEaFACTORY$<�M�^�<�M�^�<�^�o�P0 P0�)�)�)P     000�P�B ��A � ��d�B ��A � ��`�W � � ��3  8�l �iP�l �m i �m �n i �n ة��B ��A �n  (��A �m  (��A �l  (� ���W �W �0���� `� � �� �0��� �� i� � ��
�A �F�B � ���A �  (�X  ���X �X ���`�H�Q � �	�� �a��Q �R � ���R h�`Hک �� �� �� ���Q � ��� �R � ��� �h`H�� 


m� m� �� h`� �> ��? �� ��L�� �L���� �� �� �� �� ��  ͋�� �� �>�D �� �� �� �� �� �� ΅  ͋�� ��+�� �� �� �>�C � �  ͋�� �� �� �� �>�E L���� �>�E �� �� � �  ͋�� �� �� �� �>�C L���� �� �� �� �� �� ��  f��� ��  ͋�� �� �>�D �� ʎ� �� �� �� �� ��  f��� ��  ͋�� �� �>�C �� 莋 �� �� �� �� ��  f��� ��  ͋�� �� �>�E L���� �� �� �� �� �� ��  f��� ��  ͋�� �� �>�D �� 莇 �� �� �� �� ��  f��� ��  ͋�� �� �>�C �� ʎ� �� �� �� �� ��  f��� ��  ͋�� �� �>�E  ��`� �͆�[ �φ�] �ц�e �͆�\ �φ�^ �ц�f ��� � �� �[�� �]�C �eȭ� �[�� �]�D �eȭ� �[�� �]�E �e`H�Z�� �� �� �� �� �� �� �� �� ���< ��= � � �<��@��� �eZ�I ��>� �z�!z r��� ����[�A �]�B  � ʏ �� j��̢ ��z�h`�Z� ��.�� � � �
�����_ ȹ���` � �_�I �
� �Ȁ��ҩ��� �� z�`� �� �� ����� �
�����a �ņ�c ����_ ȹ���b �ņ�d ����` `Z ��� �A �� �a�B �� �c�I �J �_΄ �� � 0D΅ �� � 0:�J �8�
�H �>�G �H �>�G �!�� �� �� �� ��� �a�� �c�H �_�J ���A �� �B �� �I �J � �� �	D� �� �:�J �i
�H �>�G �H �>�G �!�� �� �� �� ��H �_�J �� �a�� �c���� �� �� �� �� �� z`Z ��� �A �� �a�B �� �c�I �J �_� �� �	D΅ �� � 0:�J �8��H �>�G �H �>�G �!�� �� �� �� ��� �a�� �c�H �_�J ���A �� �B �� �I �J ΄ �� � 0D� �� �:�J �i�H �>�G �H �>�G �!�� �� �� �� ��H �_�J �� �a�� �c���� �� �� �� �� �� z`Z ��� �A �� �a�B �� �c�I �J �_΄ �� � 04�J �>�G �J ��H �>�G ��� �� �� �� ��� �a�B �c�H �_�­A �� �I �J � �� �	4�J �>�G �J ȌH �>�G ��� �� �� �� ��H �_�� �a�B �c�¬� �� �� �� �� �� z`Z ��� �A �� �a�B �� �c�I �J �_΅ �� � 0:�J �8�	�H �>�G �H �>�G �!�� �� �� �� ��A �a�� �c�H �_�J ���B �� �I �J � �� �:�J �i	�H �>�G �H �>�G �!�� �� �� �� ��H �_�J �� �a�� �c���� �� �� �� �� �� z`xH��� ��� �� ��  �魓 ��� ���� hX`H�Z�� � �� ��B� ���K � �N  ���K �K � �� ����N  �� �� ��ة�3  8� Z����N  ��z�h`��A �
�B �  (꩑�B ��A ��  (��A ��  (��A �n  (��A �m  (��A �l  (�`� �G �� � ��G �G �0�LY��� �� �H �
�����a �ņ�c ȹ���b �ņ�d �H �a�� �c��  ���H �H � �L
�`� �G �J �� � ��G �G �0�L.��� �� �H �H � �� �� �H m� �� mo �o �H �mH mH ml �l �m i �m �n i �n �H m� �� �� i �� ؘ
�����a �ņ�c ȹ���b �ņ�d �H �H �a�� �c�� �J �� �[�� �] ͋� �> ��? �� �e�� �>�J �H �H � �Li�`�V �j ��V �!��� �9��� �Q��� �V ȹ!��� �9��� �Q��� ��� �	�� ���  ���� �� �� �� �� �� ��� ���  ���V � �� `�� �F �F ��E �D �F �D 0U�D ���]�G ȱ]�J �G ;�G �]��J �]�[�G �e�H ȱ[�I �e�J �G �[�H �e��I �[�J �e�D �E �D ���E �E �F � Ў`� �e�x��̢ 0����� �� �� � �� �G�� �� �	� ͋�� �K �>� �� �� �� ��΅ �� � 0� ͋�� �>�K �>� �� �>�K ��`� �� � ��  ͋�� �>��  ��� �� �0�� �� �	0�`xH�Z�� �G � �� H��3� �/����' Y��� � �R ��� � �H�G ��  �h��  ��L6��0� ��  E��� � �" ���� � ��G ��  �h�0� ��  U���G �� hz�hX`Hڮ� �� �� �� �� ��  ���h`�� �� �� �� �� � �� �΄ �� ��  �魎 �� �� ��  �魎 �� �� � �΄ �� �� ��  ��`�� �� �� �� �� ��� �΅ �� ��  �魏 �� �� ��΅ �� �� ��  �魏 �� �� ��  ��`xH�� � � U���� ������ U�hX`xH�N H� �N  ��h�N hX`��B ��A � �N � ����N �B ��A � �� ~�B �<�թ|�B ��A � �N � ����N �B ��A � �� ~�B �<� ���)��&  ��` ���A ��B � ���A �;�B � ���A �N�B �	 ��`�@ �����< ����= ��G �B ����> ����? �A �<Q>�>�< Ȳ<Q>�>�< ��G ��`�h ��� �0�A �d�B  �� �� �	�A i�A ��`�
�B ��A � �驇�B ��A � ���A � �� ��`HZ� �> ��? � �>� �	��	0�� ����� zh`Hh�|�B ��A � ���A �X�B � ���A �d�B � ��0�H �X�I  �`��g � �h � �Q �R �� �� �V �� �� �l �m �n �r �s �t �u �v �w �x �y �z �
�j `�� �� �o � �� �� �� �< ��= � � �<�������� ��`�� �� � �> ��? �� �� � 0+ ͋�� �>� ��� �����΄ � 0 ͋�� �>� �	� � 홀���� `�� �� � �> ��? �� �� �	/ ͋�� �>� �#�� �� ���� �	 ͋�� �>� ����� � 홍� `�� 8�	��>� ��� i	��>� ����� `�� �� �� �� � �> ��?  ͋�� �>� ��� � ���΅  ͋�� �>� ����� � ���� `�� �� � �> ��? �� ��  ͋�� �>� �%�� � �"���  ͋�� �>� ��� ����� �
�� �� ���� `�� ��>� ��� ȱ>� ����� `�� HΎ �� �G  E��� ���h�� �h��  ��G ��  ��`�� H� �� �G  ���� ���h�� �h��  ��G ��  ��`xH�Z�� H� �� �G  Y��� ���h�� ���h��  ��G ��  ��� �� z�hX`�D H�E H�� �� � �� �G  �� � �$�� �� � �N  ����N �G �� ��  �� j�ɩ �3  8 �� h�E h�D ` ͋�� �>� ��� ����� � �� `�P�B ��A � ��d�B ��A � ��s�B ��A � �驂�B ��A � ��`� ��������������������������3 ��%��������������������P��
����
����������=�����������������������������������
������ ����� 轱��� ����� ���ԍ���
����


m���� ���`Hڭ8��A �9��B ��
��&��L �&��M  �� �̩ z��  ��g �̩�A �2�B �d�@ �  \��  ��I �������A ����B ʽ���L 轀��M  �� �̭:��A �;��B ����� (� �� �� �� ���h`Hڢ� z� ������ �� ���h`Hڢ� z� �� ������ �� �� � ���h`H��������&8��������8����m i�m �n i �n �Э��8����m i �m �n i �n ����8����m i0�m �n i �n ����h`H�Z��  |ϩ2�P �� ͩР��������P�<��P��P�s�s)�խ� ��
 4ө�s�ĩ�A �N�B �= �  )��� �� �� ��z�h`H� �@ �
�A �S�B ��G �/�H  M�h`H���Q �Q � |ϭP8�Q �P��G �Q �H �  A� ���Q � z�� z�� z�� z�h`Hڽ� �	0� [��h`ڢ�s)�ɀ0 ӭ�� ��s)��s�
����#�����`Hک���� � ���	��J�� ���h`H�Z�
�����A 轉��B �
�����L ����M  ��z�h`� � � � � � � � � � � �( �) �* `Hڜr �s �t �u �v �w �x �y �z � �^�� �&����$�� �&�h`� �Q ���`H�Z�� z� �� ������ �� �� v� �� ���"�� o�� � �� �̭  ��� Y�z�h`H� �A �B �(�G ���H � �@  M�h`H���%��A �J�B �b�@  \���i��� �����p� �=��A �d�B �b�@  \�� �����������G���i`����i ��������!�"��A �t�B �b�@  \����m�i��؀	�"� �� V��h`H�Z��A ���B �b�@  \��a�@ � \������A � ����� �� �ʀ�z�h`Hک ����� �� �ʀ��h`H�Z�������N8��������8�����A �t�B �a�@ � \������A  V���i����i �� ���������z�h`H�Z���)�JJJJ�@ �����a�@ ����� \��)�@ ��������a�@ ����� \�z�h`H�Z���)�JJJJ�@ ��������� \��)�@ ������������ \�z�h`xH�Z�@ �a��$�>�b��%�6�c��&�.�d��-�&�e��(��f��)��g��*��h��+��i��,�����< ����= ��G �B ����> ����? �A �<-N �>�< Ȳ<-N �>�< ��G ���A �A z�hX`H�
�����L ����M  ���h`HZ��3  8� B� �� (� �̈��zh`Hڭ��@ �-�A �P�B  \��h`H�a�@ �-�A �P�B  \�h`H��A �f�@  \�h`H�b�@  \�h`�Z�P��������z�`HڽPm��P�h`HڽP8��P�h`H�Z� �L�$�0�a�#�b��c��d��e��f��g��h��i�8�7�@  \�Ȁ�z�h`H�Z��1 |� Hԩ�-�"�P�c�� Y��"��/� z��"��.��J� Y���1��"�B  R���A �"�B �����1�
���2��3 �2�B  R���A �2�B �� С�B�B  R���A �B�B �������@  E�  (�A������
���������m������ � ��� ����i���؍� С�R�B  R���A �R�B �����4�
���5��6 �b�B  R���A �b�B �����7�
���8��3 � e���A ���B �H ��A ���B ���@ ��G ��H  M� 5��  (� t��  ���� �) ��P�r�� 
�L%��)�'����������i������N�)����0��2������. B��)��Pi�t��"�P�)��P8��"��r�PLO��P�"� �L��2� %�L��B� ��L��R� �L��b� !�L�LO� �� �� �� ��z�h`��A ���B � �@ ��G �	�H  M�`��A �a�@ � E���`H�Z����� 3ԭ2�� �� ��� � �Ȁ��2�����z�h`H�Z��2 |Ϡ � t� t� �� t����� J�� ��ε �ީ���� 3ԭ2�&� �� ���2�����z�h`H�Z����L!��ͩ���"�B  R� 5����/��A �"�B �2 ��A ���B  i���@  E�  (� (�Lo��а��A �"�B �3 ��A ���B  i���@  E�  (� (�  ���� �) �W�)����	���L!��L���)��L�� B��)��Pi�t��"�PL!��)Ь�P8��"��r�PL!����"�����8���� � 
������L!���������8���� � 
������z�h`H�Z��ə�L���2�B  R� 5����/��A �2�B � (��A ���B  i���@  E�  (� (�Lը�� �/��A �2�B �  (��A ���B  i���@  E�  (� (�Lը��A �2�B �0 (��A ���B  i���@  E�  (� (�  ���� �) �u�)���0���L2���i��L2��)�����0�L2���8���L2� B��)��Pi�t��"�PL���)Ў�P8��"��r�PL�����3��ə�)����"�8���� � 
���ɐ��i�L������L��� �1��ə������8���� � 
���ɀ��i ؀�������0�/��ə𽭞����8���� � 
����p��i0؀����z�h`H�Z�����L㫩B�B  R� 5����,��A �B�B ��@  E��A ���B  i��P (�  (�L����/��A �B�B � (��A ���B  i���@  E�  (� (�L����A �B�B �2 (��A ���B  i���@  E�  (� (�  ���� �) �|�)���2���L���m��L��)�#����2�L�����L���L� B��)��Pi�t��"�PL㫘)Ї�P8��"��r�PL㫭��A�����6���P����*���8�P����� ��� � 
���i�������L���0����������8���� � 
���i����������2�.����𽭞����8���� � 
���i�������z�h`H�Z����L�������R�B  R� 5����/��A �R�B �5 ��A ���B  i���@  E�  (� (�Li���A �R�B �6 ��A ���B  i���@  E�  (� (�  ���� �) �c�)����	���L��i�L���)��8��L�� B��)��Pi�t��"�PL��)Р�P8��"��r�PL���������8���� � 
����L���������8���� � 
����z�h`H�Z����LK�������b�B  R� 5����/��A �b�B �8 ��A ���B  i���@  E�  (� (�L����A �b�B �3 ��A ���B  i���@  E�  (� (�  ���� �) �W�)����	���LK��L.��)��L.� B��)��Pi�t��"�PLK��)Ь�P8��"��r�PLK���������8���� � 
����LK���������8���� � 
����z�h`xH�Z��
��G��< �G��= ���H ���I �B ����> ����? �A �<�>�< i�< �= i �= ��H �H � ����H ��I �I � ��z�hX`H� �N  O����N h`H� ��������� ���������B ���A  O����q� t�����������ة��������������B ���A � �������� O��������B ���A ���������� O����D0 t��������������� t����B ������A � �������� ����i���A  O������8����A ������ O����� t���h` ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?   ?��������?�?   ?����������?   ?��� ����?   ?��� ����?   ?��� ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                                  `% Z	�V*�Z� P �
P�@�Z     <          <          <          <          <         ��        ��        ��?      ������?    ������?  ���������������������    ��        ��         �         <        <        <        <        �       ��      ��     �����   ������? ���������   ��       �       <      <      <      <      �     ��    ��   ����? �������   �     <    <    <    <    �   ��? �����  <        �� ��?� � �?�       �   �  �   �?  �������   ������  ���������������  �����+            �   0  ��g �0�H �X�I  � �� ~����
�����/�� �N  ���N �g �g �0��g �X�I ��d�I  ꀿ`.
� �
� �
� �
� �� �
� �
� ��.
� �
� �
� �
�    �� �
� �
� �� �� �
� �
� �
� �
� �<� ��    �� q� �
�    �
� �� �
� �
� ��.� �
� �
� �
� �
� �
� �
� �<�   \�����\�\���������.�}�.� �� �� �� �� �� ��.�   }�\���\���������\�����   H�Z� �> ��? �� �0� �� 
�����< 轀��= � �C �<�G �����C �<��G �>�C �C �� ��z�h`H�Z�g � �H �d�I  ���   ���d���.� �N  ���N � �g ��g �I 8��I �˩�g ���I ������� �N  ���N �g ���g �I i�I ��� �g �d�I ��� �������g � �����	�����������	����n z�h` ?� ?� ?
� ?
� ?
� G
� O� G
� T
� O
�    ?
� (� G� G� G
� G
� G
� O
� T� O
�    T
� _
� �
� (� 
� _
� T
� O
�    ?
� G
� ;
� ?
� /
� /� /� /
� 5
� ;
� ?
� � G
� ;
� ?
� /
� ;
� /� 5� ?
�    
� G
� ;
� ?
� O
� ?
� T
� ?
� _P�    
� �
� 
� �
� 
�
� 
�@
� 
�
� �
�@
� 
� �
� 
� �
� 
�
� 
�
� 
�@
� 
�T
�    
� �
�}
�T
� 
� �
� 
� �
�}
� 
� �
� 
�}
�    
� �
� 
�}
� 
�@
� 
�@
� 
�@
� 
�T
� 
� �
� 
�
� 
�}
� 
�T
� 
�    �
� 
� �
� 
� �
� 
�T
� �
� �
� �
� �
� �� ��    �	� �	� �	� �	� �	� �	� �	� �	� 	� �	� �	� �	� �	� �	� �	� �	� �H�   }	�.	��	�.	��	��	�}	�.	��	�}	�T	�@	�.	�	�	� �	�}H�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ���ة��  ��� � �T � � �U � �ߍ& ����"  ��� t ����< ��= �� � �<����= ��� ��XL �H�Z� ����#L���O �Q � ��Q �g ��S�R � �L�R �G�O ������λ�����������=�� �� �ڭ�������� ��� ��(z�h@H�Z�' )�D� ��4�����% m� [����͵� Bڜ������ �����S �# �	�O �S �# �$ �% z�hX@                                                                                                                                                                                                                 ���N  �� ɮ��3  8� ��� �� �� O�L �L �� O� ��� O�L �� O� �� O�L �� O� ��L�� Ș��7  �� �� � �� �� 8��7  �� O�L �� O� :��g �� �� /� ���� ���LE� ���� ���Lí� ��� 3��ڭ  ���� ��� ��L��� %�L��ɿ�L�����	 �� ͚L�����	 �� ��L�����# �� )��� ���5 j�  ����L�� �� )�L�����	 �� ;�L�������3  8� ��L�© �3  8� � � [��� � � f��� ���9 �L�� �� � �� ��g ���o �d0� ׊ ;�Lk­� ����o �xе���7  �� /� ��� O�L`�� O�ߍ& �l �m �n �� �� �k �� ��L�Lk©�3  8�` ᛩ�7  �� �� �� 8��7  ��ߍ&  Ο ��ߍ& �  O�L �� O�<�S  �Ω�� oΩ�  |ϭ�ɠ� Uʀ d� ������ �� ��X�S �#  ������& ��ɠ� �έ��� �Ω��������� �� �� �ҭ�ɠ� x� �� � �� (� S� �΀
������������" �� �� �ҭ�ɠ� �� � �� (� S�L�ŭ����L�� �ϭ����������  ���	������L�Ŋ�� ��L��2x���& � � �*  � �̭  ��� �X���& � �N ���N Ljĭ�ɠ���� �̩����)� �Ɗ)� EǊ)� �Ǌ)� �ǭ���)� �ȩ
������) � Wȩ8�
���� ?٭�����ɠ�
���� �� i� Tح���Ljĩߍ& � ��x ������� Lĩ�A �<�B �F ��A �X�B �G ��-�<�P�c���  (��  ���� � B��)��,�)��P�<��X��<�P�)�ϭP�<��X��<�P�� 
� ��P�<��LĜ ��L©ߍ& � ��x ��� ����� ���� L"�� H� ��L©�� �  �� �`� � �  �� ��`H�Z��ɠ���I�"�-�@�-�N�8 �������� �� ���2�� �	�2��4��  ^��#��-����-z�h`H�Z��ɠ0��I�"�-��@�-�N�8 �������� �� ����� �	�����  ^��#��-�0���-z�h`H�Z��ɠ���H�"�Pɇ�?i�P�qi�q�.��� �� �������5�P ^��#��P�Ai�Pz�h`H�Z��ɠ���H�"�P�2�?8��P�q8��q�.��� �� ���9����U�P ^��#��P�!08��Pz�h`Hڭ�ͩ�; W����4�  d����ɠ��@� �ɀ����ɠ��( iπ ����h`H����'���"� d��ɠ� #ɀ y�����8����h`H� �������������� ������ �h`H� �����$������ �ʽ���������� �����-�h`H�Z a��#��� �2� @��!� *��!� @��!������ ����8 i�z�h`H��� �	�s)��0���#��h`Hڢ"�-����� �(���#����� ������ ������ ʜ�� ���h`��� � �s)�ɀ0�-����m�8�0�0	��#�֩ ���`H�/����� .�h`H������ .�h`H�'��� �� .�h`H�&����� .�h`H�Z W������� |Ϡ"�-m��-�P�Pz�h`��! |ϩ�" |�`��! |ϩ�" |ϩ i�`Hک��@ ���G ���A  �ʭ�i�A ��G ���@ � �� ���h`�qi�B ��H  M�`H�Z���@ �8����G �m��A  ��z�h`H�#�A �ri�B �� _�h`H�
�A �ri�B �� _�h`H��A �ri&�B �� _�h`H��A �ri&�B �� _̩"�A �ri&�B �� _�h`Hڭ�ɠ�I��� �=�i�9�P�n�2 �˽-��%��!�Pɉ�Ɍ����	8�

��� ��� ����!й�h`�-��.��*�PɄ�#ɒ�����
���8���3  8��`H�Z�-8�������A �;��G �P�B �����I ���B ����> ����? �A �G �H ���
.��H �����>�>ȭ�>�>�I �I ���������A �B ��z�h`Hڪ��G �)�JJJJ z̊) z��h`xH�Z�����< ����= �G �J �B ����> ����? �A �<�>�< Ȳ<�>�< ��J ���A �A z�hX`H�Z����� ���  �� ���� ��z�h`H�  )@��h`H�Z������� ���� ��z�h`xH�Z �ͽ3��H ����G �ɀ� �̀ ��  β<-N �> ����B �H ��z�hX`xH�Z�� �ͽ���G �G 8�G �J �3��H �H ���� ����� ��L�ͭ�ɀ� �̀ ��  β<>�> ����< mJ �< �= i �= �B �H ��z�hX`�)�����	�)���`�-�A �P�B �� �ʊ`8�
�����< ��� �͍= `
�����< ��� �͍= `�G �I �B ����> ����? �A `�< i�< �= i �= ��I `H�Z  β<-N �> ����B �H ��z�h`H�Z  έ@ -N �>��I 0
���B �H ��z�h`Hک � �� ��#���h`Hک � �������h`H�Z�����> ����? � � �>��(����m��z�h`H� �@  *� M�h`H�Z� ����> ����? � � �>��(����P��z�h`Hڭ���	� ������ ��h`H�Z�����> ����? � �>	��>��(0���m��z�h`Hڽ-�A �P�B �� �ʽ���G �(8�A �G �G �3��H �8�B �H ��H �h`H�Z� W����� ��z�h`H�Z� ��z�h`�c��� ����-����P���s`H�Z� ��ɠ�l��)��1�� ��  �)� mЭ� Њ)� �Э� =Њ)� �Э��� ���J�P�)� �Э��� ���J�P���%��z�h`HZ�� �4��5��2�
�2��3���� zh`HZ�� ������
������� zh`��� ����#��`� ^��#��-�0���-� �`� ^��#��-����-� �` ^��#��P�608��P� ` ^��#��P�2�i�P� `Hڢ �� �� =р ���h`H�Z��U�@ � �A �(�G ������ ����H ���m��B �� M�������� ����@ ����'�ˢ:��z�h`H�� ������
������������� �������������������G  �рD�2���������3����������4��������
��������G  �h`H�Z�P�������m�,�B � �A ���
��� z̈���� z����mG ����z�h`HڽP���(�����m�0�B ��8����A �� z̭A �(��� z̀�mG �����h`H���������h`Hڢ �� ��J�ޯ ��� �h`����������� `Z ������� �� ���� =Ѐ Щ��� z`H�x��� �C�!0���� � x� �ʀ,��ɠ��P�n��s)�ɐ��������n� 3ԩ����#гX�h`Hڽ� � �νs)� �� 4��h`H�Z���� �����������c���ʽ������ �����	������<�(8�-͚01��͚08�J���-8��-���8�J}-�(��'�-������ ���sz�h`H�Z�� �Ԫ���G ���8�P�H �� �ʽ3��H ��H z�h`Hڽ� �ʽ��8�G ���ɀ�8�
����m��< ���i  �͍= �
����m��< ���i  �͍= �h`H ����� �Ӏ *� A�h`H�Z���-�. �����'�sɀ� )����
��� �Ԁ�� �ʽ������ ��z�h`Hڽ� �� ������ � �����������������h`ڽ� � ���	���������`H�Z�s)��� �c��� �Χ�C���s�s�� �(� *��!� rՀ'�s��-� @��!��s��-8�P��P� ^�z�h`��� ���-����!��`��� ���-����!��`�D ��8�-���
0 ր�- ��`�% ��8�-���
0 ր�- ��`8�� �������
�������s)m��� ^й-`8�� 

��ΙΙ�s)m����-`�P���� ����i���P8����� �8�P��P` ��-m��-`ڭ���� ��*͙�������`�, ��i��8�-����
0 �ր�- ��`�= �Ս�8�-����
0 �ր�- ��` �8�-��-`�Z���P�P�����ʽ3������}P͚�L���ʽ3�yP���P�7�-�-�����ʽ����}-͚����ʽ��y-���-����� z�`H�Z�� ����� ����s)�ɀ� �����Χ �� Z׀��!��z�h` ٹ-m��- �ٹPm��P`ڹ� ����ɠ��?��P�F��?��7���� �ʽ��s� d� ?��`� �� �s)�ɠ����
���ɐ�$�-���i����i ��؀���i��؀���i��عs)�����)�͚���



͚����i��ح�ͫ�����`H�Z�� ����� �*���s)�ɠ�ɰ������� �����Ψ �� Z׀��!��z�h`Hڢ��ɠ�T�� �H�s)�� �(�0�; ׽� �3�s)�
� �� Χ�"�s�P�P� ؽ� ��s)�� �� Ψ��!Ю�/�� �%�s)�� ��0� ׽� � �Ԁ ؽ� � ����!���h`H�Z�s)��� �c��� �Ψ��	 �s�� �2� VՀ 9��sz�h`H�Z�����������ݣ�08���J��z�h`Hڢ�� ��� �� ��!���h`ڢ �� ���!������`H�Z��ɠ�W��� �K�s)�ɀ�B �����; W����9���� |Ϲ� �� ��-m��(��- ���Pm��P�� �� ��!Ыz�h`�-�0�%�P�0�i���`H�Z������3�����3�08�3�J��z�h`Hڜ���� �%�s)�ɀ0����)�͘���



͘����!���h`H�Zζ���� 	ڭ���W W����P����ҍ��(��O JJJ���"������O JJJi���h |ϭ��P���-��������� �ԍ�z�h`H���������������	�� Mۀ =ۀ -��h`H��������;���� ������������)������� ���O )i��O )?i��h`H�G������ q�h`H�S������ q�h`H�����M���Ѝ� qۀJ� =ۀ -�h`H�Z������O���J���� 	ڭ���: W����3��� |ϭ���i)�P�O JJJ���"�-)����m���� ��z�h`H�Z������������� �L�� HԽs)��`� M�L��ɀ0| ��ɰ�� ��<��� &�3ɠ� �� �݀'��� �� ��������
����ɐ���� �ܽ� ��+���&�s)� 4ӽ� ��� ������� ��� �� �s��!�L�ۭ�����������	������z�h`H��

m�'��&�	h`H�Z �������-�� ��z�h`H�Z qݭ��� �� �� �>�
J� 1ݭ�ɠ�+�����#�8��}P�P���8�����P8��P�Pz�h`��J��  �)��-��)��-`Hڽs)��s�� J�ޯ �
�� �� �� �h`H�Z��ɠ��P�m��0��Pɝ�	�0 ���� �� z�h`H�Z�P�� ���� �� z�h`�-�'�� � ����������	� ��� ���`H�Z qݽ� ��y�y�Ɂ�ɉ� iހh�z�ɂ�Ɋ� }ހT�{� A߀KɃ� �߀Bɋ� n�9�|� G߀0Ʉ� �߀'Ɍ� t��}� M߀Ʌ� ��ɍ� z� � m�z�h`HڽP���P��P�h`H��P�h`H�Z�O )i���O )i����s)�d���L=߬  �)��)��-͘��-�%��-�
�-���-�)��Pɖ��)��Pɀ��P͙��Pɛ�@�P�;�P�6���
���s�%��-��� ��%�-�`�P�� ����s H�z�h`H h�h`H h�h`Hڭ  )��P�P��J�� h��h`H�Z�  �)� ���P��J��	�-��-��-��-� H� ��z�h`��	�� 8��� `��	�� i�� `H��ɠ� ��2�� ,���2�� W�h`H��ɠ� ���� ,�� ������A�� W�h`Hڭ�ɠ� ��P�� ,�� ������P�� W��h`H�Z�Pͼ��P��  )��� Ƀ�Ʉ����Pz�h`H�Z�J�B�"�P�P��P�P��P��)�-�-�!��-� �Ȁ�-��-� H� �Ȁ�-�Pͼ��Pz�h`H�Z�  �)�
���" �߀�)�
���% �߀ �J�-�-�	�%0�-� H� �Ȁ�-��-� �Ȁ�'��-z�h`Hڭ�ɠ� 3�P���  )��P��P��P�h`H�Z�  �)��)��-�	��-� H� �Ȁ�-��-� �Ȁ�-z�h`H ��h`H ��h`Hڭ  )��P�P��J�� ���h`H�Z�  �)� ���P��J��	�-��-��-��-� ��z�h`H�Z �ݽ� �L���f�� ����n�	�v�� �� �������L���e�� ����m�	�u�� �� �������L���d� 5�w�l� ]�n�t� {�e�c� L�\�k� 2�S�s� ��J�b� c�A�j� �8�r� ��/�a�� ����i�	�q�� ����ɠ��i��  ������� m�z�h`H�Z��ɠ�G�P�n� �ހC�-� HԽ-��� � �Ȁ�-��!��-� ��P���P��P��Z�� ��z�h`H�Z��ɠ� ��K�� �� ������K�� ��z�h`H�Z��ɠ� ���� �� ������<�� ��z�h`H�Z��ɠ� ��-�� ���-�� ��z�h`H�Z��ɠ� ���� ����� ��z�h`H�Z��ɠ� ���� ����� ��z�h`H�Z�Pͼ��P��Pz�h`H�Z�J�B�"�P�P��P�P��P��)�-�-�!��-� �Ȁ�-��-� H� �Ȁ�-�Pͼ��Pz�h`H�-����ɠ� �� ��h`H�<����ɠ� �� ��h`H�����ɠ� �� ��h`H�-����ɠ� 3� ��h`H�����ɠ� 3� ��h`H�K����ɠ� 3� ��h`�Z�� ���� ���" ��� ��?�� �O�-�r�P� d����z�`H�Z�  �)���� ���P��J��	�-��-��-��-� H� ��z�h`H�Z�  �)���� ���P��J��	�-��-��-��-� ��z�h`H�Z���L�孢


���O )m���������)m������� 	ڭ���M W����F��� �w���ɠ�:����� �-i�(��'�-�Pi�P�� ʭ�ɠ���i����s��z�h`H�Z�

m�$��!��


m�i��P� qݽ� �L����J�s)�	�H�-m��
�'�-8����Pm����P8��d� c�L��s)�� �L���ɠ�I�� �� 1ݬ  �)��)��J��-���-��-�� ��
�)��)�4�P��,�P�1�s)�%�� ���� ���" ��� � p��P�P�P�� �� z�h`Hڽ-���-��-�P�<��P��P�h`H�Z �ݽ� ���+�s)��� ���" ��� � p��P�P�P�� �� z�h`Hک ��  ���h`H� �筣��?��_�� �O�-�r�P�a�s�h`Hڭ�ɠ�������8����� ���������h`H�������8����`��8����h`H�����JJ���������������h`H�O �  ����O �0�h`H�  ����h`�Z �� ���)��&  �  ��� � �� �ߍ& z�`Hڪ�C�




�I ��)I �& �h`�Z� ���� ���� ��z�`�Z�P���� ���� ��z�`�Z������ ���� ��z�`H�Z�/���� ���� ��z�h`H�Z�� 
��K��< �K�m��=  ��z�h`�E JJ�F �B ����> ����? �A JJ��<-N �>�< i�< �= i �= ��F ����D ��`xH�Z�< H�= H�> H�? H�A i�E �B i�D �h ��� ����	�
�����m� ��ӆ�< ����=  ��h�? h�> h�= h�< z�hX`xHڮ� ����A �� ����B  ��hX`H�Z
����L ���M � �L�$��a��[��d�8�7�@  E�Ȁ�z�h`H�Z�< �@�= � � � �<����= ���z�h`ڭ  ���� ��`�H �A i�E �I �B i�D ���  ��`H�Z�)�JJJJ�@  E�)�@  E�z�h`xH�Z�< H�= H�> H�? H�@ �[��%��a��$��d��&�����< ����= ��G �B ����> ����? �A �<-N �>�< Ȳ<-N �>�< ��G ���A �A h�? h�> h�= h�< z�hX` �Ɯ � � � � � � � �- �. �ߍ& `H�Z� ���Q� ���.� � �� � � �  �� � �� � � �  �� � �	 � ��� � � � Y� ���.�( � �� ��! �" � � � �  s��( �( �# � ��(z�h`� �� ȱ� ȱ�	 ȱ�
 ȱ� )
��L�� �L�� Ȍ � � �	 � �'� �/� ȱ/� � �� � �� ��Ȍ � ��`� ��! ȱ�" ȱ�# ȱ�$ ȱ�% )
��L��& �L��' Ȍ �( �) �# � �#� �  �� �� � � � � � � � `� �� ȱ� ȱ� ȱ� ȱ� )
��L�� �L�� Ȍ � � � � �'� �1� ȱ1� � �� � �� ��Ȍ � ��`H�Z�
 )?	@�+ �
 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �- �� �- z�h`H�Z� )?	@�+ � 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �. �� �. z�h`H�Z�$ )?	@�+ �$ 4��-+ �+ �) �&��% )@��J��+ �+ Ȍ) �&����) �% �) �+ � �- � �. z�h`� �- `� �. `H�Z�7 

����/ ȹ��0 ȹ��1 ȹ��2 � �/� �1� ȱ/� �1� � � �� �  �� Y� �� ��� z�h`H�Z�3 
��8�� �8��  � ��*  �� s��� z�h`Hڪ�5 ���9 ����5 �9 ���8 �h`H�Z�8 ���C�5 
��n��: �n��; �9 

��:�$�* ȱ:



�4 �6 ȱ:�) ȱ:4 �( �9 � ��z�h`�8 �* ` �� �� �� �� �� �� � �� �� � �� ��    �� �� �� �� _� d� q� � �� �� ��    �� �� �0�    � �� �� � �� �� � q� � �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��    �� �� �� � � q� � �� �� �� �� �� �� �� �� �� ��    �� �� � � q� � �� �� �� �� �� �� �� �� �� �`�   \���\���\�����\���:�\�������\�:�������   }���}0�\���\����0��0���\�������\��0���\��0�   ��\��0��0��0��`�    /�  ,�  *�     G� C� q� K� O� �� Y� G� 5�    2� /� .� ,� *� .� %� .� *� &�    ��    �� �� �� ��� ��� �� �� �� � d�    �� /2�   .� �� �� �� ���.��@���� �� �� �� ���� �� ��� ��   @�.� �� �� �� ���.� �� �� ��   � ��� �� �� ��� ��@�.� �   \���\���\���\�������\��������\���   \������\���\��������\���\�\�    �    �� �� �� �� �    �� /2�   	

	�	�	�		�		��
 �

		�
	��
	�
�
�
	�	�	�

		��������
���&�0�4�������U�g���:�  ������Q�  =����  �p�  ;�z���ƴ  
�l�  ����J���  �\����  P�  ��  r�������0������  �������"�%�2�X�c�f�q�z��������t�}���  

 +.148<AGMSZahpx�����+036:>DJPW^elt|����-037;?EKQX_fnv~����/259=BHNU\cjrz�����    ���������������������������������������������������������������������������������������������������������������������������������������1�G�_�w��������$�<�S�k�����
 �� 
 ���  ��� 
 ��� 

 ��� 
	 ���� 	

 ��� 	
 �� 	
 �� 
2->:64(<20(6<&.40*3:"6.,(&0,*$.,!($/"'"$ ($"
	
           	
   !"#$% '()*+,   012345 789:;<= ?@ABCD   HIJKL NOPQR TUVW YZ[\  _`abcdef  ijklmn  qrstuv  yz{|}~  ������  ������      
          "!          





  





  





  





  





  





  ����  cB� g
 mIIUF2
2P �<diZF2 ddl_K7- dcqvvU cciZF2 cci_K7- 2<FPZ 2<FPZ 2<FP 2<FP    ��nZF2  ��nZF2  ��nZF2  2FZn�  2FZn�  2FZn�    ������� �RR���� �B/44444 ??!!!!!! /���� ee44444 ee!!!!!! ����� ����� ���� ����  dd������  ������  ������  ������  ������  ������    	 (($$   	    
    	
  
	  
  
  	
  
  113/  
 		3GGG	 	  
G 	  	 	
 	   !  
      
    ��������������A����
�P�x������A�B9S�U�������C�C�B�B�B@C���A�C�A�AB=BYBdB���A�AmB�B�B�B�B�B���A����������9MN�AB=BYBdB��SL�LmB�B�B�B�B�B���N�N�NO>O���O�O�O�O<P���P�P�P)Q��������������hQRR�CEK�K�I�C�C�����C~D�D0E�C�C�����C�I�JK�C�C�����CXE
H�G�FmE�����CXE�FxFFmE�����CXErII_HmE����  0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____PRESSaSTARTaBUTTON$NORMAL$FLASH$BEGINNER$AVERAGE$EXPERT$MUSICaAaBaC$GAMEaOVER$CONTINUE$END$PAUSE$LEVEL$TIME$SCORE$BLOCKS$aaaPLEASEaSELECTaa$ENTERaSIGNATURE$LEVELaSELECT$PRIMARY$MIDDLE$ADVANCED$HASHaBLOCK$EAGLEaPLAN$8�K�R�X�a�i�p�|������������������������������U  � ��Ѱ�����r#)0 PdxF<2(
F<2(
F<2(
F<2(


���<  0�� � �? <  ��   0@P`p��������  0@P`p��������  0@P`p�������������������������������������������������������U� ���