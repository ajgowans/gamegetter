      �    �[      �               �   �[[      �           �����Z  X[[      �-           �e���j��[[[    *  |7   �    �������X�[[[U  .  l'   �U	 ����������VX�[[[U ��  �)   @U `Y������k�[��[[[� �� ��� ��
 `Y�����������[[[� ��d�[�eY�� `Y�����U��[�[[[� ����Z�eY��[U����������[�[[[�WUuUB�[�eپ����۾��U�������[[[�WU�ݒ�����������������zww���[[[�WUuU�Z�e�������������ww�[�[[[�WU��mU�����������������{w�[�[[[���~U���������������zU���w���[[[��������������������^U���{���[[[{U�����������                                         �W                            �Y P              @U       �� �  �W P        �YV�U �V  �o��jV  ��      TP�jVfV�U T��V��j ��V�     @V���Z�UlfUg��Z��� ��U�V   ��կ��mf��V����j��^���Z��VU   ����k�����j��٪Z����j�����U  䪚�����֫�j��گ��������V���VZV��������֪j���j�Z�����~��V�Ze���������j���i�kU�����j����ڪ�fջvի��_ֺ����i��Z���������j���k���گ�몵������������꿮�g��������j��������������Zm�����Z���V������絛j�����j�����]��ګ�j����������UU   Z    Z  �        @U@U UU �V   ��  �      PUUTUUEU�U �fU   ��e  �      TUUUVV��WfVū�U  �jY  Z�  @UU@U�ZU�fYU������Z *�g� Z� �UUUEU��V��eU�jj�����U� Z� �UUUե��Z��j��������֗���f Z� jUe�է�j����������U����U Z��kYU�Z믪��k�������]U��yY�Z��UYW��������������뺫UU_m���Z���UW�U��������������kUU_[U�֫�֪�U]�U��������꯯�����UU�[]�Z���[�wUU髯�����������jVU�k��f������_�w믿�����������UY�����Y������}����������������[�����jf����������������������������������������������        �     �     �     �     ��   ���   �[-���V�? ��U�  �U�? �oUU� �oUU  �U�?  �U�?  ��90 ��?        0                                  �     �    ��   � ��3  ���   ��� �j������> ���f  �e���ki��?�k��� ���? �U�? ������ï��<��  < �   ��   � �   �     0     0        0   � <     0 �     �(   �� <��  ?(H * ji�   j�  JdT R�E"R$U"< �V�  BU�   *�    (�
�0��  <            �  � �  0                   �        "     *    �B
 �T �DR�TE�  TU�  V�Z �YDUH �)�VJ @�T&�  �FdF  �  �I   H�   @�                                              �   ��=   ��=   ��   �=�  ��>  ��n���um�� ���U�?���U�?�um�� ��n����>  �=�  ��   ��=   ��=    �                                        �   ��=   ��=   ��� �=�� ��>  ��n���um�� ���U�?���U�?�um�� ��n����>  �=�� ��� ��=   ��=    �                      @   T   T@   �  ��=  ��=E  ��P�=�U��> ��n��C�um��@���U����U��um��@��n��C��> �=�U��P��=E  ��=  �  T@   T    @    @   T   T@  �A ��=TU��= ����=��U��> ��n��C�um��@���U����U��um��@��n��C��> �=��U�����= ��=TU�A T@  T    @                      �?  ��?  \U�?  �s=?  ��� ? ���� ���� ��m����U�?��U����U�?��m������ ���� ��� ? �s=?  \U�?  ��?   �?                                 �?  ��?  \U�� �s=�  ���0? ���� ���� ��m����U�?��U����U�?��m������ ���� ���0? �s=�  \U�� ��?   �?                    @@U   P  �?E \�? \U�?�s=?@ ��� ?����A������m����U�7��U�W��U�7��m����������A��� ?�s=?@ \U�?\�?  �?E   P @@U       @@U   P  �?E \�? \U���s=�@ ���0?����A������m����U�7��U�W��U�7��m����������A���0?�s=�@ \U��\�?  �?E   P @@U                    �?  ��?  \U�?  �s=?  ��� ? ���� ���� ��]��|�_U�?|�^UU������?�ݭ������ ���� ��� ? �s=?  \U�?  ��?   �?                                 �?  ��?  \U�� �s=�  ���0? ���� ���� ��]��|�_U�?|�^UU������?�ݭ������ ���� ���0? �s=�  \U�� ��?   �?                           TUU U�_ ��U ]U�U�}U���U����W������]��_}�_U�}�^UU�������ݭ��_��������W���U�}U]U�U��U U�_  TUU                    TUU U�_ ��U ]U��_�}�U���u����W������]��_}�_U�}�^UU�������ݭ��_��������W���u�}�U]U��_��U U�_  TUU                          �   �>   �j=?  �s�� ���?  ���� ���� ��]��|�U�?|�zUU������?��������� ���� ���?  �s�� �j=?  �>    �                             �   �o>  ��  �j=?  �s�� ���?  ���� ���� ��]��|���?|���_������?��������� ���� ���?  �s�� �j=?  ��   �o>    �                UU   P@  �  �> P�j=?@�s�����? ��������P��]��_}�U�}�zUU�����������_����P�������? �s���j=?@�> P �   P@   UU          UU   P�C  �o> ��P�j=?@�s�����? ��������P��]��_}���}���_�����������_����P�������? �s���j=?@��P �o>  P�C   UU  ����                      ��    ��   ���   ��� �����������|}UU��ח���:ח���:|����������� �����   ���   ���    ��    ��                                                                      �� �����������|}U��������ח���������������� �����    ��                                                                                           ��� ����� �WUU���������������������  ���                                                                                               �� ������������WUU��ח���������|����������� �����    ��                                                                                    ? � �����>�����ͫꫪ���ꫪ���ꫪ���ꫪ������ͫ�>�������? � �                                                                        < � ?���:�?��:����:��W�:��W�:��W�:��W�:����:�?��:���:< � ?                                                                         ?  �  �  �  W���  W���  W���  Wկ�  Wկ�  W���  W���  W���  �  �  ?  �                                                                         � � <\��?\����?\U���?\U���?\U���?\U���?\U���?\U���?\����?\��?� � <                                                                    ��   ���? ���Z������>������������UUUUUUU��UUUU��UUUU_UUUU����������������>����� ���?   ��                                                    ��   ��? ���_������>������������UUUUUUU_��_UU_��_UU_UUUU����������������>����� ���?   ��                                                    ��   ���? ���Z������?������������UUUUUUU_UU��U_UU��U_UUUU�����������������?����� ���?   ��                                                    ��   ���? ���Z������>������������UUUUUU�_UUUU�_UUUUU_UUUU�����������������>����� ���?   ��                                         �     �   �   �e9  �Z�� �����Z��j9�����l����5����6�����;����������; ���� ����  ��;   ��    �    �                                   �   ��   �V9  �k��  �����k��j�����9l���������5    �6�����;쫪�������;�뫪� ���� ���   ��;   ��    �                            �    �   �Z9  �� ��V���Z���l���j�����9 ����?   �5    �6   ��; ����?�����;쯪������������ ��   ��;    �    �                      �?  ���� ���U��jU�j🪪j ����9  ���9   ��9   ��    �5    �6    �;   ��   ��;  ���; ����;𿪪����������� ����    �?                         �    ��   ��   ��   ��   �������������_UUU�믪��ꫪ����������������������   ��   ��   ��   ��     �                                      �     ��   ��   ��   �� ������������oU�UUի�����믪���ﯪ����������������   ��   ��   ��   ��                                           �    ��   ��   ��   �������������oUU�_ի���ꫪ���ꯪ���꼪������������   ��   ��   ��     �                                            ��   ��   ��   ��   �������������oUUUU�����������ꯪ��꼪���������  ��   ��   ��   ��    �                                                                           �    �W   |��  ���Z� W���U����j��ë��> ��� ��                                                                                      �    �    �6    �6   ���?  W�j�  ���  ���  ����  ��?                                                                                              �    �W   ���  ���Z� W���U����j��ë��> ��� ��                                                                                                             �����?WUUUUի����ګ����ꫪ���������?                                                                                �    ��    ��    ��  0��  0��  ���  ����  �Z�  �Z9   ���  �:   ��   ��    �     0     0     0     0     �    ��   �Z   �Z9   ���  �:   ���  ����   ���   0��  0��   ��   ��    ��    �                                                          ?    ��   ��   �V  ��j�   ��  ��  ���  k9?  �j�  ���  ���    �;    �?    �                                                                                        �    �>    k9   �j�   ���  ���   �;?   ���  �   �V  ��j�   ��   �   ��    ?                              �    �<   �� <  ��<  ����  ���� �UUU �UUU9 �ZUU9 ����: ���� ���� ����  ��<  �� <  �<   �                                               ��  ��  < <  � <  ����  ���� �UUU �UUU9 �ZUU9 ����: ���� ���� ����  � <  < <  ��   ��                                            � <  � <  �<  �<  ����  ���� �UUU �UUU9 �ZUU9 ����: ���� ���� ����  �<  �<  � <  � <                                             �    ��   ��  �  ����  ���� �UUU �UUU9 �ZUU9 ����: ���� ���� ����  �  ��   ��    �                                 �    �    �:    �:    �:    � ?  ��������Z�Z�Z��j�Z����Z����Z����Z^U? �Z^U; �Z^U; �Z^U�?��_U�: WUU�:�����:��_׫:��_��?����   �    �>    �:   ���   ��� ? ����� �:�� �>�Z ���j ���� ���� ���� ��?  ���;  ��U;  ��U;  ��U;  ��U;  ��U� ����������]���]�  ����   �   �_�   �U�? pUU��pUU��pUU�ZpUU�j�U����_�����_����Z�? ��Z�; ��Z�; ��Z�; ��Z^; ��Z^; 0�Z^;  �Z^�? ����:    �:�����:��_׫:��_��?����   �    �>    �:   ���   ��� ? ����� �:�� �>�Z0���j��������������? ���; ��U; 0��U;  ����� ���U� ���U� ���U�����U��u��U��u��U�������  �7W��7            ��   �VU
  h���  �_՟��UU}
�}UU�	`_UU�'`W��U'�W��V��U��V��U��V��U��U��U�jU��U�VU��W�VU�`W�VU'`_�U�'�}UU�	��UU}
 �_՟ h���  �VU
   ��          ��   �VU
  h���  �_՟��UU}
�}UU�	`_UU�'`WUUU'�W�kU��U��U��U�UU��U�kU��U��U��U]�U��W�kU�`W�ZU'`_UU�'�}UU�	��UU}
 �_՟ h���  �VU
   ��  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@� �� @� �� ������@� � ���� ���� ��   �� ��� �� ��� �������� � 00�� ���� ��   ,�����,�����������,��� pp�� ���� ��   M�����M�����������M��� ��� ������ �   ��� m��� ��   �   �  � � �   ��09 �   � ������ ���? ��? ������ �   �� �   � �����   � ���: ��: ������ �   ��� �   ������   � ���: ��: ������ � � ��� �   �������� ���? ��? ������ � ��� �   ���� m��� m�   �   �l� � � �m�: �   ��������������   ��� ��� ����� ���� ��������������   ���� �0�� ���� ����� ���� �� ��� ����   �� � �p�� �� � ����� ��� @� �� ����   @� � ���� @� � ����                                                                                                �� �� @� �� @� �� @� ���� �� �� �� ���� ��� �� ��� �� ��� �� ���� �� 0� 0��������,��K��,��K��,������ �� p� p��믫���M�����M�����M������ �� �������묯� ���� ���� ��� � � �� ��L���� 묷� ���� m��� m��  � � �� �뜳��: 묳� �� ���� ������  � � �� �묳 � 묳� �� ����� ����� � � �� �묳 � 묳� ������ �4��� @�� � � �� �뭳��: 묳� ��m�� ���: � m � � l��� ���0�� ���� ����   �~���� G� � ���: ������ �� �����   ��� ���� � ����� ����� �� ��� �   �� ���  � ��� �� ���� �� �@� �   @��� �@�  � �� ��  @��� �                                                                                                � ����@�  � �� @�  �� ���@� ���@� @� � 0�����  � L�� ��  �� ����� ����� �� � p���,���� ���,����� ���,�����,��,�������M��p� ������0�� ���M�����M��M���m �� ����   ����:� �   �    ��l���� p: �<�� @��}���� �� ��  �� �������� � �O� � � ���� ��� ���  �8 ��������  � 듿 � ,�� ����������� p9 ����@� ��  �� � M��<����������� 0 ���@�� � 09  ��l � �  � m���  m�m l �l  m � ������� ������������ � ���� � ������0�� ������  � ������ � ������ � ����� p�� �����   � �� ��  � �� ��  � ���@� ��� ���@�   � @� @�  � @� @�                                                                                                 ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ ����  ��� � �.� � �-� ��" ����dͩ�ϩ�Ω �Ʃ��ǥǅťƅ� `����r� ���ǀ�d�ȩ����ǥǅťƅ�dͩ�� `����ɥɅťȅĩ�Ω�� `����D� ��L\� �� ���ǅũ�Υƅĩ �� ����i�ƅ� `��ȅĩ�� ����8��ȅ� `����T� ��L����ϩ�Ω�ͩL�ĩJ�� `�  ��2 ������ `�܍ � �� � �� � �O� � � �ةv� � � � � �2� � �O� � ��	@� � � ����� � `H�Z��
��ׁ� �؁��΅ʥυ˥Ņ̦Ž҃�н���ѥ�JJ�� %���� �����Ȁ����
�̥υ��L�z�h`H� �� `�����h`H�Z�/���� ���� ��z�h`݁͂̃ ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                     0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^_____`````aaaaaabbbbbccccc��������i����!� 	� \ 'q 2!"4VDEh��h�ۻ��������������������������쇾�Ez�Fu  Q                            #42#VeVf��w����˽���������������˪��ۘ�������������������������������������������������������������̻��������˻�̻�����������ffvUDC332                          "#324D3DUUUVfgffwwgxwwwx�ww�ww��wwwwwwwwvgwfgvffffgvgwwwwwwx����������������������������˻�������������wwffeUUTDD3333""""""""""""#333DDDDUUVffwwwx���������������������������������������������������������������˻�������������������wwwwwvfffffffUUUUUUUUUUUUUUTEUUTDDDDDDDDDDDDDDDDDEUUUUUUUUUUUUUUUUUUUUUUUUUeVfffffffffffffffffffgwwwwwwwwwwwwwx��������������������������������������������������������������������������������������������������������wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww�������������������������������������������������������������������������������������������������������������g�@�KV�������o���  �   `    ���(���������������@�0���P���������             �PJm�~���������������������ٶ�
p\_��I�P                       ?o�������������������o�u� b        # @(� @          8��������������������������W�B�a       ��<P�R����)"�?��Tf����������������������&�@              $ %Sl������̞��)�50F��X��������������������o�d��Q                @�n��������������������{猃z��4sWRfGA aEf����W�h���v�6Tc�8TFr$&eVTVGC�k���������������������eW2 0            E8GU>���������������z��G��X6=U4q6G�S�xF������G��5K�1b Q3B#5F�$�3xuh�W�EGu�������ܬ��������������ʗ�cU       4!��e�����x���ݚ���������}ּ��ic{e~�3f�uId�X�x�y{v~ۅz�gxw�y����W���ggGde#Ev%dGSTFggtifkhf����������������ۻ���8CfT3$1tTSTGBx%TJe�eewsw�V�xdytxY��������������������tFC3   10SWf����̻�쬺�ʌ����ewFg4r$"%2V2eGdh��z����̽�������ܺ����wVvT%TDER2D32UcU6cxww��y��������w�j��g�w��v������̬����������˪�v�44#       !DdXx�������������껩�v�WwfvdvFvVwgwy��y�j���xvvFwDfWuwV�v�x������̫�˻����G�WeT5DVDFefV�v�����۫�ܼ�ܺ�����xwvfVfwgewffwhvw�f�wx������g�wvh�x���������v�wehdVVeF�Wxv�y��˹���������ۛ��efD3       35Txx��������������ʺ���eeEcED5ETFvfvy����������xx�fuWUeUFfWfWww�y������ܽ��̺������gugeUFeFTTFffxw�x�����˼˻�����wuUUDD3B"""4CUUvx��������������̺���xeUUDB4"31#3DDTVUWvVwvgx��������������˻������x�wudUTDTDDUEfwhh�x���������������xxwgwgfgWgww���������������������������x�x��wfwfUVTTETEDUVffy���������̻�̻�����wvuVdUDDUUCUVVgx��������������y�wvwufefVeffgww�������������������wwfvgfffVfvfVfvww�wx���������������wvwwgwvwwwwxw�w�����������whvfEVUVeeVfwww���������˼������ufUTCDC3DDDDVff����������̻��������wffTeVEEUUUffw�����������������wwvffVeUeUUVUWgxx�����������������wvfeEDUDDDTUEUfvwx������̼�̼�����wfeTD332"#333DEffx�������������̻�����fUTD4333C4DEUVfgw�����������������wwwwvfffffgwww����������������wwwfffUUUUUUVVfffwx�����������������������wwfffffffffffffgwwwx���������������������Ex���wwgw�ʇCX�wdi�g���Fwwg�vg���fx�y��eeEVX�˩��d3Vwx��fx�����gffUVy����vgw���wxwh������wwwveUffg�������vwww�weUy������UTDDy������w�wvfxweg���xwwfwy��xw�gw������Vw��w���g���eeVf�����ffT5z�vgw�V������AX�̨eTf�x̧fh��vUC$W���̩uC#Fx�������weVDT5�gx������Wy�veVfxvEX����ܻ��VD4$V���ܪzx���xH6d�f8X�șYf��z���7���Y��Y��h���G��Y��YY��e�ze��wfWd�Wx�xfx����ɧj���e�RtZ�hW�����iiU��xXE��؊xz���I���eWX����Xd�x�W��Ǚf��iHU��hS�Y���gy���J���Jv��Xf���d�H�w��˦c:�VuY���ec)f��|�yi&s7U��{�����5Qf���7t����i���5v%wtI�Ɋٸ2aH�׼��X��8�k���bVCU�y�I����7�z��h�|ٽ��x�XuudaX�i�ى�x�hsz��������R�F�fdx�jțǌ�z�7�Fw5�e|�i�w�E�x������v��hfVv5j�i����UwuF�������fz�w��evuU���wvWz�i��v��vE��y�yWw�������WUg���������Ww�DF��xh������fVvE6������fXx��v�wx��hvv����xih�w����gVG�������V6ef���wXVUvw���xfDe����z�yw�uv�����vwwfXg�����xhgvv��zxuDu�������dF7g���fXy�����iy��dE6W�����U3Sw��xx������vtfWWx���fWw����yw���xhfeuiy���tEGWx���j��w�i��udEFy�ʻ��ecfXw�����w�vVEV���hx����W���gfevx����g����hx����z����yv�whi���xYw�fgy���wvvW����h��vWy���yw�eWg�����wfew���vvy����ggfw���wvg�w��xxyx�������hffvxxwwwg����������wvvgxwveegx�������gx����xveeVg��ghw������x��vvwh��xgf���x����w������wgv�fgx������xgfwxx���wx���gffwx������ ̋�̈�����̊�����w�x��xx��x�xxxx�xx��xx�x�����޷   &��˻����0  7�쇗E�j��hz�   ��ނ6v��}���   N��@  -�����@    f�`��#����   O���   ~������     ������   {�sXh�   >�������     I�����    |�� l���  ����p    �P (�����   5 
�����       ����� ����0      W�������    ����    ���  ������   ����  ���dM����          ������0     ����  -���������     '�����   �W�  ޾������      (�� o������     L����  L���   ����b    "7r3m���   ������    ^����    ����  ,�����0     ������   ��������     �����     ����`    5e��������     j��P&�   �������       ,��� m����     �����c     ����������    TU    =����    n���p    ����  ����P    +��   ,������t       (����3���  �����  %P������     V����  ����   �ܾ���  Y����    |����������      ���   &��������  ����0   N�����     D3 ��������     9�����0       ���������      3D ,��������  �����   ������   EeCEfD{���P �����u    ����vx����      J� �����   �����P    j̦����e   8���܃  H������  ������vA    J��  ��������     DV�1L���1   =�����   h�rY���  F��̥  	�������@      h�����b   ��������Q     �������      <���  (�������      7�u16�����    �����q   �����1    Vx���16�ʪ�������      �����   )������@    ^�����P     ��˙���a   )��ډ������     i�������    W������q     G����  ��B��������b      (����uVh�u   i��������    ����������        �����@   J�������        �������v0   F��@��������     C$������̸04Ed4y��R   }���F��������b       H���̺���ܕ2   �������   ���ܹQ   ����   �������     $T!6����   H��������0       m����   �������c     �����0   ����t   ]��؊�vwwxc   �����q    )�����T1   '����ۘS     ���������d    UVx�������uUW�̺a  $��������S     }������@    �����A    k�� ;��������A     5g������0    j�������Q     {����  I��dDW��0 ���@   �����4z���̺�0    W����Q ����0   &�����  =���ۗS    4T����������1     F���̺��Vfg������ݹuB !#X����fgx����d    z������R #D1 ���������t    h����  ������S      H��������S     ;�����wA    �����0    ���r ������˅    EUUUdK��������t     �����P F����u  ������˅      X�ʙ�����0    ������@    \�����0   �������ۖ0      5����uUw����̺�0   '������r  ����ʫ̸c     h����ܩv  ��r ����Q  G�̩���ۄ   ������ܨR   y���˨S! Z����۪��@  ����uDUB   ���ʫ�˺�feT2   X���ܻ�d!F��������ܖ1   y�����Q 5xuW������ܹc   j����̻�  z��˘R  6���d"6���쩘��R   X���ܻ˧0  z�ݹvC"$h��g�����    G������t  #l�����e2  Y���˩�0 $h�������0   j���TG����  5feg����̺�1   $y��˘��d"5��ܺ�u1 k���˻�u2 "4Eh����vU1  [���fy���R   #Vy�����   G����څ1 4W�����u14h���ۅ 4Y���˪��1  ���ʆeT334Vy��u1 '�����B  z���˺��c  #Ug����ۘvDEUC 7���UVx���eDUeS 8�����332#W�����dC34Fx�̻�vTDVx����vC#W���gy��b �����eUD2""G�������x�wfg���S ����uDDDDDW����wfffw�����vT3Fy�̺�vffS|����veT34Ufgx�����wwvfg����vS 8����eUVeC3Ey���fgx�������vffffg����vefffg����vTDEy��ܹ�eEUUT2%����˘vUC34Vx�wwx���wvffg����wwvfeUUfx���fgx������vffveDDVw���ܹuUfgwwvfffx���ww�wwfx���vgx�wfUg���˩�vUUUVgw�w��wwwwvfw��˩vVffw����wwffeDV����vfx��wfffw���wffx��ww����wffgx��veVw�������vVffffgx���������wx���ffffww���vwx��wwx����wwgffgx�����vfg������wwffffgx������wfefffgx�������wffffx����wvffx������wfUC4F���������wwwfeUDEg�������wwwwwwveC4i��ʘ�x�vfffwx�veVg�������wvfffgx�����wwwwwwww������wvffgfwx�������wvfeTUg����������vfffeUVx��������wwwvfeUg������������wvfUVffx��������wwwfUUfx����������wwvfUUUh�������wvffffw�������������vfUfg��������wwwwwwfwx��������ww��wvffww��wx����������wwwfveUUx�˩�x����wfwwwvfUfx��������wwxwwwwwwwww���www�����wvfeUVw��������wwwfwx�w�x���wwx�������veUgx���w�������wfUUUg�����wx����wwwwfffx�������www��������fUUg��������wwx��www�wwwwwx�������wvffwxwwww���������wwwwwxwwx���wfffw���������wwwwwwwwwx�wfffg���������wwwwwwvgvwwx���wwwwx���w���������wwwwwww���wwwwwvgx�������wwwwwwwx��wwwgww��������www�wwwwwwwwwww�wffw���������vfwwwwwww������wwvffg����������wwwwwww�wwww���wwwwwffg����������wwwwwwwfwwwx�����wwwwwfw����w�����������wwwwwwwwwwwx�wwwx�wffw���������w����wwwwwwwwx���wwffwx����������www�wwwwwx�www��wwwwvwwww���������wwwwww��wwwx�wwwx��wx���wwwwww�����w���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������                                                                  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������                																















 @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @��    				



    !!!!""""####$$$$%%%%&&&&''''(((())))****++++,,,,----....////0000111122223333444455556666777788889999::::;;;;<<<<====>>>>???? 0333<???<???<???0333<???<???<???0333<???<???<???������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@dxآ�� 3� �� ���X� ��  ��  �� ��dxآ�� �� � ����X � � ��L��� � � ����� � � @�Ј`��������0���P���p� ��� ���@� @�  � ��  � �� 0R��R�JR�����΂7 ^ 2C ; U7 - 39 - 9 - 3E > R9 ( 8; - ; - 3? ( hB ) 7G + 5; ( ; ) ; , ���> - ; 4 ,7 ? Q> 7 )@ * = 9 '9 < T@ 1 /? ) B ; %? B ;  ? " B & 
G 6 �� �Ɇ �� �Ɇ �� �Ɇ `� �Ɇ �� �Ɇ �� �Ɇ `� �Ɇ �� �Ɇ �� �Ɇ `� �Ɇ `� �Ɇ 0� �Ɇ 0� �Ɇ 0��	$   �$   �$   ��� �                        �                        �                        �� 
��         �
         �         �� 
��
 2   2   2   2   2   2  ��  �0   �0   �	  ��  �0   �0   �	  ��ʽ�    �ʧ�    �ˠ�    ����K�  D�A�    }�z�    ����������������������������������������������������������������?<<<300030003000                           ?<<<300030003000                           ?<<<300030003000                           0123456789ABCDEF �  �  �  �     ����     U��0�����?� @��v
�F�F��o/�R"�ʢ|X7�����zdP=+����Ǽ������}voic]XSNJFB>:741.+)&$"                                                  $ ( ,   $(,  $(,      
             " $ & ( * , . ������������������������Y��������?�?�?<��??<? ?0�������??<?<?0?<?<?<?<?<? ? ?0?<�?<??? �<?<?<?<?<?<?<�?<?<?0?<?<?<? ?<? ? ? ?<� <�? �??<?<?<?<?<? �?<?<?0?<?<�? ?<��??�?� <�? ?3?<?<?<?0���?<?<?0��??<? ?<? ? ?<?<� <�? ?0?<?<�??? <�?<???3?<?<?<?0?<? ? ?<?<�?<???<?0?<?<? ?????<�?<��??<?<����?? �?<��?<�??0?<�? �<??�����<?<                                                ?<�?����?<�?�?�?��        ��UU  UU  UU  ?<???<�?<?<?<? ?  <?<?<    ���<?�UU  UU  UU  ?<�?<� < <?<�� ??<?<    ��� ?�UU  UU  UU  ��?<���?< <?< �?<    �??��UU  UU  UU  �� ?<�?  <�? <?<�?<�?        ��UU  UU  UU  �?<?<�? ?< <?<?<�?< <� �        UU  UU  UU  ��?���?� <������ �    ��UU  UU  UU                            �         UU  UU  UU    0 0     0  0 00  0      00     0   00   0 0     SHIPS SCR WAVE  MATTA BLATTA HALL OF FAME  # Q u � � U  ��xd(

7Ҹ�ӹ�3�n��ӸҀ�   �   �   �   �   �   �   �   ����������������������������������������������������� � � �d��������������  ������������������������������������  ����d � � � ���������� � � ����   �� ������������������ � � � ����������    ��� � ���� � � � �����d� � � � � � � � � � � �     � � � � � � � �  � � � �d��������� � ����������������� � d���� � � � �� � � � ����        ������������ � � � � � � � �d� � � � �  � � � � � � � �� � � � � � � � d� � � � � � � � � �            � � � �� � � � � � � �                  � �d � � � � � � � � �MONTANA!    MR. SOSA    FRANK LOPEZ GINA        CHICO       ERNIE       MAMA        ELVIRA      OMAR SWAREZ MANOLO                            P      P   %    P          ABCDEFGHIJKLMNOPQRSTUVWXYZ. ?!Great Score! H�Zح' J��$  �Հ	J��%  ��z�h@���# `�`H�Zإ�K� � JրA��  I��'��!) ���')���')��� �P� H�H�H ���h�h�h� �Qz�h@�����`�EH� �ץ �עdd &&&8������������ ���h �צ� `�EH� �ץ �עd d! &! &��e � �e!�!���!� h |׆!� `�SI��S�UI��U8�R�T�S�U`� � ����`� ��`
� ��e � �i ��� �� �� �` �l  � Z� �� � ���� ��0��z����`Z� �� �L�N����L�N�M�O�0��z����`	 I�i`H� |�h`H�I���I�����h`�e � �`�`�e��`�`�eL�L�`�M`e(�(�`�)`eN�N�`�O`H� I�� �I��� ��h`H�I���I�����h`ڢ �JJJM
j.
....����` �׆��
�L ؊H |�8�����8��������h |�`� I�� �I��� ��`�� H�H�&H�1H�� d ۩  ��h�1h�&h�h� ``���H�K)�Kh




K�K�& `H�Z� ��  	 � �� � ȱ � ȱ � ��� z�h`�'��Q�Q������������`dQ�Q��`x �ة�X`�X�Yd1�
&1
&1
&1
&1�(�1�)�(
&1e(�(�1e)	@�)�JJe(�(��)ڊ)�1��>ͅ5�0�:�%5�4�1�`�{�G�a��a`�[�<�A��A`�:��0��`�.��$`�,��%`�'��&`�"��'`�?��(`�!��)`�`��H�Π� ׎�h�	i


����I�,�� ��� ��Z ��z��m��I��JL��H�m�h�`lH �ة ��h E٢͠� טi �L�i��M�1
i����	��&�	� ��L� � (�(�� ������(�(�(i0�(��)�Li0�L��M�&��`H �ة  ��h� ���L�� E٢Π. טi��L�i΅M�1
i���&H��	��&�	� ��L� � (�(�� ������(�(�(i0�(��)�Li0�L��M�&��h�&`�� �L�(�(��)ȱL�(�(i/�(��)����`�')H���H�*���G�Hh`� ����Z �آ�
� �(���(i0�(��)���z���&�&HZ�.*.*.*.*)��
��� Y�hzi�h�&�&��`�')����')���`�Q�
I|�I5�	�I�` �إ4�(`�(H�)H�e1iJJ�
�
ڦ1�B�I��he1)��F�I��	��� �(%�(� �
�ȑ(���(%	�(�(i0�(��)���h�)h�(`�Z�(H�)H�	�e1iJJ��ʆ
�0�N��O� �(�Nȥ)�Nȥ
�Nȥ	�N� �צ	�
�(�N���(i0�(��)� �����h�)h�(z�`�0�(�1�)�2�
��3�	�4�L��M�	�
�L�(���(i0�(��)� �����`�(H�)H��1�>�I��	��(%	4�(�(i0�(��)���h�)h�(`��e1JJ�	�1�B�I�2(�(�0�:�=B�(�(��0�:��	��(��	���e1)��F�I�1(�(ڦ0�:��=F�(�(`�+�,�X�)�Y�*� �ܭ*m,8���) �خ+� �ܮ)�* �ج, �ܬ*�)m+8�� �ج,L�ܩ `�X�Y�� �* ���Y0�X SޥYe-A��8�Y�-�8�Ye-�`��-8�� ��-�,JJJ�dd �֘e*�*�e+�+�X�  Sޥ1
i��i��Ƞ �� ���.0 �إ,iJJ�	�(8�	�
�-�&�	� �(I���*���� ��� I��(ȱ(I�I���֑(�(i(�(��)�*e	�*��+�&д`�X�Yd1�
&1
&1
&1�(�1�)�(
&1
&1e(�(�1e)i�)�JJe(�(��)ڊ)�1��>ͅ5�0�:�%5�4�1�`��`�چ[�
�\�J�-�I�\�]^�A�\ie�� � ���0�[�J�-�&�\�ef��[�0�\�],�]��^)�ߠ� #׀Ѐm)����
I

��@�  !��TH�[�	��h}���I

�ڹS͝ ��͝ �\i]� ��ڦ[�)� zߊ�\�e�f�	@�� �[�	@� ��0L��`H� � �֡ �  ��he � ��)�Ff Ff Ff �[�)���� `������n����!�K���;�`�[
i]�� �[�L�֦[�J�I�-��� � ��� ���� ���( `�)������ ��� �( �`�\i]�ڦ[�)� zߊ�\�e�f`�\�]�]��^�[�`�\i]�� H �֡ � �֡  �֪��h`hL�ح8�


e\��\��˙] ��˙^ �[�`���� ��� �( �* ��L�


�� ��˙] ��������etf������������`Matta Blatta Press start to play Get Ready! �F� o� ����� �� ���0� �  �آ���  ��0�� �آ���  ��0�� �آ���  ݩ�I���J�(�� �٩�I���J� �"� �٩
���I���J��P�  �٢ � �إ'�)��0���P �آ�� �ۢ � �إ'�)�����л�'�)��L� ���P �آ��
 �۩�I��J�(�P�  �٩< �ة `�X�Y�/� ڦX�Y �آ���hH�/���0�M�L �ڥYi�Y�����`Pause � ��')��`� ��� ��+ c�  �إ')����')���� L_܆J�I� �I�����



�2��8�2Jm.H8���-i8�Z �إ2i�ڠ  �� �۩�0��   �hi���L�� �� _� �� �񢂠 �:�9 /� 1� ,� �� �� �� ��� ��
 � ���r�ح�
���ѭ�
)�ʭjk��
�2��
�����
�s�  ����
�� �� � �� Q� p� p� J� �� O� #� � �� �� � �� ��L>�?����	 �׭
)�ް	���p	��ѝ�	�0
 �׭
�0	��` d� �䩐�l��m�ȍj�k�t�i�u�
�p
�F�~
��
��
��
��
��
��
��
��
��
��
��
��
 	� � � ��&�|
��}
�p��
���
��=��;��<���
`��
���S� �jk�`�k��j�Z�ک ����j��k�j�jk�	��jJ���i

�
��Wɍ�
�Xɍ�
`�lm�&�l��m�l�lm����n �׭
)?i �o�nɌ�X�n�n�L��nJJ��o 孀
0;��
8�nI�i��)��
8�oI�i����j��k ����L��`�čl��m���n`�>� ���(�>���?��@�A�B��C�n�oLuݩ>� �����>���?��@�A�B��C�p�qLuݜr�q���p`�r���r���p �׭
)i@�q�pɌ�`�p�p�Ld�pJJ��q 9孀
`��
8�pI�i��x��
8�qI�i��f ��i���t����
�	���
�t ���t��i�i

��jk���jJ��e��
��Wɍ�
�Xɍ�
 d���L��` +� Q��
���
`�')0�9��
04� ��
������&Z�i��Ս�
��ɠ� ��z��
i��
��
iD��
`���
���
��
��
��
 ����`8`���
J�/J�,��
8�8��
I�i�
���
8�8��
I�i��8`���`���
J�)J�&��
8��
I�i����
8��
I�i��8`���`� ��
��
��
��
���
�܅I�хJ� �� �٩օI�хJ�d� �L�٢ ��
 ���
 ���
 ���
 �瞅
��  �آ8� �۩��I�
�J�� �L��HJJJJ	0��
�h)	0��
�`��

����m�
��
� �m�
��
��
i ��
��
i )��
�LP����
i%��
��
i ��
��
i )��
�LP� P碔�  �آ� �ۭ�
	0��� LYک ��
��
��
��
���
��J	��
` l��
��	��
��
�8�ҝ�
�� ��
���`��i��
�y��ɠ�� ��
��`��
� ���
����`���
J����`��
8�8ɀ���
��
��
i��
`��
i���
i�	��
J�4J�1���
�'8�8�I�i�
���
8�88�	I�i�
�8`���`��
01��
�,�|
��}
�|
�|
}
��
���
�d�~
���
i��
�`��
��	�s��s`���
J������&�|
��}
��
02�~
�,�
��
�	��
� ��

���ԍ9��ԍ: �� ��
��
`��
� �L&ɩȍj �� ��
��
��
��
��
�t���t�t�i�t`� � � � � � � � � � � � � � � � � � � � � � ���`�'����D����D����D��E�@�@E�h�pE����E����E��� F��0F�0�`F�X��F����F����F��� G���PG� ��G�H��G�p��G���H���@H���pH���H�8��H�`� I���0I���`I����I� ��I�(��I�P� J�x�PJ����J����J����J��K�@�@K�h�pK����K����K��� L��0L�0�`L�X��L����L����L��� M���PM� ��M�H��M�p��M���N���@N���pN���N�8��N�`� O���0O���`O����O� ��O�(��O�P� P�x�PP����P����P����P��Q�@�@Q�h�pQ����Q����Q��� R��0R�0�`R�X��R����R����R��� S���PS� ��S�H��S�p��S���T���@T���pT���T�8��T�`� U���0U���`U����U� ��U�(��U�P� V�x�PV����V����V����V��W�@�@W�h�pW����W����W��� X��0X�0�`X�X��X����X����X��� Y���PY� ��Y�H��Y�p��Y���Z���@Z���pZ���Z�8��Z�0L�`� �N��O� ڽp	�	�0	ɠ��JJ��)��	�:ͦ=>͑N�P �����@��`�?��	��0
��	��	}0	�0	��`���i�� �i�����A�� ��[�����A�	� �
�[���� �����
��� ������� 8� � �� ��  �ץi0����i0����i0���	�
i0�
���П`�=�`��= P��;�z��;�9�i�� �:�i��<�<� �� �<H ��h �ש���A��(��[��� ���� 8� � �� ��i ����i0����i0������`�N�A�'~�A�����N�A�'~�A�����NB�'~�A�����N8B�'~B�����NhB�'~@B�����N�B�'~pB�����N�B�'~�B�����N�B�'~�B�����N(C�'~ C�����NXC�'~0C�����N�C�'~`C�����N�C�'~�C�����N�C�'~�C�����ND�'~�C�����NHD�'~ D�����NxD�'~PD�����N([�'~ [�����NX[�'~0[�����N�[�'~`[�����N�[�'~�[�����N�[�'~�[�����N\�'~�[�����NH\�'~ \�����Nx\�'~P\�����N�\�'~�\�����N�\�'~�\�����N]�'~�\�����N8]�'~]�����Nh]�'~@]�����N�]�'~p]�����N�]�'~�]�����N�]�'~�]�����`�ک}� �Ʌ��
8�:��{���
�8����� u����آک}� �Ʌ��
8�:��{���
�8����� u����`�~
�`���I�хJ�0�P�  �٭�
JJJJ	0��
��
)	0��
��
���I�
�J�X�P� L��H���ȕ�H���Ȟ�H� � �@�`�  � � ��
��h�������	��`�Z����
J�;�>� ����
�>��
�?��@�A�B��C��
8�:���
8������h u�z�и�>� ����
�>��
�?��@�A�B��C��
��
Luݭ�
)�C��
0>�')��� ��m�
��ɀ���
�*� ��m�
ɨ��@���
��
��
��
8�@��
`ڮi��

�` @Xp�����
`��

����!�)������
����
����
� �1�	 �׭
)?	�����
�)i���
�ж`��
�>���
J�3�=	���)���	��	����)�!��
	)���
��`���
J�L�J�<�!�r�)�!�����
)���
�0��
���
 W�N���
i���
���
�;J�8�!�3�)�!��
i���
���
�������
8����
��
���
�0L��`ک�ɠ� �����
	��
� ��
����
� ���!�)`��

��%҅ �&҅���
J�u)�q�1� �d�� �1L[� ���
)��}�
��
��
q ��
Ƚ�
q ��
��
)���
0��
8��
��
��
���
��
Ș�1��
)�����1��`�� ��
J�n)�j��
i��`��
�
��
)���
�Q ���u�u���u��
i


��)����
	��
�)J��
)?i�e��
�)
i0��
�1����`��
)�X��
�`� �1�	����
 �׭
)i



��
 �׭
	���
	��
��

�����
����
�����!�)`� ��ԝ ������ �i՝���,��` � ��� �L��M�0�N��O�
�� �N��L�N���Li�L��M�Ni�N��O��٩�� ���=����
�&� �  ����  ���� � ���� � ���� �� i� ���i����&���0�I��J�
�&��<�&H�Z�IH�JH�  ��h�Jh�I�Ii�I�Ji �Jhi
��h�&�&�Щ=�I��J�
�&�f�<�&H�Z�IH�JH�  ��h�Jh�I�Ii�I�Ji �Jhi
��h�&�&��`HJJJJ	0��h)	0�`�'�`hh�'��`��� ���
�8� ��
���� 8�� ������F`�
���D�
8�D�E��F`�
�


8�i�X�

�

ei`�Y�X�Y �آ�L � � &��  �� ��'����K��d�g�h ���g�h��0 E��
 �إ'��Hd0�g�h E���)��LN��)0�&�)���mg0�
��g�*�mh0���h��� ��h
�

emg���Յ�?���ʩ �K���KH�
�

ei��Mh Y� ���')0����?�����L���������')����F�E�&�w�� �ʈ���&��E�&�'�����ʈ���&��D

�
e�� �K� ������D

�� ��
�������`��0�d0�
�

ei��Y �آ
L�ܩ � �A��	� �� +ש@� �B������ +ש`� �C�����U +ש�I�хJ� ��  �٩�I�хJ� � � L�� �����I�ՅJ� �@�  �٩���Յ�d�Y��
�X�
ZڦX�Y���� YڥXi�X����z�Yi�Y��ө�0��V �آx �ܢ�K �آx �ܢz�� �آ� �ۢz�� �ةG�L�ɅML�ڜ���� ��� �0�0���`���  � � � ���#  �������K�& ` �� � � � `� � � � `H�Z� H�H� � �@�� �  )�h�h� z�h`� � ����  )ע t ���`�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������