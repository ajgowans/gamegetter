                                                                  UU  UU  UU  UU  UU  �W  �W  �W   W   T   T   T   T   T   T   TUUU�U=U�U�U�U�U�U���UU��UU��UU��UU��UU��U���U���U���U���U���U�PUUP�UUP�UUS�UU_�UUU�U�U�UUU�UUU�UUU�UUZ�U�Z�UUZ�UUZ�UU[�UU_�UUU%  U�  U� U�
 U�* ���@U���U���U��U�������U���U���U��U���U��� UUU@WUU�WUU�WUU�WUU�W���WUU�WUU�WUU�WUU�W���WUU�WUU�WUU�WUU�WUUT@Wp�W|�WU�WU}�WUu�WUU�WUU�WUU�WUU�WuU�W�U�W�W�W�_�W��W��UWUUWUUUWUUUWUUUWUUUW�VUW�^UW�_UW�_UW�_UW�WUWUUUWUUUWUUUWUUUWU�                U   U   U   U   U   U                      �   �                                                        ������������� ��� ��� � � � �                                  ����������������������������                                ����j�㪪�㪪�⪪�⪪jb��������                                ��������������ꩪ�������������                                ���������������������*���
 ��                                ꪪ*���
������ ��* ��
 �� ��                                    @�  ��  ��  �  �   �   �   ��  ��  ��  �   �  ��  ��  @�     �� ���A����?������  � �� �������������� �� �� ��       �? �� �������?���?���??��??<�?? �?? �?? �?? �?? �?? �    ����������  �  �  ��� ��� ��� �  �  �  ���������     ��  �� ��? ��?�? ��? ��? ��? ��? ��? ��? � ��? ��? �� ��     �������������������������?���������� �?� �� �� � �    ��?���?���?�?  �?  �?  ����������?  �?  �?  ���?���?���?�    �  �?  �   �   �   �   �  �  �?  �  �  �?  �?   �   �                                                                                                                 	
                             !"    #$%&'(    )*+,-.    /01234                                               56789              :;<=>?@A            BCDEFGHIJK          LMNOPQRSTU         VWXYZ[\]^_`         ab cdefg                                                                    � � � �          
  � �                    ( ( �$*    % )      �                          ���jC)N`��V�R�*�B�B   �>���٩U�e��V��B	 � �R�ۗ�F ��	`)j(A
A�
               ��  . ~ � � ��
,-N=HPJ�����(z~^�^�Y0e� ��*�?K�I,l o �试����T��@@         .      ������ R             �                �           ���_y       �  7 0 ��(
*
�
�� �  
� ��b�����(�\�^@�A���V � �$J  @]@�@�U*��
���� � P�@=
=H.�
�
�#��(�? � K H , ` � � 8 6�U��V�O��@?P�WVP UP�T�U�zU����z�^����*5 ;          �   � � p { /  _w~>yT�� �¯�� ��)��|��%X~hzkA���R���?���)YRP�*� P!R                             � (����V������   UP������o����_�Vo����    U�U� @��        (�
��         ��B�� 	�
    	             |���l�l`�
� � � � 0   (    
X�� X   �            (      � ; � � � � < ��������������  ��5J:����ꪾ        ��6o钿       � ���Z�         � ��j� � ��ꯖj�������������[�o�l����+��k����
�Bk���j�
  U�����ꪥAU �@����VW__ ^��Z�UUUU@U U U� jW5y9y:��l���� � � k������k�k�������֮�k��F��k�[�F��k�Z��V�V������U�P���~�W~W _    @ T@UT� UP�T���-�Mj:���� : : �𮯫k��F  � �V������          � k�������          ��� � � � �������FU UUUUVU���__  PUUU�����@ TPUU�U����꪿��=�5������o��Z�뫿���������UUk�[�W�竾��ꩪ�k���k���寿�>�� : � ��:�:�:       ���Z�\A � �����Q�t�>�W���>�>    ����          ����? � ����kAV����Z�A�A�>�> �����> � � [�B������VjA�A�>UU�����>�>    �>h����        �)�          �T������?      �:            � � �          ��>�                         �B �            �?                                                                                  	
      !"#$%&'    ()*+,-./0123456  789  :0  ;<=     >?@ABC@A        DEFGHIFG                                                                                                                                                            ���������������������������������������������������U��E���W����������������������_gW�ַ��U�U������������������������+�J����+�����������������u�V�g�_ݿ���������������������������������������U�k�^�{v�U�֪�TOt�WUMTu�U� ���5�U�U]UUUU�   �V]��Z�W���T�����YU     �������+�
���
��@�P�P�T�T�P�����������/�/�/U_�WUU�U��   W�T�U~�����{�~�z�W՗�YUUY�   �SW^Ԕ���� �������������������������������������,���������     /  
`� �     �������n�} ~ �   "� ��kp/@ @�� ���
�+������������@� U TP
@+@�@�P�������~�������
�*@: �  � )���d�@��� ���@  �;�. > ; �  �*� ������������������_jW�]��������U�]�Qꕪ��������������������˫��� � *�� � ���������������j j���
� �@�������������@�������������������������+P+T+�
�
�B�������������������������_��U������P*��`��������ù��N�*@�@������� ���� �+ jYZ_
 : @2 |������������������������������
�. � ���������������������������o��������������W������������A�U��������������������������������������������������������?��������������?�������������? ?�?�?��������������������������?������?����� ��?����� ����� ������������?��������������?����������������������������������? �      ?���?���?���?�  ?�  ?�  ?��??��??��?�  �   �   ��� ��� ���    �� ��� ����������������� ��? ��? �� �� ����                �P �� ��� @��.����j�y��                             �  OZ �  �� P��j� �                                                            @  ��  ��  �u  �y  ��  �  ��  �n                T   �  �  G+  �  �  �  t  m�� �� J�  �j                                            ��       �  ��~  '� �
�                                             @  �  @* �
 ��                                                  �� mi  �                                   �j  Y�   ����@F `@� X�� ع�     	                                      i  '
  g  	      �*          �P �� ��� @�  (�  U� @�9   �   �   �   �   @            �  OZ �  �� P��j� ��  ��� jW j)  j  �  �          @�   �   m   �  @  �  �  p@   �   �   �   �   �   �   @    �   
   �  Z  �=  y=  X<  i>  �>  �>  i?  �  �               `VZ�����9 `�M �� @�� � 8@f   �                            �  [� �� �� �  ܪ ߤ
 u@*  �   @                        �V� U��  �.  �
  �
� V��@i��� �  l  �                                                     
   (   �?  �  (  8   �   �   �    (�� ��� ��  � �� @�* �K^ ��� ��� �	� হ �[> @�  �         ��  ��  @�   �   ��  �  
�  ��  ��  �  ��  ��  ��   �   �   �        �P �� ��� @�  ��  �  �X ��� p�� |�� �)p �  �              �  OZ �  �� P��j� �                                         P  U ����� ��Y ��b @Ub ��i��� ��  �  �                �   +   �R �� ���
Z�j�Y ��Z ��R ��X �� �j  V         
   8   �  �
 (�o� ��J�Z n*V �)e 8�Y (� �% �� �Z �        �  �  �    (  
�  n� n��k���I�J��^���a �j  P  0     0     .�     .�  n� �{��b��b��{���v@*� �V  P       V  �j �� ��X ��R ��Z�j�Y��
Z � �� �R +  �           �  �j �� �% (� 8�Y �)e n*V�J�Z� �(�o�
  �   8   
      P      �j ��a�^��J���I�k� n� n� 
�  (   � �  �      P  �Z @*���v
P��
P��
@��@�� ��  .�     .�     0     0       �     @  @
 �@
�*����	]@ͤ���@
�* �  @
  @     �              �   
 �@	�%T��*9�A3Tj�* � i �@�                                   P   $  @ �*��Z���PU��  �*                                       @ �@� � )Tj�*9�A3T��*@	�% �   
  �                                  �*PU���͐�Z�@�*  @   $   P                                           �   �   �   �   �   �  @�  �                     �   * ��� �G��������_/[ �F: �
 9]. {}�                              �?  �?                                                     T  �?   �                                                     T   �  �   /                                                 P   P  �  �      /                                         @  @  �  �  �  �  �                                         �  �  �  �   �                                                P   T     �  �  �                                                    P   W  �  �                       �                                                            ����Fk Z � { ��+ �%* �O �� ��; ��<   �                                          �  `  P	  �                                                  �  p  �9  X%  P  �                                      �  �:  [�  W�  W�  U�  X9  �                                  �   �  \  �+  �  �  �                                       �
  X=  �  �  �   �   $  @                  h)      � ����������F��ê�����*�����
�������� �  h)  h)  � ����������F��ê�����*�����
�������� �  h)  h)  � ������������F����3����*�����
�������� �  h)  h)  � ����������F��Ϫ���?�*������
������� �  h)                                  �  �                                                     �   �  �                                                     �   �  �                                                �   �   �  �  �                                             �  �  �  �  �  @  @                                             �  �  �  �                                                  /  �  �  T                                                     �/  �  �                                                                        �   �  �  �C   �               �   (   
  ��  �  �n���N|��n���V��E	�E��Z|��n                � kU+�
  &  P�@kUP �                                  0  ;�  *�  &�  &�  T                                               �   �   p  Z)  p  �   �                                       �   �  [  [  �  �                                              8  �  p  �  8                                        �   `  |  �	  �/   �                                   �  ��  �7  `~ |��� w�  �}  �  � �          
 ��8�#���*�	�f�hB�3�4F>�J���b
�R��ME>��`���I���*(
  H����N  �n  �  ��   
   (   �                                    ���0����?�������      �  ��������?0�����                    �  �  �            �  �  �              ��� �� �?  �  �  � �? �� ��? �  �  �  ��? 0�� ���    ��� �� �?  �  �  � �? ��  �?  �  �  � �? �����        0  �  ��������? ��  �?  �  �  �              ���    0�� ��? �  �  �  ��?  ��  �?  �  �  � �? �����    ���0�� ��? �  �  �  ��?  �� ��?��������?0�����    ��� �� �?  �  �  �            �  �  �              ���0����?��������? �� ��?��������?0�����    ���    0����?��������? ��  �?  �  �  � �? �����                                                                     ��D(\� ͰcfeY�}� �Z��Yp9 ���!�� (]�Ͱc�feY}� �Y��Yp9 ��� ��0\� B�c�eY"إ 3X�H@p9�� ��\��@�c�eY� 0X�@@s9 ��  $    R  L� @1`  !I @�$  P    ��     �  �@  `Y  !  � @@	  ��           �   �   `          H   F   �  ��  ��  `�  `�  ��  ��i   �   �   �   �   �   �  ��  `��?X�_�k�@� ?��Է���P���� (   � �Q
 `�* �. F� Q�
 �� �� ��  �  �/  �+  �  �
  �                                     �   �   �   �   \      |   �   \  ~�  P �  �T�U�CuU��U�^���~��mp�j{r�j�}�j�}�k{n�m�W���Aݶ]@����@���U����Wj�[~U����������������\��\�����u��_��� ��� �  �   �   /   +      
                �   �  w  3  3                                                                    ��   �   �                 ��� pt�����빪���@ǥ��ǔ���P��@]�����z�Gۯ��n�Х�0n��psk�pn�W���A��9?�z���ސm�^W��F�.��Ӯ���n��[n[��_���u�Z�Z�k@���Uz����E����Ѫ���V[�ZV��UV�VV�XVx `W� ��w       �  �             	   /   �   �
  ��  �� ��5 �k� �[U�VU ����uհy�e,u�\�eYkYe�G]�SWmYW[�G��QWk�U[lՖ�ey԰u��[�e �Zey�eu�Y�eYeYe�G]�YVmYGY�GV�QWY�U[�Q��U�Q�e�U�e�e�y�eYu�eY�G�eYW��GY�YV��GY��V�Q�Y�U��Q��U�Q�e�U��e��y�e�u���eY�Yem��  !  ��
��W)�UU�jAU�j �n �nA��U�������������W���V5��]��]���V��Z��k�:鯿:���鿪�鿪������������꫿��Z���V��?�k�:�Z��V�  ��                                                            �����@]��P�ǔ��ǥ����@빪����� pt� ���                   �   ����  "  .��n�Ӯ�F�.���l�^W��ސ?�z�A��9���pn�Wpsk�0n���Х����nz�G�} ��y �W��V��V���V[�UV��_V���������F�U��k@��Z麪Z����u[��_�VU�_U�~� ��5 �� ��  �
  �   /   	             �   �  w     \   �   |      \   �   �   �   �                            �A�  #  ��W��n�m}�k{}�j�r�j�p�j{~��m^����U�CuU��U� �T �   P  ~���� ��� ��_���u�������������������[~U��Wj�U���@������]@�3  3  w  �  �                
      +   /   �   �   �    ��  ��  `�  ��  ��  ��   F   J      (   `   �   �   �        ��  $  �P�����Է ?��@��_�k��?h�  `�  ��   �   �   �   �   i   �  �
  �  �+  �/  ��  �  �� �� ��
 F� �+ `�. ��
  �  (                                                              	
	
	
	
	
  %                                                               ! ! ! ! !                    "#$%"#$%"#$%"#$%"#$%&'()&'()&'()&'()&'()                    *+,-*+,-*+,-*+,-*+,-./01./0  &  1./01./01./01                ��������������������������������������������������������������ﯪ�ꖪU�U�U�� ������Z�ZiVUTQP@�����������UQU 믫������V�UeU��E�fwV3Fwe����R����wW3wW����U��ݪ�U� vUު���Tuݥ�a�owm�o�eݩwJUK�-�UUUUUUUU��U�U��� �U�U�Uժ*tUD  '  U��  tUDUTU���R�t?E@UUUUUUU���fo��V�z�~A목k�k����꪿Un���A� �E������UoA��U���Z��n�����������?�������k�����?�A�������m��cA�����n�z�o�����?��к���m��cA�������?���ᑻ����A�?���꾑k����cA�m䯿����?����o�z���n���~Ay���U�o�f��n  (  ��Uꪥ����k�k��oA�U����E� �A�������nZ���U���  UUUUUUյ-UK�* �U�U�U��� �Uժ�  tUDUTU��  tU��  UUUUUU?u�D�R�R�wDwfwV3Fwew�wU�w�w�wW3wWw�w�Du�ݪ�U� vUު���wJݩ�%�owm�o�aݥ �U�U�U������P@TQVUZiZ������� QU�U����������eU�U�V������믪������������������  )  ��������������������������������������������                                                                  UU  UU  UU  UU  UU  �W  �W  �W   W   T   T   T   T   T   T   TUUU�U=U�U�U�U�U�U���UU��UU��UU��UU��UU��U���U���U���U���U���U�PUUP�UUP�UUS�UU_�U  *  UU�U�U�UUU�UUU�UUU�UUZ�U�Z�UUZ�UUZ�UU[�UU_�UUU%  U�  U� U�
 U�* ���@U���U���U��U�������U���U���U��U���U��� UUU@WUU�WUU�WUU�WUU�W���WUU�WUU�WUU�WUU�W���WUU�WUU�WUU�WUU�WUUT@Wp�W|�WU�WU}�WUu�WUU�WUU�WUU�WUU�WuU�W�U�W�W�W�_�W��W��UWUUWUUUWUUUWUUUWU  +  UUW�VUW�^UW�_UW�_UW�_UW�WUWUUUWUUUWUUUWUUUWU�                U   U   U   U   U   U                      �   �                                                        ������������� ��� ��� � � � �                                  ������������������  ,  ����������                                ����j�㪪�㪪�⪪�⪪jb��������                                ��������������ꩪ�������������                                ���������������������*���
 ��                                ꪪ*���
������ ��*  -   ��
 �� ��                                    @�  ��  ��  �  �   �   �   ��  ��  ��  �   �  ��  ��  @�     �� ���A����?������  � �� �������������� �� �� ��       �? �� �������?���?���??��??<�?? �?? �?? �?? �?? �?? �    ����������  �   .   �  ��� ��� ��� �  �  �  ���������     ��  �� ��? ��?�? ��? ��? ��? ��? ��? ��? � ��? ��? �� ��     �������������������������?���������� �?� �� �� � �    ��?���?���?�?  �?  �?  ����������?  �?  �?  ���?���?���?�    �  �?  �   �   �   /    �   �  �  �?  �  �  �?  �?   �   �                                                                  	
                     !"#$%&    '()*+,-./0123456        789:;<=>            ?@ABCDEF             GHIJKL                    0                                                                                                                                                                                                                        @ P T U     VPe�Z�ZjTU @UUUUQU  �DUD  1  YPB U  �     UE%XU �`             U                                                                    @  	   	  @  AB  !I  "� "�+� +� 7��u
h�v)iMti�O� �     ����h)'� �,9��,9�	'�`�'�/daI�J����'�@.� .�  d             ��
*�"����Fr���z��F~���z��F����������  &�  *           
� �
�`$	���*)h$�
���S��Ɠ�	`��*���Z$�)h�	` 
�     �  ��  �7  p  �
 3k��3��?�����?�[��k� `	  �  �  �  @ `	��#�$d�Z�j&�X%&�X%@&@Z� f  X%  `	  �  �  @ ��:0���3� s� ��ot0���t����t0��o�S�          �  &�  "�  � �{�����3�9�����)i�0)i��k`/�	0� �  @  �(02���������D��F)��'`C��� � � �	 �	                 �  �?  �?  �?  �?  �                                      �  h*  X%  �  �  X%  h*  �                                               �
  Z�  � �@�@�@�@ �  Z�  �
                  �
  Z� �P`P	`$		`$@$@$	`$`$	`P	�P Z�  �
      �
 �Z� ��h @
  	  )  $  $  $  )  	h @
���Z�  �
                    P   �         P   �        @ @       �  P ��_@��@?������7��7���@�@?���_ P  �         �
�
h5\)�*$�$��_&�p��?�<������_ �  �*          P  	 @�j �����h|
e�q!�1e|h�
����@�j  	  P              �  ?� �t���������? �? �����t ?�  �                                          � �W� p�k߽߽5�������V����             � �9 �� �� ��� �����������������:[�V�             ��  l� �� k� ���ZP:�?�?��p:��p:���?�����V�k���                                 �?  _���Op~�4\~�4�w3ӕ73ӗ3s�  P8  |I  ��  ^W  ��  �_  S'  <                                 � � lp		�$�	X+l0��                                            @  �@  �  �>  p�  \��� �  �  |�  �C�          
 ��(�"���*�QZ	j@	hA�*h%X*�
%��	$	h!%j(X&hPi)�������*(
  ��Ͻ�߽��km U{pP��WE���F{��Fnp�G�p�G�p�A�p�ep��p����W���^������[��k���n�\�m�\�m��Ю���S�������[~����knV���z����[�o  �  �>  ��  ���Z�����j�R�~�
��U+��my1�zL�.tW��������ꫪZ���Z_�@�ky�5�y�5����@��Z_Wo�޶����ojk�����F�����^>��z~��y�/4�U 5�P�Q��Q}�QG��Jn�gAY@V@V�V�FV�F   �  �V  ZV �UV VV XV@ `W� ������
�RT)�PU�*PU�
����V/�V��   �
  ��  �� ��5 �k� �[U�VU�V��Z�Υk�����������������������?hP)���?�P:�����������o�����g��_�t��c����Z���N   �  �V  ZV �UV VV XV@ `W� ������
�RW)�PU�*PU�
����V/�V��   �
  ��  �� ��5 �k� �[U�VU�V��Z��k�:���:�������������� G�� �� \�W pA �WG  |S  ��   �   �                            �Vz����@�� y��U�9u����_0bupt�|}p�� 0   0   p   �   p   0���o]�_������O�o4o����G��҇������҇��҇������҇��҇������ڧ�^����v��3w� �v. M�KU��������-H�-���> �               Z�� �j� �5 �A �� �=  �  >                                  �V��V_��~���TպZT5�ZP�[P��@ ��@ �W �V �V ��V  UV  PV   ��������������������k���Z�n�V�o�VU[�_UK�~���5h�����  �
 ��  ����N����ʪ��˫�����n���
���o�o���Z�j�J��K����  K�  ��  k�  [�V��V_��~���WպZV5�ZY�[Y��e ��a �W4�V9�V��V UV PV  ������������������?�k�:�Z��V��VU�_U�~� ��5 �� ��  �
  �      p   �                                                        �֗��S�k�C�W��������[�[��?�?                                                                                              �  ��  ��  7�  7�  �  �  �                                         �   �   �   �   �   �   �   �   �   �   �   �  @�  P�  T�    �?  E�  E�  ��  Ei  ��  Ei  ��  � � �: �: �� �� ��       �� �� �� ��� �� ��� �� ��� �� �� �� �����������                                   :   �   �  �  �:     �     �   0�  �  �� �  0\ r ��q� p0\Wr��qE�pQ�WT? �?� 9��������������*iW*�oW)YU%�WU%FU  TQ%@E% %V �V �� �l� ��
������J���i�������e�l���\UU�\U� �\E �\Q �\T �?   �   @  z  �5  S�  �X 4u @�5 MS� �X�4u�@�5QMS�ET����   �        �����pU%%pU%%p���pU)T�A�B T) �A�  T  �A  �  �� Z�� ��� ��������SI��QI��Q���QU���U��ST��QB��Q)��Q����T��SA��Q����QU�]UmU�m�Pi[�Pi[]B�VW�UUC�UU�UXUXYC�YWAY]@�j5P�V�UE�Uu��WuU]]yUyu]U�u]���W��WU��WU��WT��WT��gdU�gdU�edUu���� �Q� oE� k��j����E�aE�aEꪪ�jU��jUE�jE�j�E�*h�V��jE�jA   �   �   �  ���XXUXXU��Vh�VAh� VA �  A  �  �  �1ݗE��Ѭ��4����A��A��E��F��G� � � ,� x� �  � QVpEVPVVV�V��pVY�pY�V��Zi�k
Ѭ�Ѱ����� �3 l3 l������C���C��՚��u�C���C�w�_p~�G�y�G�w?G�G��W�� ��> ̠> �u�0��QM�?GM���p=pA-pEpQp�p�p� p� p< 0-  0  p   �  �  ��  �_  ��  �5  ��  ��  ��   7   _   �                ��Q���Q�������S}�QM�Q��E�Z}XYM`e���?  V   X   `   �    �j�P�kU��kU
h T
(U�%��IꯥF�T��Q����CV��W��������O��_U]���W�@U� )�oU(��jX���ad���Z�_F�_FE�{P�{Y��륪��j��������E�*�E�Jo������VE��}E�pMQ������4�:p}��M��W�  �:             �  �  �  �  �  S  �  4  _  �   �                       �  �                                                      l l� l�  p~  �_  �   ?   �                                �> 0�>  �. �  �
  �  �   +                                    p  �  �   �   0                                               ��� �F �F �F  G  [�  [�  \n  �^  �  �  �  �C  �Q  �   ��� �� �� �� ��  ��  ��  �:  �:  �:  �  �  �  �  �  �                                                                    @  	   	  @  AB  !I  "� "�+� +� 7��u
h�v)iMti�O� �     ����h)'� �,9��,9�	'�`�'�/daI�J����'�@.� .�  d             ��
*�"����Fr���z��F~���z��F����������  &�  *           
� �
�`$	���*)h$�
���S��Ɠ�	`��*���Z$�)h�	` 
�     �  ��  �7  p  �
 3k��3��?�����?�[��k� `	  �  �  �  @ `	��#�$d�Z�j&�X%&�X%@&@Z� f  X%  `	  �  �  @ ��:0���3� s� ��ot0���t����t0��o�S�          �  &�  "�  � �{�����3�9�����)i�0)i��k`/�	0� �  @  �(02���������D��F)��'`C��� � � �	 �	                 �  �?  �?  �?  �?  �                                      �  h*  X%  �  �  X%  h*  �                                               �
  Z�  � �@�@�@�@ �  Z�  �
                  �
  Z� �P`P	`$		`$@$@$	`$`$	`P	�P Z�  �
      �
 �Z� ��h @
  	  )  $  $  $  )  	h @
���Z�  �
                    P   �         P   �        @ @       �  P ��_@��@?������7��7���@�@?���_ P  �         �
�
h5\)�*$�$��_&�p��?�<������_ �  �*          P  	 @�j �����h|
e�q!�1e|h�
����@�j  	  P              �  ?� �t���������? �? �����t ?�  �                                                �   Z  �U  ZU �UU Z  ����                            �  �  U* U�
UR�UiIU�J UUi�T�   @   @   @   @   @ �
@ �P �������/��/��&���	�V�	�R�	���               �
 j� �� �Z�����W��_��j��kj��W*��W*���                              �
  j� �UT��UTj�UTaiUT�VUTiUU V��                                    
   �   U
  U�  UU
   � ���
  P8  |I  ��  ^W  ��  �_  S'  <                                 � � lp		�$�	X+l0��                                            @  �@  �  �>  p�  \��� �  �  |�  �C�          
 ��(�"���*�QZ	j@	hA�*h%X*�
%��	$	h!%j(X&hPi)�������*(
  ������                                                            �R�W J5~ +�� �T� �R� �J5 �(� ҠT ҰR �0J � ) < �   �         �����������|��l0��l�����Ҽ5�Ҵ6����������{��D���D<��E���E*��k*w�W*w��*}��
y���y��p{�+\~�˜n�s�o�_�k�W�k��j���j���j�+�j��s���\� +W� �� r�� \�� W(� 
� �� �� (� *< "           �   W  k�  �V h� �V�h��?�V��h0�>��x� �> �S� 0N� �8�  �T           �  �  �  ��  � �� ��V�oh��[�V�^h��>�����ݩ>��        �  ��������P���*��U�VU��VG�������E�vQ����F^��        �   �  �  �  P  � �* _����_)����_)����w��w��j   �  ��  _� �� _)���_)�˕��)��2���k-�� ��2 Z� V, �    `  �                                                        �FG�JG��G� �G' �G �XG  X�  Xg  X\( `\�`��*` �b �Z �Z �j����u�t�� y�� v*? q*  �*  �*  �
 ,�
��
��ʿ ��/ �� �� `  �                                                            �C  0  �8   �   �   0   �                                    �:�]U:�]T9�]@5�]4�]0�]�?�^ �^KU�^K��_KS�^KS�^KC�^K�^K�@^KU{��������V�B��K����/��/�V�o���oX��oX��o��oX��o`i�[a�[ai�[u�Zu�Uu�lu�\u��u�����/� �WU�����V��V��V����_���U��2  �  ,  �   2                                               j  h  `  @                              @   @   @��  �-  �  �  n   f   j   j                           ������~�������Q��Q �Q �Q  � �A  � �F  �  t   t   d  �������?���ј�G�����V��V������������ ��  ;�  ,8  � ������������ `� `� `� ��  p� ��  �� ��              �  �� ��� ����������� ��� l�� ����զ�pU����n�������ꦫ���  ��  |�  � ����U�VuU�@������������A���A��zP��zP�zT�ZT�V   � �W pA @: �? O>��@�W7@�U7�U_O_U]CWU�QUUu�UUuM=@�WWEU�?  ���WUpAU:@_:���O���@��7@��7��z]O�z]C�{�Q�^u��^uM��W�^�?   � �U �U: �_: ��� ��?���տ��U���U��zU��{Uկ^UU�^UU�W@�U]�  Z=  �  �� [U��ZU]�j t���_zA�UnA�U�UW�UW�T]�T]�ZPu�ZPu  �   �  �E _E�U_UUUEUU� UU4 U� UEWU�UU����:E��:Ѫ�ꫪ�n����TU�T��@uW{ ��wQKwQ�]Tp�]T�uU {U �EU �  �UU ���U��U�uUUju��j]UUi]PUY]UUYWUUYWUUZWUUV�UUVUU�VUU�VU �VUU�V���WuUEU}UEU�UEUUU� TU�UTU�UTU�UTU��TUEUU�OUUUUUU��UU��_U��zU}��Ut�W~�~}_�z�UZ�UU�U��W�V�W�Y�We��_%��_e��_���������iQ�i@�i@�~U]U_U]UUU]U� \U�U]U�U]U�U]U��_UUU]UUU��UUUUUU�WU��~U���U����yеTkA�QoA�Q�UUE���E�UUE� �EU�FU�U?�UU�UU�[TU�[TU�k W�nU^ծ����꭪�ꫪ��UU�� �U[�UmE�U���U�u4U�U�]U�� UU7 UU7 UU� ���  bWU�`]U�XtU�X�U @W`@]`PuXP�XTiXwT���Q��UG��T��Tu��T���TUGU�W�U�WmU�W}U�_5U�_�U�uUU��W�z\}�z1ԝ~qP�~l���V���j����������5�^}��^��Z_YUiW �e_U}���W�UUU5WUU��UUUU���UUUU����]TU��QUUT @dQ�������T��d�_oUU�oUU�pUU_UU�UUUU����UUUU����QUUUGUUU  �uvԴ������k�eU�Y[ �[}U�[��_\UUUWUU�UUU���UUUU����UU�GUU} PWz�^Uz�zU}�{U]�{UW��UU��U���U}��WWM����wA��T���:�^=�^���z��zU�� UuMU�5U�5��7u�w]��W��5Q��5P%�5@EW�@�U� t� ]�AW��U��TU�QUu�@�ꪪ�ꦪ����������KU��+ ������oU����� �� �T� �� ����� k�� ��? �?  �?  �  �  �  �  �  �  �   �   =         A������j�����P����                                            ������������UPU����                                            ������P����@�����                                            ��z� �:> �z ��  ��  ��  ��  ��  ��  ��  ��   �   �   �   �   �tU�]UE�W ������ZU���������?VU�? �?���WU������ U�? � �?                                                                   @  	   	  @  AB  !I  "� "�+� +� 7��u
h�v)iMti�O� �     ����h)'� �,9��,9�	'�`�'�/daI�J����'�@.� .�  d             ��
*�"����Fr���z��F~���z��F����������  &�  *           
� �
�`$	���*)h$�
���S��Ɠ�	`��*���Z$�)h�	` 
�     �  ��  �7  p  �
 3k��3��?�����?�[��k� `	  �  �  �  @ `	��#�$d�Z�j&�X%&�X%@&@Z� f  X%  `	  �  �  @ ��:0���3� s� ��ot0���t����t0��o�S�          �  &�  "�  � �{�����3�9�����)i�0)i��k`/�	0� �  @  �(02���������D��F)��'`C��� � � �	 �	                 �  �  �  �  �  �                                      �  h*  X%  �  �  X%  h*  �                                               �
  Z�  � �@�@�@�@ �  Z�  �
                  �
  Z� �P`P	`$		`$@$@$	`$`$	`P	�P Z�  �
      �
 �Z� ��h @
  	  )  $  $  $  )  	h @
���Z�  �
                    P   �         P   �        @ @       �  P ��_@��@?������7��7���@�@?���_ P  �         �
�
h5\)�*$�$��_&�p��?�<������_ �  �*          P  	 @�j �����h|
e�q!�1e|h�
����@�j  	  P              �  ?� �t���������? �? �����t ?�  �                                                            �   [  K�        <   �  L=  ,�  �T  �R   K   ,   �   � ��  l� �� k� ��                   =   �  I=  U� TJ=�RE5KU5,U5��T��R� [�                   �   |  �K  |I �KU|I4\I��\U��\U8�_�_��_�      <  �3  |1  W8    �  �   8          � �9 �� �� ���                                                    �   �  ��  _�  P8  |I  ��  ^W  ��  �_  S'  <                                 � � lp		�$�	X+l0��                                            @  �@  �  �>  p�  \��� �  �  |�  �C�          
 ��(�"���*�QZ	j@	hA�*h%X*�
%��	$	h!%j(X&hPi)�������*(
  ��KU KU� UUlTU��QUU�FUU UU lTU �Q� �F�  �  l�  ��  ��   �  �~�ZP:�?�?��p:��p:���?�����V�k���Z���Z_�@�ky�5�y�5����@ �� _���Op~�t\~�t�w3ӕ73ӗ3s�^>��z~��y�/��U ��P��Q�k�Q}��QGk��? �W� t�k߽߽5�������V����Ͻ�߽��km U{P��WE���F{��Fn�����������󯪪^���z[�V������[��k���n�\�m�\�m��Ю���S �U� _U��UU�_U9UUEUU�UU� U9 WE ^� ^�  9  N  �  �   �    ��  �  x  {L  .t  ��  ��  ��  �o  _�  �  �O  o4  �  G�  ���Z_Wo�޶����ojk�����F�����^����v��3w� �v. M�KU��������-H��J�n�mgA�Y@mV@�V�mV�F�V�FWZ����jԬ�5[�A����Ž�ǃ�Z>����G�x�G��A�x�e��x����W��^��G��z���]�W�{A��WG��S��������������[~����knV���z����[�o�Vz����@�� y��U�9u����_0bup�  U;  �m  1�  �  W�  ��  ��  ��  ]�  �  ��  �  o�  ��  ��                                                     �   `      \  ��  ��  ��  ��  ��  ��  ��  ��  ��  S�  C�  �  ��  �  [�  �?�-���> �                                             ��� ��� ��� ��� ��j ��Z �� �� ��Z @k @� @� @V�  V�  Z�  Y����� �� �� �� �� �� �� �� �� �� �� �� ��  ��  ��  t�|}p�� 0   0   p   �   p   0   p   �                        ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  k�  W�  ��  �  [�  �?                     �   �   �   �   �   l  �o��n������Z������� �? ����U�?kU��ZA��Z ��Z ��YA��iU���U�������������������������                            ?   ?   �  �> ��������j_��Z��W                                                   9   �   �     X  h  d  `  �  �  �  �  @               $   `   ��?  �?  �/  �  �  �  �  �  �  �   �   �   9   -                k   �   �   �   �   l   o   �  �  �  �  �? ��� �U� kU��_���kM�:[p��� 5�� ���P��~Y��� ��6�����  ��  j? �j� �Z�����������?�� 9  l9  �?  �� ���.j���VU��UU��P��@�� U�Wp�k=�;�_���kq� �� �� �Z� kkC k�E ��L��p�>/�[�  k� �� ��  �  �  �   �   �   �   �   �   �  �  �  �  �?  �� U�?                                    �  �W  pA  \@  @  @  @  @                                           �  � �� �� ��                                 �� ���������������\��6                                   �   �   �?  ��  � �? �� �                                ?   �  A  5  4  �  �  �  �ZA��Z ��Z ��YA��iU�l�U�l���l����劢�)�����갮�����������o���o���[�8[�Z��j��i��j���j�zК�՚���Z���Z��j��h���������� U^ U
@U�P��UU��UU��VU�^j��
꫾�����z���*�������������������� k�?�Z�?�Z�?�Z���Z{��j���������W�������������?���?���?��� �U�� A�� �� ��A��U��?U��?���?���?���?���?�����������   @  @  @  @  @  @  @  @  @  @  @  T  U  W  �  ��� ���  ��  �� �W= �W��WU=�CUՃ+TU��BU��(T���B���*�������������o�����g��_�t��c����Z���N���N����ʪ��˫�����n���
���o�o� ��  �>  � �� |��W�|U��WU�~U�WU��W(�W���*���������«���  �  �  �  �  �  �  �  �  �  �  �  U�  @�  ?�  ��   �o� �oQ ��A  �E  ��  �>  �   [   �   �   �   �   �  �k  �Z  �Z� ��: ���  �����6���ƀ��R�z�S�A���� ֗� �P���������>P��o�������������������? �  X)  �? ������?�U��jU��ZA��Z ��� �� ���k?�?�������e��j���jk� �_P �>� �ť�����S��>_�E�? A� Q:  �  �  �  �  �   �   �   �   �   �   �  �  �    ��  �  ��  ��  ��  �  ��  ��  ��   �                        ��>�����>  �  �   �   �   �   �   �                           F���Fz��V~���_�& �  �  ��  �  <<  �  �  �  �  �  @  @ ������  �?  �?   ?   �   �   �   �   �                        ��  ��  ?�  ?�  ?�  �?  �?  �  �  ?                             �         \   �                                            �^�T�l��Zm���n��n? �o   �   �   �   �   �                    Y ��YA��hU���U��������������ê�Â��ê����:���>�����?��� �?     @�?��V��Zꯪ�>�� �?                                   �  �   �   5                                                  AB1/00CAB1/01:set8bit
CAB2/00CAB2/01:s2bit
CAB2/00CAB2/01:nb2
CAB3/00CAB3/01:super_vision
CEC3/00CEC3/01:sachen
D527/00D527/01:get_scr_adr
D562/00D562/01:minsert_channel
D571/00D571/01:meffect
D5C8/00D5C8/01:pausemusic
D5FB/00D5FB/01:replaymusic
D616/00D616/01:waitsong
D61E/00D61E/01:mdismusic
D630/00D630/01:mplaymusic
D661/00D661/01:music
D9DA/00D9DA/01:song1
DBC4/00DBC4/01:song2
DD1A/00DD1A/01:song3
DDDB/00DDDB/01:song4
DE60/00DE60/01:rndx
DE8A/00DE8A/01:lr_sc
DEB1/00DEB1/01:rl_sc
DED8/00DED8/01:rl_scc
DEFF/00DEFF/01:d_sc
DF37/00DF37/01:u_sc
DF6F/00DF6F/01:auto_wait
DF82/00DF82/01:push_space
DFAB/00DFAB/01:pause_str
DFB4/00DFB4/01:pr_sprite
E01D/00E01D/01:draw_pic_all
E01D/00E01D/01:prdata_m
E01E/00E01E/01:draw_pic
E01F/00E01F/01:inc_cursor
E05A/00E05A/01:draw_sprite_all
E05B/00E05B/01:draw_sprite
E05B/00E05B/01:inc_sou_adr
E05C/00E05C/01:inc_sou2_adr
E05D/00E05D/01:xor_sprite_all
E0E4/00E0E4/01:xor_sprite
E2EE/00E2EE/01:act_set_data
E37A/00E37A/01:act_set_data1
E3FA/00E3FA/01:power_display_press
E421/00E421/01:power_display_press_inc
E457/00E457/01:time_display
E4D8/00E4D8/01:init_sr
E4F4/00E4F4/01:s5
E5A4/00E5A4/01:init_sr1
E5BB/00E5BB/01:s51
E65C/00E65C/01:over_pic_press
E780/00E780/01:game_over_press
E87E/00E87E/01:babo_press
E983/00E983/01:plan_press
EBC5/00EBC5/01:plan_move_contral
EEDF/00EEDF/01:move_8_direction
EF53/00EF53/01:plan_lab
EFF7/00EFF7/01:print_scoress
EFF7/00EFF7/01:print_scoress1


### symbol table by name ###
0EF3:01:act_bull_fl
0085:01:act_bull_power
0EF9:01:act_bull_us
0EE7:01:act_bull_xx
0EED:01:act_bull_yy
0EE4:01:act_flag
0084:01:act_move_speed
0EE6:01:act_pic
0EE5:01:act_plan_num
0F08:01:act_power_h
E2EE/00E2EE/01:act_set_data
E37A/00E37A/01:act_set_data1
0F07:01:act_ship_powre
0EFF:01:act_xd_set
0EE2:01:act_xx
0EE3:01:act_yy
0016:01:addr
0018:01:addrx
DF6F/00DF6F/01:auto_wait
008D:01:ba_fl
008A:01:ba_index
008F:01:ba_mode
008E:01:ba_onf
008B:01:ba_xx
008C:01:ba_yy
E87E/00E87E/01:babo_press
00B1:01:back_counter
82DF/0002DF/01:back_ground_press
82EF/0002EF/01:back_ground_press1
0023:01:basecolor
090C:01:beat_adj
001C:01:bgbase
02D0:01:bgbuff
0F02:01:buff0
0F03:01:buff1
0F04:01:buff2
0F05:01:buff3
0F06:01:buff4
105E:01:calcul_yn
00AF:01:cheng_mo_pl
C88A/00C88A/01:chk_imp
0014:01:clock
0022:01:color
CAA4/00CAA4/01:colt
C815/00C815/01:cos
105F:01:counter
C141/00C141/01:cur2addr
0010:01:cursor
DEFF/00DEFF/01:d_sc
0ADD:01:data_buffer
0200:01:dbuff
8000/004000/01:demo_press
C73A/00C73A/01:div16
C73B/00C73B/01:div32
C739/00C739/01:divay
E01E/00E01E/01:draw_pic
E01D/00E01D/01:draw_pic_all
0EDF:01:draw_spr_clk
E05B/00E05B/01:draw_sprite
E05A/00E05A/01:draw_sprite_all
006B:01:eff_sel
0928:01:eff_sw
C058/00C058/01:enable_sound
003A:01:enx
003C:01:eny
C558/00C558/01:flash
E780/00E780/01:game_over_press
D527/00D527/01:get_scr_adr
C11D/00C11D/01:home
C79A/00C79A/01:htod24
C8FC/00C8FC/01:htod32
C73D/00C73D/01:htoda
C751/00C751/01:htoday
C739/00C739/01:idiv16
C73A/00C73A/01:idiv32
C739/00C739/01:idivay
C6C8/00C6C8/01:imul16
C67D/00C67D/01:imulay
E01F/00E01F/01:inc_cursor
E05C/00E05C/01:inc_sou2_adr
E05B/00E05B/01:inc_sou_adr
C0AA/00C0AA/01:init_def
E4D8/00E4D8/01:init_sr
E5A4/00E5A4/01:init_sr1
C0A9/00C0A9/01:jirq
C000/00C000/01:jnmi
0EE1:01:key_delay
0000:01:lbuff
C9BB/00C9BB/01:line
C157/00C157/01:line2addr
CA60/00CA60/01:line_45
C889/00C889/01:line_div
C889/00C889/01:line_divx
C889/00C889/01:line_divx16
CA32/00CA32/01:line_xay
CA02/00CA02/01:line_xly
C9D8/00C9D8/01:lj0
C9E9/00C9E9/01:lj1
CA5B/00CA5B/01:lj10
CA2D/00CA2D/01:lj5
DE8A/00DE8A/01:lr_sc
104C:01:m_bull_fl
1034:01:m_bull_xx
1010:01:m_dirr
1004:01:m_fl
00A5:01:m_index
101C:01:m_sida
1028:01:m_sida1
0FEC:01:m_xx
0FF8:01:m_yy
007B:01:mask_addr
0CBD:01:mask_buffer
CAAC/00CAAC/01:mask_c
CAA8/00CAA8/01:mask_s
84FD/0004FD/01:max_plan
D61E/00D61E/01:mdismusic
D571/00D571/01:meffect
D562/00D562/01:minsert_channel
0020:01:mkbase
0FDC:01:moon_bg_move
0F8C:01:moon_bom_numh
0F8B:01:moon_bom_numl
0FA8:01:moon_buff
0FA5:01:moon_fl
0F99:01:moon_gum_fl
0F8F:01:moon_gum_xx
0F94:01:moon_gum_yy
0F8D:01:moon_move_speed
0F8A:01:moon_pass_time
B58D/00358D/01:moon_press
0FDA:01:moon_times
0FA3:01:moon_x
0FA4:01:moon_y
EEDF/00EEDF/01:move_8_direction
D630/00D630/01:mplaymusic
C70F/00C70F/01:mul16
C6A9/00C6A9/01:mulay
D661/00D661/01:music
004E:01:music_sw
CAB2/00CAB2/01:nb2
C66C/00C66C/01:neg_ay
0988:01:old_clock
0F0A:01:old_time_contral
0FEB:01:open_counter
84D8/0044D8/01:open_screen
E65C/00E65C/01:over_pic_press
DFAB/00DFAB/01:pause_str
D5C8/00D5C8/01:pausemusic
0077:01:pic_addr
EF53/00EF53/01:plan_lab
00B0:01:plan_moon_yn
EBC5/00EBC5/01:plan_move_contral
E983/00E983/01:plan_press
0FEA:01:plan_str_conter
E3FA/00E3FA/01:power_display_press
E421/00E421/01:power_display_press_inc
DFB4/00DFB4/01:pr_sprite
C195/00C195/01:prasc
C5B8/00C5B8/01:prblk
C182/00C182/01:prbyt
C580/00C580/01:prdata
E01D/00E01D/01:prdata_m
C18B/00C18B/01:prhex
84B2/0044B2/01:print_moon_p
EFF7/00EFF7/01:print_scoress
EFF7/00EFF7/01:print_scoress1
BB13/003B13/01:print_stage
C17C/00C17C/01:prword
CA7F/00CA7F/01:pset
DF82/00DF82/01:push_space
B9CC/0039CC/01:read_moon_pic_data
0460:01:reflash
D5FB/00D5FB/01:replaymusic
DEB1/00DEB1/01:rl_sc
DED8/00DED8/01:rl_scc
098A:01:rndbuf
DE60/00DE60/01:rndx
CAB0/00CAB0/01:roq
C812/00C812/01:rotx
C813/00C813/01:roty
C814/00C814/01:rotz
CAB0/00CAB0/01:round
0030:01:rx
0031:01:ry
0032:01:rz
CAB2/00CAB2/01:s2bit
E4F4/00E4F4/01:s5
E5BB/00E5BB/01:s51
CEC3/00CEC3/01:sachen
105A:01:score
1058:01:score_kine0
1059:01:score_kine1
0048:01:scr_adr
001A:01:scraddr
0012:01:scrx
0013:01:scry
CAB1/00CAB1/01:set8bit
8000/000000/01:ship_bull_press
C81A/00C81A/01:sin
D9DA/00D9DA/01:song1
DBC4/00DBC4/01:song2
DD1A/00DD1A/01:song3
DDDB/00DDDB/01:song4
004C:01:sou2_adr
004A:01:sou_adr
05F6:01:sound_end
05F5:01:sound_oft
05F0:01:sound_sw
05F1:01:sound_val
001E:01:spbase
0079:01:spr_addr
0290:01:sprh
099D:01:sprite
0A9D:01:sprite_sum
007D:01:sprite_sw
0270:01:sprnh
0250:01:sprnl
0987:01:sprsize
02B0:01:sprv
0210:01:sprx
0230:01:spry
C73C/00C73C/01:sqra
C73D/00C73D/01:sqray
0086:01:stage
0071:01:str_adr
0036:01:stx
0038:01:sty
CAB3/00CAB3/01:super_vision
00AE:01:sys_clock1
0008:01:temp0
0009:01:temp1
000A:01:temp2
000B:01:temp3
000C:01:temp4
000D:01:temp5
000E:01:temp6
000F:01:temp7
0033:01:tempx
0034:01:tempy
0035:01:tempz
0F09:01:time_contral
E457/00E457/01:time_display
DF37/00DF37/01:u_sc
0024:01:va0
0025:01:va1
0026:01:va2
0027:01:va3
0028:01:vb0
0029:01:vb1
002A:01:vb2
002B:01:vb3
002C:01:vc0
002D:01:vc1
002E:01:vc2
002F:01:vc3
C65C/00C65C/01:wait1
C663/00C663/01:wait2
D616/00D616/01:waitsong
C559/00C559/01:wprint
C559/00C559/01:wsprite
E0E4/00E0E4/01:xor_sprite
E05D/00E05D/01:xor_sprite_all
00A6:01:xx
00A7:01:yy
    Qv�.wm  GRAPHICSOBJ           �F�r/  HTOD32  OBJ           �{AN�  IO      LST           ���SE�  IO      O             �r�?N�  C       BAT           �J�>NP   IO      EXT           �d�+v  NUM     OBJ           �Y�En�  GRAPHICSASM           �[�M�  SCREEN  ASM           �Q��I�f  ���x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l���  �U�`LX�� ;�� ��������������� ��L[�`dd� Z��� ��z���Z����� ��z�����`H ;���I���hdi��
&
&
&
&e��e�� �� ��������0����1����`����a�����������������	�����
����������� ����!����P����Q��`����`������`�$�%� 8�$H� �%�h`H�$E$�$�I�i�hI�i ��$$� 8�,H� �-�h`H���,
�-hJH��e-�-hf-f,��,�-`�%E)H$%� 8�$�$� �%�%$)� 8�(�(� �)�) 	�h� 8�,�,� �-�-� �.�.� �/�/`� �/�.�,���-F%f$��.e(�.�/e)�/f/f.f-f,��`````��8��
��i
�$�



$`�$�%��$�tǥ%�uǐ
�%�$�tǅ$8&,&-���,�-`    
  ( P d � � ���@�E�$��ǥ%��ǥ&��ǐ�&�$��ǅ$�%��ǅ%8&,&-&.����`        
    (  P  d  �  �   � � � @ '  N @� �8�Ń�`����	 &� &� � �� Á�� |�Lw��������d���h�� �l��LW����p���t�� �x���������`    �������p����������l��)�D��������0�  ) ��  )����$��d�L̀�  ) ��  )������������������
���������� � ��`�o�`����� ��o��`JJ��������
��̈́��΄�� � ��`�  )���8������  )���e�� ����  )���8儐���  )���e�ɇ���`�������������������������
����������� ����`	  ���ɠ������ ��o������������`�  )�`����G�����`���0��`ڮ���}:����}>����������������`�   ���o����o����o����o����o�`��i������������i����������������������`�������	��i����`�����������}ق����`�� �}��������d�
�ڽ?���@����d ���G���H����dL��� ����������L�ZH A�h ��z�L�`��O���K�!�y�̓u���*+,-*+,-*+,-*+,-*+,-�./01./01./01./01./01�	
	
	
	
	
��"#$%"#$%"#$%"#$%"#$%�&'()&'()&'()&'()&'()���� ! ! ! ! !�                    �                    �                    �                    �``������Ǆ������	�  ��  ��  �*+�45�
��݄�������  �  �L�M�N�O�P�Q�  �  �����@�9�                                                                @� ��� ���A���� ��� ���  �������������� �������������@���    � ��?���?���� ?� ?� ??��??��??��?? ?? ?? ?? ??     ��� ��� ��������������������<��� �� �� �� ��� ��� ���    � �������  �  �   � � � � � � �   �   �   �������� �    ��?�������������������?������������� ��� �?? �      ?���?���?���?�  ?�  ?�  ?��??��??��?�  �   �   ��� ��� ���    �� ��� ����������������� ��? ��? �� �� ����            �P �� ��� @��.����j�y��                             �  OZ �  �� P��j� �                                                            @  ��  ��  �u  �y  ��  �  ��  �n                T   �  �  G+  �  �  �  t  m�� �� J�  �j                                        ��       �  ��~  '� �
�                                             @  �  @* �
 ��                                                  �� mi  �                                   �j  Y�   ����@F `@� X�� ع�                                       i  '
  g  	      �*          �P �� ��� @�  (�  U� @�9   �   �   �   �   @            �  OZ �  �� P��j� ��  ��� jW j)  j  �  �          @�   �   m   �  @  �  �  p@   �   �   �   �   �   �   @    �  �  Z  �=  y=  X<  i>  �>  �>  i?  �  �               `VZ�����9 `�M �� @�� � 8@f   �                            �  [� �� �� �  ܪ ߤ
 u@*  �   @                        �V� U��  �.  �
  �
� V��@i��� �  l  �                                                 
   (   �?  �  (  8   �   �   �    (�� ��� ��  � �� @�* �K^ ��� ��� �	� হ �[> @�  �         ��  ��  @�   �   ��  �  
�  ��  ��  �  ��  ��  ��   �   �   �        �P �� ��� @�  ��  �  �X ��� p�� |�� �)p �  �          �  OZ �  �� P��j� �                                         P  U ����� ��Y ��b @Ub ��i��� ��  �  �                �   +   �R �� ���
Z�j�Y ��Z ��R ��X �� �j  V         
   8   �  �
 (�o� ��J�Z n*V �)e 8�Y (� �% �� �Z �    �  �  �    (  
�  n� n��k���I�J��^���a �j  P  0     0     .�     .�  n� �{��b��b��{���v@*� �V  P       V  �j �� ��X ��R ��Z�j�Y��
Z � �� �R +  �           �  �j �� �% (� 8�Y �)e n*V�J�Z� �(�o�
  �   8   
      P  �j ��a�^��J���I�k� n� n� 
�  (   � �  �      P  �Z @*���v
P��
P��
@��@�� ��  .�     .�     0     0       �     @  @
 �@
�*����	]@ͤ���@
�* �  @
  @     �              �   
 �@	�%T��*9�A3Tj�* � i �@�                               P   $  @ �*��Z���PU��  �*                                       @ �@� � )Tj�*9�A3T��*@	�% �   
  �                                  �*PU���͐�Z�@�*  @   $   P                                           �   �   �   �   �   �  @�  �                 �   * ��� �G��������_/[ �F: �
 9]. {}�                              �?  �?                                                     T  �?   �                                                     T   �  �   /                                             P   P  �  �      /                                         @  @  �  �  �  �  �                                         �  �  �  �   �                                                P   T     �  �  �                                                P   W  �  �                       �                                                            ����Fk Z � { ��+ �%* �O �� ��; ��<   �                                          �  `  P	  �                                              �  p  �9  X%  P  �                                      �  �:  [�  W�  W�  U�  X9  �                                  �   �  \  �+  �  �  �                                       �
  X=  �  �  �   �   $  @                  h)  � ����������F��ê�����*�����
�������� �  h)  h)  � ����������F��ê�����*�����
�������� �  h)  h)  � ������������F����3����*�����
�������� �  h)  h)  � ����������F��Ϫ���?�*������
������� �  h)                              �  �                                                     �   �  �                                                     �   �  �                                                �   �   �  �  �                                         �  �  �  �  �  @  @                                             �  �  �  �                                                  /  �  �  T                                                     �/  �  �                                                                    �   �  �  �C   �               �   (   
  ��  �  �n���N|��n���V��E	�E��Z|��n                � kU+�
  &  P�@kUP �                                  0  ;�  *�  &�  &�  T                                           �   �   p  Z)  p  �   �                                       �   �  [  [  �  �                                              8  �  p  �  8                                        �   `  |  �	  �/   �                               �  ��  �7  `~ |��� w�  �}  �  � �          
 ��8�#���*�	�f�hB�3�4F>�J���b
�R��ME>��`���I���*(
  H����N  �n  �  ��   
   (   �                                    ���0����?�������      �  ��������?0�����                �  �  �            �  �  �              ��� �� �?  �  �  � �? �� ��? �  �  �  ��? 0�� ���    ��� �� �?  �  �  � �? ��  �?  �  �  � �? �����        0  �  ��������? ��  �?  �  �  �              ���0�� ��? �  �  �  ��?  ��  �?  �  �  � �? �����    ���0�� ��? �  �  �  ��?  �� ��?��������?0�����    ��� �� �?  �  �  �            �  �  �              ���0����?��������? �� ��?��������?0�����    ���0����?��������? ��  �?  �  �  � �? �����                                                                     ��D(\� ͰcfeY�}� �Z��Yp9 ���!�� (]�Ͱc�feY}� �Y��Yp9 ��� ��0\� B�c�eY"إ 3X�H@p9�� ��\��@�c�eY� 0X�@@s9 ��  $R  L� @1`  !I @�$  P    ��     �  �@  `Y  !  � @@	  ��           �   �   `          H   F   �  ��  ��  `�  `�  ��  ��i   �   �   �   �   �   �  ��  `��?X�_�k�@� ?��Է���P���� (   � �Q
 `�* �. F� Q�
 �� �� ��  �  �/  �+  �  �
  �                                 �   �   �   �   \      |   �   \  ~�  P �  �T�U�CuU��U�^���~��mp�j{r�j�}�j�}�k{n�m�W���Aݶ]@����@���U����Wj�[~U����������������\��\�����u��_��� ��� �  �   �   /   +      
                �   �  w  3  3                                                                ��   �   �                 ��� pt�����빪���@ǥ��ǔ���P��@]�����z�Gۯ��n�Х�0n��psk�pn�W���A��9?�z���ސm�^W��F�.��Ӯ���n��[n[��_���u�Z�Z�k@���Uz����E����Ѫ���V[�ZV��UV�VV�XVx `W� ��w �ZHM� �� �m� �� ��� ��  g� '����hz�@���+� ��� ������m������� � � � ��`
��
m��� �s����������`�,
� � 8� � 
�@@ 
�S�V}S�( �  �S����@d ��� �� ������ �󩠍  � � � � � � � � � � � �	�& ��"d#� ����/�O�o������멀� �`������_���`� ��@����'� ����0e�� e����`�


 Q��
e�� e�`d
&
&
&
&��
&e��e��@e�`H� |�hHJJJJ ��h)	0�:���H�Z�Z�Z ��z�z�z�h`8� d
&
&
&iN���e�� Z��
 ���� ��� ��0e�� e�z����8��~����`�"�NŅ�#�NŅ	F
�	F	*F	*L�F*F*F
�	F	*F	*L'�F*F*F
�	F	*F	*L:�F*F*F
�	F	*F	*LM�F*F*`        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l���  �U�`LX�� ;�� ��������������� ��L[�`dd� Z��� ��z���Z����� ��z�����`H ;���I���hdi��
&
&
&
&e��e�� �� ��������0����1����`����a�����������������	�����
����������� ����!����P����Q��`����`������`�$�%� 8�$H� �%�h`H�$E$�$�I�i�hI�i ��$$� 8�,H� �-�h`H���,
�-hJH��e-�-hf-f,��,�-`�%E)H$%� 8�$�$� �%�%$)� 8�(�(� �)�) 	�h� 8�,�,� �-�-� �.�.� �/�/`� �/�.�,���-F%f$��.e(�.�/e)�/f/f.f-f,��`````��8��
��i
�$�



$`�$�%��$�tǥ%�uǐ
�%�$�tǅ$8&,&-���,�-`    
  ( P d � � ���@�E�$��ǥ%��ǥ&��ǐ�&�$��ǅ$�%��ǅ%8&,&-&.����`        
    (  P  d  �  �   � � � @ '  N @� �8��@� 5```I�8i@�@�!���"

JJ(�I�i )?��C�(�I�i � `�� `����` 	"%(+.0369<?ADGILNQSUXZ\^`bdfhjlmoprsuvwxyz{||}~~`�)�(�JJJJ�)�
)


8�(�$�
)�J8�)�%�)


�&�)�J�'�e$f,8��jE,.�$e&8�(�,�,� �	e%f,8��jE,�%e'8�)�,�,�8``�|�$�5ɥ%�6ɥ&�7ɥ'�8ɐ�'�$�5Ʌ$�%�6Ʌ%�&�7Ʌ&8&,&-&.&/�����`            
      (   P   d   �   �     �  �  �  @  '   N  @�  �8 �� @ �  5 @B ��  	=  z ���  -1 Zb ������� ��8���I�i���8�	��I�i������������LZʰ0�Z� ��� y��e�8�����e��e � z���`Z� ��� y��e � 8�����e��e�z���`Z� ��� y��e � �e�z���`�"���H� Q��)��JJ����1�h=���` U��0����?```�ɍ& ���  ��� � � � � � �� � �( ����M�F�̅G ѩ@�KdJ�� �J����K�K�`�������� �ϥ)��������)�S����L�Pˍ������W˘ �ˬ��^ˍ�� ���e˘i ����Ll�@@@@@@8  0@P`8@@@@@@p�����Т ��	�
8��
�����p���	�
i�
�����������i����ɀ�L�d�ɴ��  ����  ����`

��̝�̝�̝�̝����i�����
�i��� �	���`	
+,)*78'(56%&34#$12!"/0 -.                   P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������)���`������0'� �	�������
���� Z f�z�����۠ ����	�	�
�
���Z N�z�����ة �`�������	���
� ���� ѭ JJeH�H�Ii �I���



eF�J�Gi �K�JJJJeK�K� )����J���J��
..
..���QH�HȭQH�HȭQH�H�Hi0�H�Ii �I�Ji�J�Ki �K��L��`e���`� ����`H)��,хHhJJJJ�I
eIi@}<хI` 0`��� P���@p��      � �H�@�I��H����I�I�`���	�[�		�
	�	d�	��	���	 �� uҭ
	����	����i<���`

�� ��љ � �����`� �/ ��	��	`��	�
	�@�]�<��8�
	 ѥHi0�J�Ii �K�
	�����J�H���J�Hi0�J�K�Ii �K���
	���  %ӭ
	�a�1�]�-�D Ѣ���HȑH�� ��� �H�Hi0�H�Ii �I��ߩ�	� �
	�_��a�Ș �ѭ
	�a����
	`�
	`�		��		`�	�M�]�I��8�	 ѥHi�H�Ii �I�Hi0�J�Ii �K�	�����J�H���J�Hi0�J�K�Ii �K���	��� %ӭ	�a�1�]�-�D Ѣ�ȱH��H��'��� �H�Hi0�H�Ii �I��ߩ�		�	�a����	`�	`



}VӅJ�W�i �K�J��� ѹZ�eH�H�Ii �I��J�H��`\�\� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �	���ȑ����� ��i0��i ���L\�`��ȱ����	��� ��i0��i ���L��```�	���
������	`��'�����0e�� e��0e�� e���` PAUSE  `

����	� �
��7����BɎ��d

&$
0%�	��!	��	�� 	����i�f
L��Ȟ	�	� 	�!	L)֥	��m	�f
L��``H)��wօVhJJJJ�W
eWi@}�օW` 0`��� P���@p��      ````�)�� �`� ��05�?Z�^ �)�

��) �� �	���	��	��	 <�z�͠ Z�^ �.� �^ �

��	���	� � 	��!	�� 	)	� $�z��@�Ʃ ��`�	�	�	�	� 	�	�!	�	�	)i�	�	)Ji�	�0��d��	�	m	:H����E���h \֭	JJeV�V�Wi �W�	�



eZ�N�[i �O�	J�jJJJeO�O�	)�	�	� �	,	p��N�	��0�� �Nڪ�.���	��	�!	.	.	.	.		.	.	.	.	��߬	�	QV�V���Ve��V�We��W�Nm	�N�Oi �O�	�L��` @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��� �"�!�����  �-� �!�y��-���� �� Z���Iw� z������� ��� S�L��`�������������_^FNNEzz#W4W2Yw� ��� ;��k��څ �٩
��� ;��3��ۅ ���.L�٩(H� � Z� �z�����e�����/����C��/�����`e����.h:м`��� ��.Jjj(**HJ~2~1~0~/J~2~1~0~/hJ~2~1~0~/J~2~1~0~/�з����`            x   �   ?�  ��   ��   �� ��� ��?� ��� aÁ� aÃ� aÃ� Ã� �Ç� ���� ���� ���  ��  ��� ��� ���  ?�  �   �        �   �  �               � ��������  0�                   p   | |  | >  ><>  <><  80  ?0  ? g�� ����� � |p 0w� 8�����~s�  s�  � 8��������g   w   �   �  ��` /�p x<x |x|~ <x|g <y�g�s�c��`��`� � �?  �   �   �    @      ��� 6��	�& ��X����� zũ �"��#�����,��ޅ Sũ����3��ޅ Sũ����9��ޅ Sũ ����D��ޅ Sũ��� ;��  ������ ;��* ������ ;��W 7� |���"� �#�H�e�� e������h��  ����  ���� �� .٩ �"��#�X�Lݭ  )��  )���W��W�  )��  )���W�W�
��W�  )�*���� ;��* ������ ;��  ���  )���X�  )�*���� ;��  ������ ;��* ���  )���X�X�L�ܭ  )��L�ܭ  )��� $���"� �#���H�e�� e������h�� ��@�� JJ����PJJ�	 �թ ��@��PJJ�����JJ�	 \�����)�& ��� ��L��W��� �Z�X���[�Y`�W�����Z�X���[�Y`� �Z�X���[�Y`STAGE: START (C) 1992   Thin Chen Enterprise �  I���H�e�� e������h����  I���`��"� �#����� �	��� � �� �֠� YފH�e�� e������h�`� ����X���� Sũ��� ;��W |������^�
i�


8������� Kǅ������
��������� �թ��� ;���� v�����$ ���% �@��( �7��)  	ǭ�m, ����m- ����m. ����m/ ���, �$ �- �% �. �& �/ �'  �ȩ��� ;��/ �.  v��- �,  v����� ;��X ���
��� ;��= ���0L�ޭ��$ ���% ���& ���'  �ȩ ����m���� Sũ ����I���� Sũ��� ;��/ �.  v��- �,  v�`         





TOTAL SCORE = �***** STAGE    ***** ******************** ZZ22222222PP@``Pp�PP@00@@0@P0P�W�
��W �� #� $� ��)������W����������������������������������������� ���o�� �����������?��^�� �֭]�`�W
��F�G�L6�`S�����S�����S�����S��_����\�_�ţ�`����)���\  ⥤� ��L�� M� �� �� � a�`�\%��^ �Z��[�� 
�������� � ��`�o�`�\�\���o�\`JJ���^ �Z��[��
�������� � ��`�  )��[8奐�[�  )��[e�ɖ��[�  )��Z8奐�Z�  )��Ze�ɖ��Z`�  ) �`�l�o�Y�m�o�R�n�o�K�o�o�D�p�o�=�Zi�[���`�f�l�a�g�m�b�h�n�c�i�o�d�j�p� X�`��lIo��f8��f���
�`}��`��`��  �  ) �`�Y��Y`��r0��`�[�f�Zi�`��r�Y���l�LX�`����[����^ �`��f������ 
��������� ����`��`ɠ��fɠ��o�l���r���f��```������������� ���
��� ��ŧ�`����Ũ�d� �㥮 �� A� �� $� �� � H��`���z����������������������`�����z��������������������`�x��x`�����o�����x�y橥�)�� b�` H� q�`�\#���Zi8����[i8����\d�`��l���`��f� ����`�8���,�8���#�o�l���r�`d�ڦ���������� X�`��i���^ ����������
��������� ��`�o�`����"��������
��������� ���`�o��`����ɠ�����ɠ�`�o��d�d�������`�yŨ���)����y���y`
���������������������l �������������d�d�`��������`��������`��������`��������`������������z������{������|������}������~����`
#A_}�������������z��捏������{��捐������|��捑������}��捒������~��捓����`������������z��捏������{��捐������|��捑������}��捒������~��捓����`��
�����l `�@�g�~������氥�


e� �ɀjiP����


 �ɀjɀje�i
��`氥�

 �ɀjɀje�i
����


 �ɀjiP��`氥�


 �ɀjiK����
��`氥�


 �ɀjɀje�i����

 �ɀjiP��`氥�

e� � �ɀjiP����

 � �ɀjɀje���`�\!�)�/����Z����8���`��i
��`��i��`��L襱L�
�����l *�2�A�I�X�`�o�w襬i	��`��i	����8���`��8���`��8�	����8���`��8�	��`��8�	����i��`��i��`��i	����i��`����������������	����������� �����	d��o�����l�`�r�m�a�s�n�b�t�o�c�u�p�d�v�q�e�w���\�^�Y�P�Z���[�	�o��� ������y��xd������o�������ǅȅ�dĩ��ȅɅ�d�d�dˢ���������������	�]�?�_``���������������������������� 
7&
7   
7&
 
7&
 
7&
 
7
&
" 
7
&
" 
7
&
" 
7
&
"�ų�`�����Ƶ�ƴ�H�e�� e������h�`沥�)�` �� t� �뭻��¢� 6���Ż�d� a� �� .� �� �� ����� X� �� :� s� ���`��������������`��������������`�\#���Zi8����[i8�����\d�`��l���`��f� ����`�8����8�����o�l���r�`d�`��ɖ��o��`���o�`�W
��y�����z�������m����m�������`����i��`��ie�����^���������
��������� ��`���o��`����������
��������� ��`��l���`��f� ����`�8�Ź�)�8�ź��o�l���r�`��8妅���� �����`��03����!�o���H�e�� e������h�`�dLYީ��\� 5쭹�����������L�� i�)��W���o�LK�k�� i�)?Ÿ�`�������	Ɏ���``���`���Ʒ�ƶ`��0`��i���� �ɀjɀji(���� � �ɀjɀjɀji��`���o�`�W�	� � ���W����� �	������� �� ��L������ �	��� ����0�����0�	 �ɩ��p�����p�	 �ɩ��0����p�	 �ɩ���0�����p�	 �ɩ��5�����5�	 �ɩ��k�����k�	 �ɩ��5����k�	 �ɩ���5�����k�	 �ɩ��� ;��W |��W�	���������� S�L���������� SũH��P��������  ���^ �֩��� ;��X ������ ;��] |��� YފH�e�� e������h����H�e�� e������h�� ��@�� JJ����PJJ�	 \թ ��@��PJJ�����JJ�	 ���������� �	���L�STAGE  : FINAL STAGE ������^ ���`�W
���������ȱ��I���`�������������������� ���-�<�X�o������� � �&'()*� 012 �!"#$%�+,-./�  3  �89:;�BCDE�LMNO� 4567 �<=>?@A�FGHIJK�  PQ  �� !"� ()*�  12�#$%&'�,-./0� 345 �6789:;<�=>?@ABC�DEFGHIJ�KLMNOPQ�� !"#�$%&'()�+,-./0�  56�<=>?@�FGHIJ�PQRST�*1234�789:;�ABCDE�KLMNO�UVWXY�����`���� �� ���)�	 �� � ��`�\P��L�Zi8����?�[i8����2� X��o�ǥ��	�����`�����`��	���
��`��d�`���eʅ�E˅˘�̅�&�Eͅ�m  M  e`��` i�ɖ���)��dƩ��ǅ�`���o�t�`��ɠ�	��������`�o�ǩ���`��e�e�i����^ ���o�	�

��	`�Ņ�ƅ��
������� ��`���������	�& ��"� �#� ���� zũ �Z�X���[�Y��	����� �	���������0����ɠ� (�H�e�� e������h�L`�H�e�� e������h� ��L��P� 1�H�<e�� e������h� ���L��)�& L��� ��@�� JJ����PJJ�	 \թ ��@��PJJ�����JJ�	 ��`�� ��@�� JJ�����JJ�	 ��`����  f��  \����� O�L�֩����� L�թ�^ ���`
��������ȱ��I���`����	
 �� $��	�& � �Z�X���[�Y��	��������� �	��������� ����v�d��H�e�� e������h��  I�����ߢ�� ��@�� JJ����PJJ�	 \թ ��@��PJJ�����JJ�	 ����ʊH�e�� e������h�`������
�������2� �թ������������������ �֊H�e�� e������h�L���� ��ͅ�� Sũ����ͅ�� S�`                �  ��%���������	����	���	`�`������������v�����  ?	  	  		 
           	 # $#    &'���  $
00		 
                 $00&'���������  60 "     (   '���  &"   ��                                 �Y���B���  6
		�  	#�  �  
	 	 	

  	 	 	
#  ��  "	"	
	
      		
        	
          	                                         ��6�����  6			
					
		%

"		
	��  #				
���!�b���  				
#($��  2000000 �Hژ���
�h��h��`��� ��H
������������ ����&`l�������� �� �����`� �� �����`� ��( ���������`� �Ν8� ����)�� �
�a� �
��"�� � � �( ����`d� ���!�a�
���(�8����` 6�����`�(t����!�
��L���
�׆ؠ � �ו���������ܩ �ٝ&���߅�����`���`����Lr���������`� �ߥ�m
����
���	���� Lb������υյЅ֦ߠ ��0L!����L$����L=����� ������� ���Յ�m
�� ��L����� ���Ս*��8�*�ե�� ��L�����LD�������}�����չ�� ��L�����- ����H ����H�}����ՙ�֙��h��h��L�����' ���߾��� �՝,�������i�թ eօ֦�L����� ����HȱՅ�h��L�����2����.)��.:�.� �/� ��ը����ߕ�LV� �� ��L������߾��)��.)�.�.�. ����L��ɀ�(逼��

�����,����-����.����/ ����L���߾&�������� �O�� �.� �/�  ��� �ը����ߕ� ����
��Օϥ֕��ߢ�&��&��`���������Lb�� ������ ��L~���� ���Ӎ6��8�6�ӥ�� ��L��

� ���Ө����� ������( ����) ���)�* 	�* Lb�   �����`�����`H���*
�+hJH��m+�+hn+n*��+�*`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   xآ�� �� $� � $� L� �� �� �۩�	�  b� ������ �	�����������d� #��	������\ :���"� �#�  )��v ���x Q������� Q� �թ �"��#�������Յ Sŭ  )����H�e�� e������h��  )����  )��� ��� Q������x Q� �� Z� �� �� �� �֭\�� X��\�o�?�]� $� �� ��L�� $� �� � ��d������� ��O�_����� �	��� � ���L(����������������`� ڎ� M� �������`���� f������������H�d	
&	
&	
&	
&	��	�

&
e��
e		@�	hHJJ�h)����Q��0e���	���Q�`8உ��}���ɠ� i�)i���� i�)��`)




H����)��h��& ������ ������& `l� �������`�������d� #��	������\ :���"� �#�  )��v ���x Q������� Q� �թ �"��#�������Յ Sŭ  )����H�e�� e������h��  )����  )��� ��� Q������x Q� �� Z� �� �� �� �֭\�� X��\�o�?�]� $� �� ��L�� $� �� � ��d �����