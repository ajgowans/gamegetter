     �   `  X	  V% �U� `UUXUU	U�U%W�W9^�^>���?��?��?��?��?��?��?��?��?��?��?��?��?��?��?��?�?�?����� �          @   P  T  U @UU PUUTUUUUUTUUPUU@UU  U �V� �Z��j����?��������� �� ���������?���������  �?  �  �  �           �   �  �  �: ��� ���������������Ѫ�A�z��PPdiAj�j��j��j�ij�i��f�@Z}  i  d  P  @           @   P  T  U @UU PUUTUUUUUVUU%ZUU-jUU/�U�/�V�/�Z�/�j�/���/���/���/���/���/���/���/���/���������  �?  �  �  �           @   P  T  U @UU PUUTUUUUUVUU5ZUU=hUU�U��V��Z��j�������������������?���?���?���������  �?  �  �  �           �  \	  W% �U� pUU\UU	\UU	\UU	\UU	lUU�U�\V�\��\��\��\��\��\��\��\��\��\��\��\��\��p�����  �  �                      @   @   @   @   @   @   p \w7�M�qCp���5�}E��u�}��w�7�_�=i�}��v�@Z}  i  �  �  @           �   �  �  �? ��� ���������?���������i�	�	�	�	h	`	`	`	`	`	`` `  `  `  `  `  @   @            � ��� �`��lk���5���5p�}=\�^?\��?t��?�u�?TW�?T��?T��?���?���?���?������T�� T�? T� �� l�  ;5       :   ;       �   � �7 �� �Y �� ֚5���5py~=\o_?\��?t��?�u�?TW�?T��?T��?���?���?���?������T�� T�? T� �� l�  ;5       :   ;               7  ��  �] �o���5���5pi}=\o_?\��?t��?�u�?TW�?T��?T��?���?���?���?������T�� T�? T� �� l�  ;5       :   ;               7  ��  p] \_ ��5���5p}}=\__?\��?t��?�u�?TW�?T��?T��?���?���?���?������T�� T�? T� �� l�  ;5       :   ;            +   �  �  � @@� @ � @ � C ��@��>��z��:��: ��: ��: ��:��:D��:��:��:��z 0�:  �:  �:  �:  �:  �:  �:   :               +   �   �   �  @� @� @ � C ����>��:A��:��:��:��zA��:��:��:��:��:��:0�z �:  �:  �:  �:  �:  �:   :               +   �   �   �  @�  �  � ����>��z@��:P��:D��:��z��:��: ��:@��:��:��z0�:  �:  �:  �:  �:  �:  �:   :               +   �   �   �   �  �  D� ����>��z ��: ��:U��:��zA��:@��:U��:��:��:��:0�z �:  �:  �:  �:  �:  �:   :          �   �  l  �9 �f� ���lff����f�$�9$l$�$�$�$�$�$�$� $�$�$�$�$�6���������_����  �;  �  �  �   �   �  l  �9 �f� ���lff����f�$�9$l$�$�$�$�$�$�$� $�$�$�$�$�7����������_����  �;  �  �  �   �   �  l  �9 �f� ���lff����f�$�9$l$�$�$�$�$�$�$� $�$�$�$�$�7����������_����  �;  �  �  �   �   �  l  �9 �f� ���lff����f�$�9$l$�$�$�$�$�$�$� $�$�$�$�$�7����������_����  �;  �  �  �       @   �  �  � @jj �ک���������&�ک-jjj/���/���/���/�j�/�j�/��/�j�/��/�n�/��/�j�/���/�j�����j�  �;  h  �  @           @   �  �  � @jj �ک����ݝ���&�ک-jjj/���/���/���/�j�/�j�/���/�j�/��/�o�/���/�j�/���/�j�����j�  �;  h  �  @       �  �  �?  �7  ? @�} �~����������&�ک-jjj/���/���/���/�j�/�j�/���/�j�/���/�o�/���/�j�/���/�j�����j�  �;  h  �  @           @   �  �  � @�j �j��ک����ک&�j�-j�j/���/���/���/�j�/�j�/���/�j�/��/�o�/���/�j�/���/�j�����j�  �;  h  �  @         �5  q�  ]U }U �U: ]�� ]�� ]�� ]�� y�� �� ��� u�� u�� u�� ��� w�� |�+ \� p� �� � �� �� �� �� ��  �  �  �  �   <  �  �U tU �U5 tW� t]�t��t��t��䕺���T�����ԥ�ԝ�ܟ��ݯ�ݫ p�+ ��+ ��; ��> ��? ��? �� ����_             �  \ W �U5 �W� �]��u��ժ�U��U��W�P^�Py�P�P��Pw�p�pw��w��u�  w�  _.  :  ??  �?  �?  �         ?     � @p @\5 @W� @_U@w�@ץ:@W�:@W�:@W�>@^�;@y�:@�:@��:@]�:@��:���:���; �� �� �� |�  ��  ��  ��  ��  ��  �?          ?  �   W �U qU ]�7 m�7 ��� ��� ��� ��� �ڟ �ڧ iڹ �Y� ��� �� �z� ��� �{� ��� �{; �� �� @� @� @� @� @�* @]*  U
  T      p  \  W5 �U5 tU� ��� ����{��z��~�jtj��i��f��Z�������������� ��  �;  �>  �>  5� @=� @?�@?� @}(  T         �  p5  \� W� �U}�V�������j��j�Ъ�	Щ}
�������ky�o���w�����w �� �� ��  ��  ��  ��  ��  Ի  ԫ ԥ P�  @      7  ��  pU@\U@W�@[�@k�7@k�7@��7@��7@��'@��)@�v.@j�/@��-@�y/@��-��~� �ޭ �~� ��. �� �� P� P� @� @� @�  @   ]        @7  @�  pU pU �W5 �_9 �: �: ��: ��: ��: ڧ6 n�) �e* ޖ. ~�/ ޭ/ ~�/ ��/ {� �� �� �� �� �~ �~ �~ �~ �u �U        �  P5  \�  \U �U �W�������������������i
�o�
�������w�����w���� {�  �?  �?  �^  /\  /|�*� *� (}           t  T  W5  W� �}U���p��p�p�p�`��}j�v��[��m��������������� ��>  �>  �>  �  �  �  � �� �Z  Z  P  @   �   U �U �U5 p_� p� ��� ��� �{� �� ؟� h�� ��� ��� x[� �m� x�����z������������� �� �� ��  �  �  u   T       �   \C  WM �Uu pU} �Uw ��u �zu �Zu �Zu �Zm �Z[ ��V �] �k] ��] ��� ��� ��= ��5 �� �[ �� �� �� �� �� � �  �  �      <   � �U pU \U k���u��^��V��V��V�������o��Z��v���7��w7 �w �w �w �� �� �� �� ��@��@�� �� 0              �5 p� \U W��Zu�j]��W��U�U��������m������������������ �] ��  ��  ��  ��  ��  ��  �� @�0 @�   �   �   0   �  p \5 W��U��V��Z�����j��j��j��km�n[��v��u�ow�o�ow�o� �k� �k7  j=  k?  �?  �  �  �  � @�  @�   �   �       @   P  T  U @UU PUUTUUUUUVUU%ZUU-jUU/�U�/�V�/�Z�/�j�/���/���/���/���/���/���/���/���/���������  �?  �  �  �                   @   P  T  U @UU PUUTUUXUU	hUU�U��V��Z��j�������������������������������  �?  �  �  �                                       @   P  T  U @UU �U� �V� �Z� �j� �� �� �� �� �� ��  �?  �  �  �                                                                       @   P  T  X  h  �  �  �  �  �  �                                           �?  ��  l� �U �V9 �[� �o� 쿕 ��� ��� ��� ��� ��� �}� ��� ��� W��e��p���\f�Y�[ff�k���efְ��%�Zf- kY/ ��; �� ��  ;         T  � @�@_�@_�@�@U�@U�@��@U� ��  U�  �*  �;  �+  �;  �+  T:  �*  T:  �*  T:  �*  T:  �*  T:  �*  T:  �:  �
                  P  T  U  �*  U  V%  Z)  �*  �
  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �       �
+ �
+ �
� �
� �
� �
� �
� ��*  �*  �
  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �                          �   �  �  �? ��� �������������������� ���  �?  �?  �  �  �  �  �   �                                                   �   �   �  �  �  �  �?  �? ��� ��� ��������������������  �?  �  �  �                                    �  �  �  ,        �+  k�  [�  [� �[� �[� ��� �� �� �� �� �� �� �� �� �� �� ��/ �� ��  �                      �  W  p  P  |  W  @  @  @  @  @  @  @  @  @  @  @  @  @  �=  $�  	�  	� )�  ��  P=  �                          ��  |U ��5����@���@���@���TUU�UU��}U��MU��MU��MU��MU��MU��MU��tU��PU��@U��@U��@U��@U��@U�� U�; T� @�      � ��
 ��* �jU �ZU�VU�VU�UU�UU�UU�UU�UU�VU�VU�VU�VU�VU�VU�VU�VU�VU�VU�V� VZ	 �U% `U �UU UU  VU@ T�  T
 @�     �   �  �?  W?  ��  ��  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��  �  �  �  �                    P  T  �  �/ @�/ @�/ @�/ P�/ P�/ P�/ P�/ P�/ P�' P�/ P�/ P�/ P�/ P�/ P�/ P�/ P�/ P� P� P�  P>  P  P  @       �  �  �  �  �  �  �  �  �  �
  �  �
  �.  �:  �.  �:  �.  �:  ��  ��  ��  ��  ��  ��  ��  �� @��@��@��@@         P   � P�_ ���]������u�__o���j���o���{���~���k��n���j���~���k���z鯩k��z�����j���~���k���z���k���z���oP��� �� P]          �7W��7    �΄�慇 F��� � J��� � F��` � F��� � J��� � F��` � F��� � J��� � F��` � F��` � J��0 � J��0 � J��0 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������@� �� @� �� ������@� � ���� ���� ��   �� ��� �� ��� �������� � 00�� ���� ��   ,�����,�����������,��� pp�� ���� ��   M�����M�����������M��� ��� ������ �   ��� m��� ��   �   �  � � �   ��09 �   � ������ ���? ��? ������ �   �� �   � �����   � ���: ��: ������ �   ��� �   ������   � ���: ��: ������ � � ��� �   �������� ���? ��? ������ � ��� �   ���� m��� m�   �   �l� � � �m�: �   ��������������   ��� ��� ����� ���� ��������������   ���� �0�� ���� ����� ���� �� ��� ����   �� � �p�� �� � ����� ��� @� �� ����   @� � ���� @� � ����                                                                                                �� �� @� �� @� �� @� ���� �� �� �� ���� ��� �� ��� �� ��� �� ���� �� 0� 0��������,��K��,��K��,������ �� p� p��믫���M�����M�����M������ �� �������묯� ���� ���� ��� � � �� ��L���� 묷� ���� m��� m��  � � �� �뜳��: 묳� �� ���� ������  � � �� �묳 � 묳� �� ����� ����� � � �� �묳 � 묳� ������ �4��� @�� � � �� �뭳��: 묳� ��m�� ���: � m � � l��� ���0�� ���� ����   �~���� G� � ���: ������ �� �����   ��� ���� � ����� ����� �� ��� �   �� ���  � ��� �� ���� �� �@� �   @��� �@�  � �� ��  @��� �                                                                                                � ����@�  � �� @�  �� ���@� ���@� @� � 0�����  � L�� ��  �� ����� ����� �� � p���,���� ���,����� ���,�����,��,�������M��p� ������0�� ���M�����M��M���m �� ����   ����:� �   �    ��l���� p: �<�� @��}���� �� ��  �� �������� � �O� � � ���� ��� ���  �8 ��������  � 듿 � ,�� ����������� p9 ����@� ��  �� � M��<����������� 0 ���@�� � 09  ��l � �  � m���  m�m l �l  m � ������� ������������ � ���� � ������0�� ������  � ������ � ������ � ����� p�� �����   � �� ��  � �� ��  � ���@� ��� ���@�   � @� @�  � @� @�                                                                                                 ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������jUUUUUUUU�������������������������������j        �������������������������������j        ��������뫪�������뫪����������j        ��������뫪�������뫪����������j        ������������������뫪ﾯ�������j        �������ꫪ�������뫪����������j        ��������ꫪ�������뫪����������j        �������������������������������j        �������������������������������j        �������������������������������j        �������������������������������j        kUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUj        k                              j        k                              j        k                              j        k                              j        k                              j        k                              j        k                              j        k                              j        �������������������������������j        �������������������������������j        �������������������������������j        �������������������������������j        kUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUj        k                              j        k                              j        k                              j        k                              j        k                              j        k                              j        k                              j        k                              ������������������������������������������������������������������������������������������������������������������������������������������������������������������ ���  ��� � ��� � ��� ��" ����dͩ�ϩ�Ω �Ʃ��ǥǅťƅ� �����r� ���ǀ�d�ȩ����ǥǅťƅ�dͩ�� �����ɥɅťȅĩ�Ω�� �����D� ��L�� �� ���ǅũ�Υƅĩ �� �i�ƅ� ���ȅĩ�� �8��ȅ� �����T� ��Lކ��ϩ�Ω�ͩL�ĩJ�� ���܍ � �� � �� � �O� � � A٩v� � � � � �2� � �O� � ��	@� � � A���� � �2 ���� ��� `H�Z��
���� ����΅ʥυ˥Ņ̦Ž��нΊ�ѥ�JJ�� %���� �����Ȁ����
�̥υ��L��z�h`H� �� ������h`H�Z�/���� ���� ��z�h`�	�� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                     0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^_____`````aaaaaabbbbbccccc��������i����!� 	� \ 'q 2!"4VDEh��h�ۻ��������������������������쇾�Ez�Fu  Q                            #42#VeVf��w����˽���������������˪��ۘ�������������������������������������������������������������̻��������˻�̻�����������ffvUDC332                          "#324D3DUUUVfgffwwgxwwwx�ww�ww��wwwwwwwwvgwfgvffffgvgwwwwwwx����������������������������˻�������������wwffeUUTDD3333""""""""""""#333DDDDUUVffwwwx���������������������������������������������������������������˻�������������������wwwwwvfffffffUUUUUUUUUUUUUUTEUUTDDDDDDDDDDDDDDDDDEUUUUUUUUUUUUUUUUUUUUUUUUUeVfffffffffffffffffffgwwwwwwwwwwwwwx��������������������������������������������������������������������������������������������������������wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww�������������������������������������������������������������������������������������������������������������g�@�KV�������o���  �   `    ���(���������������@�0���P���������             �PJm�~���������������������ٶ�
p\_��I�P                       ?o�������������������o�u� b        # @(� @          8��������������������������W�B�a       ��<P�R����)"�?��Tf����������������������&�@              $ %Sl������̞��)�50F��X��������������������o�d��Q                @�n��������������������{猃z��4sWRfGA aEf����W�h���v�6Tc�8TFr$&eVTVGC�k���������������������eW2 0            E8GU>���������������z��G��X6=U4q6G�S�xF������G��5K�1b Q3B#5F�$�3xuh�W�EGu�������ܬ��������������ʗ�cU       4!��e�����x���ݚ���������}ּ��ic{e~�3f�uId�X�x�y{v~ۅz�gxw�y����W���ggGde#Ev%dGSTFggtifkhf����������������ۻ���8CfT3$1tTSTGBx%TJe�eewsw�V�xdytxY��������������������tFC3   10SWf����̻�쬺�ʌ����ewFg4r$"%2V2eGdh��z����̽�������ܺ����wVvT%TDER2D32UcU6cxww��y��������w�j��g�w��v������̬����������˪�v�44#       !DdXx�������������껩�v�WwfvdvFvVwgwy��y�j���xvvFwDfWuwV�v�x������̫�˻����G�WeT5DVDFefV�v�����۫�ܼ�ܺ�����xwvfVfwgewffwhvw�f�wx������g�wvh�x���������v�wehdVVeF�Wxv�y��˹���������ۛ��efD3       35Txx��������������ʺ���eeEcED5ETFvfvy����������xx�fuWUeUFfWfWww�y������ܽ��̺������gugeUFeFTTFffxw�x�����˼˻�����wuUUDD3B"""4CUUvx��������������̺���xeUUDB4"31#3DDTVUWvVwvgx��������������˻������x�wudUTDTDDUEfwhh�x���������������xxwgwgfgWgww���������������������������x�x��wfwfUVTTETEDUVffy���������̻�̻�����wvuVdUDDUUCUVVgx��������������y�wvwufefVeffgww�������������������wwfvgfffVfvfVfvww�wx���������������wvwwgwvwwwwxw�w�����������whvfEVUVeeVfwww���������˼������ufUTCDC3DDDDVff����������̻��������wffTeVEEUUUffw�����������������wwvffVeUeUUVUWgxx�����������������wvfeEDUDDDTUEUfvwx������̼�̼�����wfeTD332"#333DEffx�������������̻�����fUTD4333C4DEUVfgw�����������������wwwwvfffffgwww����������������wwwfffUUUUUUVVfffwx�����������������������wwfffffffffffffgwwwx���������������������h��������������������������������������������������SUQc3Cc"c2!!37egVfWWwV�X���{�������TL˨�z�������ٙ����X���wfgSn��d���w�������κ��߻����d~ٶh�{�Ȧ�޼�˽�����ׇ��T�ǆ\�̺��������Ȭ��ʨ���C��u~���ɍ�����������ʻ��uK��e������������ݻ��ˬܼ�T6��Cm��خ��̻��ݷy���d%�ޖV��4Vgu7�Y������w���UuR��S%h��!'t!�R[��c$���c7�bL݇fh��1"�;��s#���C'��D���SFwa��vi��ECc�!J��R&��B9�لW���!!�rj��B$����e8��tz��v4�ۇwy��c3��!8��!jt�cDl�3{��R��V�̧B��R���BL��<��骼�˩�R��U���b~�b���C+���i������#���y���b��!]��s$����쪜�QN��f���t�� +��~���X���z�an��U���P��
����!�욝�߸��!o����� ��%���m�a-�쨧��C����r=�{��!8�1M��$x��1��[�� ���x���Wg1=�����2 ��!��L�1��tu��t
��8��1h1����rEx!=�v�� 
��J����	޶Vv���1��@z����)��14����67�������q80����c&v M�#d�� 
Α [��&�a��Vg��v!����a #ͳ ;ͦ!5� l�qEw��K߁ ���7� M�sF���f ��H��AU�� *��1Fv m�A5gʴ k�1���H�@�wu��e 	޴j��!t�[��W�m�qVv�� [�Q��G�Q	��He���!��)��PG��I��@7�@��f��Aα \���� ��eH��A ��Q���am�!��b����Bwkݣ ��
��Q|�0-��U��� �����1�1��{̨sI�0=�H���1 L� ��6�� ���r6��! l�q���'�0��t����ib��x��$̔ JͶ �� ��dq9��" ��a���9�q	��gG�ܖA ��@���:��S���Ri�l��4Fݶ J�a k������1��0�� 8��1��κ�����x1��Y��1&��	ޘW��܅�A��I��1xޡ8��a(�P	Φ%#��A ����Q:�q [ܢ�� )�a (�����̩�k�م�j��!'ʹ��톇q��G��ai@��E�ʄ�� ��SC[ݱ �Q )ݵ��	��A��R ����a}�A.�ʨg��wb��`���|�Q^������yu�q{��I�p>똹���yf^�j��H̒x��VS�J��!7̵�˚g�ݧUA߷��P��1Nݨ�W��e1��A���Zܢ��Uk�B�u��1��A-�ڕW��dA.�qK��H��^G��T ��1��Z����ez��u1��A$��$��������c�����p���y���eA��(��`��1o�ʧ����f�S)��17��!^�ʨh��vB�Q;��G��1��E��0 
�s)��1&��q����Q�s:��A&�����T}��Q�*��Q%�����e���s����'������w|��t��!���k��+��f6��~�1���h��a��Q\��A���Q%���	��DE����1=��!y�� ^��TI�����!������@���V���A�S=��`h���N��w{���1��@���������v���r��ޱ8~��1��tE���!�s+��QI�����EG�� �]��!y����DY���^��"y�޴��"F����A,��1Y���
��#%���<��1Y�����3F���#�����(���!��a$~�� 1��������@~�#l��1$f� }��0x�����G���$1~�������@��${��@#S�]��!g��o�A%{��U�<��Pg����5}�$R>�������R!��y��axA.�#������t1��!F�� $@n�!������u!��1G���Ut����D��̨0��BW|��!6c-�"���3y��A.�r���25�p߳@;��i���Sn�s7���B6�E�TA;��{���vS��5��ޤF���G!���v����c��dh���Dg�A��b���9���v!��Fy��sT��#���h��s����Vj���z��̪��遼>��f���u���a��bF��Em��!N��wy��vx�u�FS������f!���7���WX��1��tH��#F!^�0&z�"��T4{��vz�﷚��b��SM���z���e3_�!4Z������%���uH�!��C|���V��a>�$���i���wb��bW|�Ft�$:윒z��Ȇf5�݄Y�ʆ3��a�ʂ+���Y���S/�i��!#{s�y3Gܜ����ɖXC��W���ʙ����b���7���BXqn�TX��tUB�U(작W�ܘ�Y���SF���v��a�Y@^��j��6R�2g��aFb�7ی�w���uyS��2X��u���1�XP<��9��CgR.�UI�ˆTe��Q���Fi��wVwc��3j�̵V���A,��I��Dgv϶vuY�R#3.�"L�#f��eT��P��Ey��R5�ʄ���z�ݥVi���vf��QV���~�G���g���vA��s6��V���UVA=�d5���2W�v1� '�܄E���h�� ��uh��4�ژB ��a'�ۓH��n�0Iδv��R�dY��Bh�ܧ4b�S~�Ry��dDd!��BX��bg�� ��1&{˒z�T"�!;��SH��Cz�6�Xh���d�xxb!�D|��Sh�ܗUxx4��V��ܕW�˨d ��R,��Vz��eFT~�BHg��x��do�c��E{ܹfW�t�HX����gxxuA~�@9�ʄ%x��UFd�C$���Ri��vfv"ބ1]�ti��uUyd>�t8f��&U��T2��19̺tH�˗gy��U2��dx��egwS��bYh��%g��e31o�1�ʆF�˘fx�Q>�D'޻�V�ʈgw�d�fs�y��Vi��uU1.�3�˨E���ww��!��s|۬�W���wwvS	�G'���dg���ffs�E%�ʪu�������B>�u;���f���wg�t ��cxw��Eg���WgR�D)���ew��wh��R�vW�z��Ux��UfeA=�TX���Uf��vVwvA<�Vhw��Ufx�wUgvR&�Wfvx�tUwwveffS&�Vfwx�uegwwwwx���w�������������wwwwwwwxw�������wwwwwwwwwwwwww������������������������������wwwwwwwwwwfg��uUGxx��wffh����c���eEevS5Wz�������ܪ�������wwveVffUDDDDD4DC334DC3DVfffgx������������̻�̻������������wwveUVUUEUDDDDDDD33V�fDDg����ww�����z�˙x���x����������wx���x��w�wfg���wgwwwwwwwwxwwwwxwwwwx�w����������������������www�wwwwwwwwwwwwwwwwwwwwwwwwwx��w������������������������w��wwwwwwwwwwwwwwwwwx������wx����������������www���������������wwwwwwwwwwwwwwwwwwwwwwwwwwwwww�������������������9��t�~�ؚ��fEx��w1Fhr  3EeFg�xw����ʘ��������������ܺ�����wwffUUUUDDEUTDC!D343!"#4Ufgx�����������������������ܻe#Vwb3gu$DgC"5efec4fxvwTVx��fx�wg�����wx���w����w�����������������������wwwx�vgwwwvfwfffvfffvfgwvwwwww�����������������������������wwwwwwwwwwwwwwfwwwwwwwwwwwwwwwx���w��������������wwwwwwwxw�������wwwwwwwwwwwwww��������������������wxwwwwwwwwwwwww�www���wwwwwx����������������������������������vww�����������������vffUTDDC3333DEgg��������������x������̼�������xwfeUTDDDUVVfgw�������������˻���wgvfUUED4C3CC3DUVfVfwwf���������������˺�������������wwwfUT3"""#3DEgfwg���������������ܺ������wx��vffeEETC""#5gx���������x����������������������������������vfeT3D2""#EUffffffggwx�������˻��������������������˻�����fUDC332!!"""333DTCEVfvveTTUggx��������������������������������̻���eD"               #Dfw�������������������wx������������������ۼ�����wvfgvfgffeUUEUUffffUDDDC3333"""335UVfgvxwx����������������̻����̻������������������www����������������˺��veB"  ""34DDVfffw���������������̺�������������������̼˻���������fUC2!               ""3Efx�������������ܻ����������������������������������������������vfVUDDT43DDDDDEVffffeUUUUffffggffwwwfvffw���������������������������˩���fffDC#34DDDUVfvfvfffTUUUUfgwwwwvfffgx����������������������˺��weD"   ""#3DEUUUUffeVefVffffwwy����������������������������������˻����vTD3"!           """#"33"#4DDUVeffgwx���˼�����������������������������̺����wweTC"!              ""23DDUUUfgw�����������������������˻�������vfgVUUDD2"  "33433EVx��������������̻��˻��www��vfffvfvfVgwxwx�wfwww���wvw��������������������̻������������wfUDC3"! "35Vfwx���������������������̻���˻�������wfUDC"""""#4DDUTDDDEUVfwww����wx�������������������������ܻ������wffTDDDDUefgwwfeffgwveUC32"#333C43DUUgwwww�������������������˨�wveD32!"#3VfVfw��������˺������weUTDCDDDUVfwx��������������˪���wffDDC333#"#4DDEDDEVw��������������wwvwwwwx��������̼̻����̻�������wwwwfUUTUDC33DDEUgwvfwwx���������˺������wfffgwwww���������������wvfeUDD333332"344Efgx���������������������ܻ��������wwvgvffUTDC""""33DDEUUVUUUDDUUgx����������������������������̻������wwwwvfeUUUUUUD3333333333333CDDEVffgwwwwx�w���������̼����������������������̻��������wwxwvfeTDDDCC3"""!"34DDEUUTDTEVffgw�������������������������̻��������������̻������wfUT3333"""""""!"""334DEUUUfffwwwwvffwgww������������������������������˻�������w��wvwwwwwwgfUTCC33333333333DEUUVffgwx������������������˻���������������������������vffeUTDTUUgwwx���������www�x�wwwwgw���������˻������������wwwwgvffUUUffUfeDDEUVfgww�����������������������������˻���������wwwwwwwffffvffffffwwwwwwx��wwwwwwwx���������������wwvfwwwwwx���������������������������������x��wwxwwwwfffffwwwwwwwwffffeUfffffgwwwvwwwwwwwww������������������̻��������wwwwwwwwwvwwwwwvwwwww����wwwwxwxwwwxwwwwwwwwww�wwx��������������������������wwfffUVfffgwww������˻��������������������������wvffeUUUUUeUDDDDDDDEUTEVfgwx���������������������������������������������������wwwwvwwgvfUUUUUUUfUUUefgww�������������������������������������������������wwwwwwwwwwwwwwwww�wwxxxwx������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������dxآ�� �� c� p٩�X� �� @��  ��dxآ�� �� c� p� N���X O��� p�L��0�����䎖Τr�����	$   �$   �$   ���                        �                        �                        ���            �            �            ��  �0   �0   �	  ��  �0   �0   �	  ��  �   �   �  ��  �   �   �	  �v�t�    ^�^�    W�:�    ���  t���    ����    ����������������������������������������������������������������?<<<300030003000                           ?<<<300030003000                           ?<<<300030003000                           Directional A Directional B Rotational Select control Chimera Pause �  





	
	
			





			

               	$ 	
 "$%()-24=HUNHGC@?=<:9632-*)($ 
   ��  YOU HAVE !FOUND A !YOU MUST FIND A !FORMED A WARHEAD  TAKE IT TO A DARKER ROOM !YOUR FOOD IS RUNNING OUT FASTER!WARNING  RADIATION!FOOD RESERVES RAISED!WATER RESERVES RAISED!UNLOCKED A DOOR:!ELIMINATED !ACTIVATED A WARHEAD AND THE BREAD SUBSTANTIALLY INCREASED YOUR FOOD RESERVES!CONGRATULATIONS; YOU HAVE ACTIVATED ALL FOUR WARHEADS  TO ESCAPE !DARK ROOM NEAR THE BEGINNING!AN ELECTRIC FENCE!A BOX THAT USED TO BELONG TO PANDORA!A TOASTER!A REVERSE FLOWING HOURGLASS!THIS IS A !TORCH!KEY!PADLOCK!SPANNER!BOLT!PYRAMID!PYRAMUD!DARK ROOM!LOAF OF BREAD!MUG!FIND A STATIC OBJECT EXCEPT FOR WATER OR TERMINALS!DOOR!WELCOME TO CHIMERA!CONGRATULATIONS    YOU HAVE SUCCESSFULLY COMPLETED MISSION CHIMERA!DUE TO A MISCALCULATION YOU ARE NOW DEAD!DARKER ROOM WITH A WALL IN IT WHICH HAS A GAP IN THE MIDDLE IN WHICH YOU MUST PLACE THE MISSILE!�ėĠı������%�;�L�Xť�����;�E�a�l�r�v�~ƆƋƓƛƥƳƷ������E�n� 	! &%*
$)-#(,/"'+.0	
 "#'()*+,-./023456789:;>@&=<1 415447,52543554-655, .7454064/55544&% &	
&'	'&		$	/!0 &(		0123456789ABCDEF �  �  �  �     ����     U��0�����?� @��v
�F�F��o/�R"�ʢ|X7�����zdP=+����Ǽ������}voic]XSNJFB>:741.+)&$"                                       ��������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������                                                                  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������  0@P`p��������                																















 @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @�� @��    				



    !!!!""""####$$$$%%%%&&&&''''(((())))****++++,,,,----....////0000111122223333444455556666777788889999::::;;;;<<<<====>>>>???? 0333<???<???<???0333<???<???<???0333<???<???<???������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������           $ ( ,   $(,  $(,      
             " $ & ( * , . �������������������������ڋ������?�?�?<��??<? ?0�������??<?<?0?<?<?<?<?<? ? ?0?<�?<??? �<?<?<?<?<?<?<�?<?<?0?<?<?<? ?<? ? ? ?<� <�? �??<?<?<?<?<? �?<?<?0?<?<�? ?<��??�?� <�? ?3?<?<?<?0���?<?<?0��??<? ?<? ? ?<?<� <�? ?0?<?<�??? <�?<???3?<?<?<?0?<? ? ?<?<�?<???<?0?<?<? ?????<�?<��??<?<����?? �?<��?<�??0?<�? �<??�����<?<                                                ?<�?����?<�?�?�?��        ��UU  UU  UU  ?<???<�?<?<?<? ?  <?<?<    ���<?�UU  UU  UU  ?<�?<� < <?<�� ??<?<    ��� ?�UU  UU  UU  ��?<���?< <?< �?<    �??��UU  UU  UU  �� ?<�?  <�? <?<�?<�?        ��UU  UU  UU  �?<?<�? ?< <?<?<�?< <� �        UU  UU  UU  ��?���?� <������ �    ��UU  UU  UU                            �         UU  UU  UU  H�Z�' J� �֭$ �	J��%  ��z�h@���# `�`H�Z��X� � s׀N�m�m��dm��  I��:��!) ���:)���:)��� �c� H�H�H � 9�h�h�h� ��dz�h@�kH�lH�DH�;H�<H�HH�GH�_H�`H c�h�`h�_h�Gh�Hh�<h�;h�Dh�lh�k`�����`�EH� �إ �آd3d43&4 &��e3�3�e4�4���4�3h E؆4�3`� � ����`� ��`
� ��e � �i ��� �� �� �` ��l  � Z� �� � ���� ��0	��z��L��`Z� �_�a����_�a�`�b�0	��z��L�`	 I�i`H� E�h`H�I���I�����h`�e � �`�`�e��`�`�e_�_�`�``e;�;�`�<`ea�a�`�b`H� I�� �I��� ��h`H�I���I�����h`� I�� �I��� ��`�� H�H�9H�DH�� d �۩  A�h�Dh�9h�h� ``���H�^)�^h




^�^�& `H�Z� ��  	 � �� � ȱ � ȱ � ��� z�h`dd�d��`x ٩�X` cٜ � � � `� � � � `H�Z� H�H� � �@�� �  ��h�h� z�h`�k�ldD�
&D
&D
&D
&D�;�D�<�;
&De;�;�De<	@�<�JJe;�;��<ڊ)�D��+ɅH�C�'�%H�G�D�`�{�G�a��a`�[�<�A��A`�:��0��`�.��$`�,��%`�'��&`�"��'`�?��(`�!��)`�`��H�Ӡ� �׎�h�	i


����\�,�� |�� ��Z ��z��m��\��]LW�H�m�h�`lH �٩ ��h �٢Ӡ  �טi �_�i��`�D
iʅ��	��9�	� ��_� � ;�;�� ������;�;�;i0�;��<�_i0�_��`�9��`H �٩  ��h� �
���_��`� �٢ӠH �טi��_�iӅ`�D
iʅ�9H��	��9�	� ��_� � �;�� ������;�;i0�;��<�_i0�_��`�9��h�9`�� �_�;�;��<ȱ_�;�;i/�;��<����`�:)H���H����Z�[h`� ����Z �٢�
� �;���;i0�;��<���z���9�9HZ�.*.*.*.*)������ ��hzi�h�9�9��`�:)����:)���`�d�
I|�I5�	�I�` �٥G�;`�;H�<H�eDiJJ�
�
ڦD�/�I��heD)��3�I��	��� �;%�;� �
�ȑ;���;%	�;�;i0�;��<���h�<h�;`�Z�;H�<H�	�eDiJJ��ʆ
�Ʌa��b� �;�aȥ<�aȥ
�aȥ	�a� �ئ	�
�;�a���;i0�;��<� �����h�<h�;z�`���;���<���
����	�ͅ_��`�	�
�_�;���;i0�;��<� m����`�;H�<H��D�+�I��	��;%	G�;�;i0�;��<���h�<h�;`��eDJJ�	�D�/�I�2;�;�C�'�=/�;�;� �C�'��	��;��	���eD)��3�I�1;�;ڦC�'��=3�;�;`�����k���l��� iݭ�m�8���� �ٮ�� iݮ��� �٬� 9ݬ���m�8�� �٬�L9ݩ `��`�چn�
�o�7�-�I�o�pq�A�oix�� � ���0�n�7�-�&�o�xy��n�0�o�p,�p��q)�ߠ" �׀Ѐm)����
I

��@�  �߀TH�n�	��h}���I

�ڹ@ɝ ��ɝ �oip� ��ڦn�)� �ފ�o�x�y�	@�� �n�	@� ��0L�`H� � �ס �  ��he � ��)�Ff Ff Ff �n�)���� `6�6�7���G�rߏ߹��ߩ�`�n
ip�� �n�L�צn�7�I�-��� � c��� V��� ���( `�)������ Sٜ �( �`�oip�ڦn�)� �ފ�o�x�y`�o�p�p��q�n�`�oip�� H �ס � �ס  �ת��h`hL٭8�


eo��o����p ����q �n�`���� Sٜ �( �* ��Lr�


�� ����p ��������xty������������` pٜ � ��\�Å]��� 0ک�\�Å]��8�  0کޅ\�]�(�P�  0ک�\�]�(�`�  0ک��\�]�(�p�  0ک  ��d���P�� �:���:��)��8�:)@��i��� ��  ��ͥ:)�����e������Ņ�  �����ک  �h`�k�l��� ڦk�l �٢�� hH�������`�_ qۥli�l�����`� ��:)��`�  �� �à w�  �إ:)����:)���� L�܆]�\� �\�����



�E��8�EJm�H8����i8�Z �٥Ei�ڠ  �� ?ܩ�C��  ��hi���L0ڜ"�#d&d'd%��������������������������1��2���/��0�(�-�#�.����)�$��#��$��"����� ������?�����O�������;�CȨ��ș���ș�� j�� �ة �_���`���a�V�b�(�'�_�a���( mة0 �����  �ة�  ��U�T�_�k�t���r � �� G� �� E� �歩���$�$��� �  ��/i-� �0e.� & &� m"�"�m#�# ��2 A٩  �ة  � A٭���� A٭  I���L"��   ����N ٩����!�  ��� [� A����� A٭���L"�� �;�@�<�x�'�; z�;���0 x����`څ�d	� FjFj�8�@F	F		�	���	�`��dd	d
�&��e��	e	�	�
e
�
����� HJJJJ	0���h)	0���歼�0�� ��`ι�`���8�-��-��.� �.�0. �� Q������8���8�/��/��0� �0�0 ��Lp� �  �� Q�L%� �  �� p�L%�x�� �٢(� ?ܩ��\��]�x��� L0ڢL�� �٢(� ?ܩ��\��]�L��� L0� �٢ � � �� �;ȱ �;ȱ �;ȱ �;ȩ, x����`� �;ȑ;ȑ;ȑ;ȩ, x����`������������`��+���,�����+��,����$��� ���� � �� ������ � � �+��,� ���� � �+������+`8�
���ǅ ��ǅ� � �+��!����e+�+��,�L%孮�`���2��� ��γ�%����1���� ���1��2�1�������1��2`�^�[�~�[���^�[�~�[���^�[�~�[���^�[�~�[���^*\�~*\���^*\�~*\���^Z\�~Z\���^Z\�~Z\���^�\�~�\���^�\�~�\���^�\�~�\���^�\�~�\���^�\�~�\���^�\�~�\���^]�~]���^]�~]��`�#J8� 2ت�$J8� 2ب�H�yHĢ��0	�O����j�`� `Ψ�����\�9����9��
`�9�\��`���\`�9�\ b�� *�	8�-��-�.�	�.������� L��DFFFFFDF     FF     FF     FF     FF     FDFD DFD @@" "@@"            ""            ""      @00 00@ @`@`@`@@     @@      @`@`@`@       @`@`@`@@`@`@`@ d     dd     d@     @   @  @@  @  @`  @  ``  @  ` 	
@ @G@GD@     @@     @@     @G      D     @DG@G@G@                            PPP PPPP     P�     ��  w  ��     �P     PPP���PP 44444444      4      4      4      4      4 44444                                  		  C  C  C     C     C     C     C     CCCC 
'G     G             G  @@@@G      G       G     G 	EEEEEEE  @E@  E ��� @E     @E�����@       E@@ @@@ HhhhhhH       H`````HH      H     H      HHhhhhhH  � � �       � �       �   �   �   �   � � �      G0G G0G0     0G     G0      G     G0     0G0G G0G DGG GGD      D            D            DGGGGGD DDDDDDD  @   @  @   @      @  @   @  @   @DDDDDDD """"    "           "         """" U@U U U@   @ @U   P P@  P@ @U  @  P@  P  @U@ @ @P  D f  p  f  p  f     f  p  f  p  f  D   H  H  HH  H  H   @  HH@@@  H      HH     HH@@H@@H f"f"f"f"     "f      "   "f"f      "     "f"    f �� � ��   �  �   �  �����         �      �������� �������� �   �� �   �      �� �   �� �   �������� xxxxxxx              xxxxxxx              xxxxxxx  D  D@@D      �      �D���� �      �      �D@@@@@D 
D      D                     $d$d$d$                 ppp               $d$d$d$ 3333333  0   0  3   0      0  3   0  0   03333333 U U         U U         U U         U U   UU p    U p    U ppU UU     UU     UUUUUUUU W W W W    @      @  GGGGGGG              PPPPPPP % !���       �@�@�@ �@�@�@��@�@�@        ��� !!" 3`0`0`3        p0p0p0tp4p4p4 p0p0p0       3`0`0`3 ""#!@@@@@HD                 @HHD              @@@ @HD #)$"DHHhhhDF`     F`     F`     F`     F`     DHHhhhD $$$#GGGGGGGW      W      W      W WWWWWW W   WG G G G % %&UUUUUUU  P   P  U   P      PU U   PU P   PUUUUUUU &&%&Cp p pC   p  �   pp �      �      �      �C�����C ('
'D"3UD"3U  U  U3  U  D"  U  "D  U  3U  U  U3" U "D ('((D�D D�D�     �D     �       D     ��     �D�����D # *<D     D     DD           DD     D      + )"  "  "                    "  "  " *,  5  5  55  5   5  55555      5      5      5555555 +  -DD DD       D@@D                     DDDD . ,/DGGDGGD  D    @                 DGD DGD  -  DgDgDgD      gDgDgDgD      g      D       DgDgDgD   -0�T�T�T�U      U      U�� ���U             �T�T�T�   /1��             ��                �� 2 0; f"f"f"f      " " " "f      "      f      "f"f" "  1 37 7   7      d7d7   d  d   d  d   d  d   d7 7   7 4;2 EpppppET      E ppppET p    E p    T p    E E   E  3 5aaaaaaa       a`a`a`a  A A                DD DD  647" "                     5         � �   � �   � �   � �      85 P P P P� � � ��   � �� ����P� �    � �    P P     79  W WWWWW      W     W     W     W     W    WW      8 :  ff"`` f      "D         D  "D     f      "ff"``    ;9    $     (    $             $      ($($($($ 3 1:UEEEEEUE  E  @E  E  @   E   E  P  @E     @U@@ @@U  =)?@@@ @@@@     @@     @0      0     @0     @0000@@@ <  >                 0     03      0                  ? = ���PPPP��P    PP    P   p  PPP   P���P P����P P��  ><@`````      ` `    ` `  0 ``  00 ``     ` `````    ?  S٢?�%���$ ���5� �%���$ʽO�V���\��[�0�%�șe���[�ȍ� �� ���V���	���  ��\��`�[��Í��č�`� � Jv 	��`�\0�8����)���)�\�V� � � � � � � � � � � � � � � ��Ӡ � � �Å!Z̛��\0	�:��9 #�hH�)� ��zZ�eJJJJ /�zZ�e /�z��1�ɢ� ��A� ��A�@��A�`�B���DB���tB����B����B� �C� �4C�@�dC�`��C����C����C���$D���TD� ��D� ��D�@��D�`�E���DE���tE����E����E� �F� �4F�@�dF�`��F����F����F���$G���TG� ��G� ��G�@��G�`�H���DH���tH����H����H� �I� �4I�@�dI�`��I����I����I���$J���TJ� ��J� ��J�@��J�`�K���DK���tK����K����K� �L� �4L�@�dL�`��L����L����L���$M���TM� ��M� ��M�@��M�`�N���DN���tN����N����N� �O� �4O�@�dO�`��O����O����O���$P���TP� ��P� ��P�@��P�`�Q���DQ���tQ����Q����Q� �R� �4R�@�dR�`��R����R����R���$S���TS� ��S� ��S�@��S�`�T���DT���tT����T����T� �U� �4U�@�dU�`��U����U����U���$V���TV��L|�`�\�  ����H� i� �!i �!h)�`8��  ��� � i �ȱ i��8� ����� �
� � ��=�� �ȱ ��=�� �ȱ ��=�� �ȱ ��=�� ���i����
н`ڪʥH�H� d�6�� � zטi� �i�h�h��`�#e$J)i��#i8�$��(�� e%��'����I��




��'

e%e"�  ��Lh�               ����L����-��&���()�L"� P���L��)�L���)��'��'L"���&���()�L"� P���L��)�L���)��7��'L"���&���()�e P���	����L��%(J�!����'�')�'������R� ���L����J�!����'�')�'������V� ���L����J�L���%�#JJ����R����V(������&�-� ���� ٥%i���'���e#�#���e$�$� �%L���'�#����Y�$d%��#Lj������Z�$d%d#Lj��$����W�$d%��$Lj������X�$� �%�$Lj� F���%JJJJ�L���[��\��%� ���� �L��JJ�L���$J�


8���#Je���)��#J��$J�� �e%�&�$J��)i�)�#J��)�)�ȅ)`���'��}B�`� �:�)���)���)���)���) ��``H���\h`�/i܅/�0i�0�� �  ��`�-i܅-�.i�.�� �  ��`�   ���Z� ٩( ���) ���* ���+�\ ��Ly��d d�>��  ��hm"�"��#��| �� � *�L���#�" ��,�� �٢ � ?ܩ��\��]�,��� L0ڮ$ʭV�O�\���[�`�Vɠ�L���U�`���8�`����`�  ੠�V�8�\������� ��������� ��	���  ���/ią/�0i	�0�>��L��.=44544������������`���`hhL��L�� ���  � A����L�� F��[��\0��5��� y���  �� x��5�
L���4��� y���  �� x��4�L���-������ �� y� x��-�KL����L%��8�L���6��7���  ��L���,���  �� y��>�L���8�9��L%�H8�.������� �� y� x�h���KL�� F�����[��\�����5�,�)�����
� �� ���4�\�5�L�� ������>L���4� ������>L���)������/�L%��
� �� ���/�L�������3�L%��
� �� ���3�L�������0�L%��
� �� ���0�L����4� �� y����L����5� �� y����L���8�9��L%��6��7����3���	�  �� ����3L���,�% y����8��"�8�-�������  ��
��L�����-��V���V��� ��8���dL����J���8�,��L���L��JE�L%��� �� y��8���dL������� ��`���  � � � ���#  S٩����& �^`� � ����  �ע t ���`����������������������������������������������������������������������������������������������� ���