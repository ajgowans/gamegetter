UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���������������������������������������W�                                      W�                                      W�            ��?         ���           W�           �WU�        \UU+          W�           pUUU        WUU+          W�           pUUU5        WUU+          W�           \UUU�        WUU+          W�           \�WU�
       WUU+          W�           \�_U�
       WUU+          W�           �^U�
       WUU+          W�           ��^U�     WUU+          W�           �*WU�
       |UU+          W�            �UU�
 <     pUU+          W�            pUU�
 �    pUU+          W�            _UU�
 �    pUU+          W� �0<��  �UUU� ��   pUU+   ?��0  W� 3�0�0   pUUU�  ��U� pUU+   �3�0  W� ��0�<�  \UU�+ �U�UW� pUU+   ���?  W� 0�0��3   \UU�
 �U�UU� pUU+   ?�0  W� 3�0� 3   \UU�? �U�UU� pUU+   �0  W� �0<��  \UUU�
�U�U}� pUU+   ���0  W�           \UUU�
�U�Uϵ pUU+          W�           \UUU�
�U�U˵ pUU+          W�    00   \UUU�
�U�U˵ pUU+   ����? W� ��   ��   \UUU�
�U�U{� pUU+   00�0 W� ��� ���   \UUU�
����� pUU+   00�0 W� ��   ��   �����
 �
��� ���+   �0�� W�    00   �����
       ���*   �0�0 W�           �����
       ���*   ?0�0 W�                                      W�                                      W�                                      W���������������������������������������WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������W�                  p5                  W�                  p5                  W�                  p5                  W�                  p5                  W�  �?<�?�       p5 �?������<��� W�  ��<���?�       p5 ���?������<��� W�  ��<��<<�       p5 ��<<�< ��<�� W�  ��<��< �        p5 � <<�?���<�� W�  ��<��< �       p5 � �?����<�� W�  ��<��<<�       p5 ���� ��<�� W�  ������?       p5 ��<?������<��� W�  �?��?�       p5 �?<<��?���<��� W�                  p5                  W�                  p5                  W�                  p5                  W�                  p5                  W�                  p5                  W�       ������?��? p5                  W�       ������?��� p5      ��         W�       ����< �� p5      pU         W�       �������� p5      \U4         W�       �������� p5      k4         W�       ���� �? p5     ��4         W�       �������� p5     ��:         W�       ���?���� p5     �j :         W�                  p5     p)�<         W�                  p5     p �         W�                  p5     ����?        W�                  p5     �����?       W�                  p5     p��'X�       W�                  p5     p��%V	      W�                  p5     Le��V      W�                  p5     SeUU�      W�                  p5     WYUU�0      W�                  p5    �TYUUe�      W�                  p5    �TYUUeU�     W�                  p5    0T]UU�V)     W�                  p5    LUUU�Z0     W�                  p5    S�pVU���     W�                  p5    W5�V�U�U�     W�                  p5   �V�Z�V9�    W�                  p5   �h��jU50     W�                  p5   ���ZU��*    W�                  p5   ���������    W�                  p5    ��? �����    W�                  p5     0?U�����    W�                  p5   ���*����     W�                  p5  �PU���       W�                  p5  ��<"��V      W�                  p5  ��� ��Z      W�                  p5    ����j1      W�                  p5    ����f1      W�       �?��?      p5     �����f1      W�       �ʫ��      p5     �?���j1      W�       �ʫ��      p5     �����f1      W�       �ʫ��      p5     �������      W�       0�<�      p5    ��?�����      W�       �?��?      p5   �?�?�곾�      W�         �       p5  ��������      W�         �       p5  ���������      W�         �       p5  ���������    W�         �       p5  ����������    W�                p5 ���������?L    W�         �       p5�� �������0   W�                  p5�? �?������   W�                  p5�? ?<�����+   W�                  p5�?��|�����Ce   W�                  p5����������   W�                  p5@����������   W�                  p5@�����������   W�                  p5 ������������W   W�                  p5 ����������?��  W�                  p5 ���?���������   W�                  p5�����?���W<   W�                  p5���<������@   W�                  p5@|������?    W�                  p5 ���?�����    W�                  p5 ��������?   W�                  p5 ��� ����V�� @  W�                 �s5 �<  �������  W�                 �|5 |_   ��������  W�                 �|5 ��  ��������  W�                 �|5 �����������/ @ W�                 |5 ������������  W�                 �s5 �� ������?0��   W�    �?           �s5 �� �����?���  W�    ��           �|5 ��� [����?Z��  W�    ��           �|5  �����  ���h5�  W�    ��           �|5  ��U�  ������  W�    0�           |5  ��]�?  ����Z�  W�    �?           �s5  �U�  ����Z�/  W�   ��?�         �s5  ��w�  0���k�?  W�   +�ʫ         �|5   ���   ������?  W�   ��ʫ         �|5   � @ ������?  W�   ��ʫ         �|5      @ ������?  W�   <�         |5        �����7  W�   ��?�         �s5        ����p  W� �?��?�      � �s5     @   �� ��}  W� ��+�ʫ      � �|5        ����7 W� �ʫ�ʫ      � �|5       @ �� ��  W� �ʫ�ʫ      � �|5         ����  W� 0�<�       |5         ���? W� �?��?�      � �s5         |���? W���? �?��?� �?��?�s5         ����� Wի�� �ʫ��+ �ʫ�ʫ|5         @�����@ Wի�� �ʫ�ʫ �ʫ�ʫ|5          ��� Wի�� �ʫ�ʫ �ʫ�ʫ|5          ��_� W�<�  �<� 0�<�|5          �ǥ�  W���? �?��?� �?��?�s5           ���   W���?��?��?   �? �?�s5           ��?   Wի�ʫ�ʫ��   �� �ʫ|5           ���   Wի�ʫ�ʫ��   �� �ʫ|5            �   Wի�ʫ�ʫ��   �� �ʫ|5            �    W�<�<�<�   0� 0�|5                 W���?��?��?   �? �?�s5                 W��������������������������������������WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ����������������������������������������                                      �                            �  @QEQEQEQEQEQEQ  @DDDDDDDDDD �  PUUUUUUUUUUUUUUUUUUUU    �  T                      @D�OO�O��tD �                         �1�1� �  �
���*�* �����  @D�tO�tO�GD �  � (
���  <<<<<<<<<<   ��1� �  � ( 
���  <?<?<?<?<?  @D�tO�tO�GD �  �
( 
�*�
 �<�<�<�<�<   �1�1� �    ( 
�"�  <<<<<<<<<<  @D�O��O��pD �  � (
���  <<<<<<<<<<    �  �
�����* �����  @DDDDDDDDDD �                         ����?� �  T                      @�tO�tt�DOG �  PUUUUUUUUUUUUUUUUUUUU   �1�1� �  @EQEQEQEQEQEQE  @�OO�Ot�O�D �                           �1=1� ��������������������������@�tOw|t�DOG ��������������������������
 ���1�? ��                        
@DDDDDDDDDD ��                        
  ��                        
@DDDDDDDDDD ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@          ��                        
@          ��                        
@  �
��  ��                        
@  � ((  ��                        
@  � 
(((  ��                        
@  � 
(�  ��                        
@  � (   ��                        
@  � �(   ��                        
@          ��                        
@          ��                        
@�������                        
@<<<<<<<<<<��                        
@<?<?<?<?<?��                        
@�<�<�<�<�<��                        
@<<<<<<<<<<��                        
@<<<<<<<<<<��                        
@�������                        
@          ��                        
@          ��                        
 UUUUUUUUUU ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@          ��                        
@          ��                        
@��*(�� ��                        
@�� (
� ��                        
@�� (
� ��                        
@��
(�� ��                        
@�� (
� ��                        
@��  
� ��                        
@���*� ��� ��                        
@          ��                        
@          ��                        
@   ��   ��                        
@   <<<<   ��                        
@   <?<?   ��                        
@   �<�<   ��                        
@   <<<<   ��                        
@   <<<<   ��                        
@   ��   ��                        
@          ��                        
@          ��                        
 UUUUUUUUUU ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@          ��                        
@          ��                        
@��
�* ��                        
@��(
�� ��                        
@���
� ��                        
@��(
� * ��                        
@��(
 � ��                        
@��(
�� ��                        
@���
(�* ��                        
@          ��                        
@          ��                        
@  ���  ��                        
@  <<<<<<  ��                        
@  <?<?<?  ��                        
@  �<�<�<  ��                        
@  <<<<<<  ��                        
@  <<<<<<  ��                        
@  ���  ��                        
@          ��                        
@          ��                        
 UUUUUUUUUU ��                        
            ��                        
            ��                        
            ��                        
            ��                        
            ��                        
 UUUUUUUUUU ��                        
@��                        
@DDDDDDDDDD��                        
@��                        
@        D��                        
@�
**�*��                        
@

 (
�D��                        
@*
  ���                        
@�
  �D��                        
@

� � ���                        
@

  �D��                        
@

  ���                        
@

 (
�D��                        
@
�
**���                        
@        D��                        
@QUUUUUUUU��                        
@        D��                        
@�?�?�?�?��                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@������                        
@�?�?�?�?D��                        
@�?�?�?�?��                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@�ʫʫʫ���                        
@�ʫʫʫ�D��                        
@������                        
@�?�?�?�?D��                        
@        ��                        
@DDDDDDDDDD��                        
@��                        
@DDDDDDDDDD��                        
 UUUUUUUUUU ��                        
            ��������������������������
            ��������������������������            �                                      �                                      �                                      �                                      �                                      �                                      �                                      �                                      �����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<3<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  ��V�V�V�V�V�V���??��??      �    �              ��           �v�      �3� 6                                  ���������������������~����������                           � ����������������������~����������                                ffff���$"�f�Eb%b����Yb)"�����   �   �   �   �  ��  ��  ��  �� ��? ��� ��� �����?��������������?�����:������?�� ��: �� �� ��  �:  �  �  �   :               ?   �   �  �  �?  ��  �� �� ��? *�� ���������?�*����������������*� ��� ��� ��� ��*  ��  ��  ��  ��   �   �   �   �                                ����������������!!!!HHHH�������������������� ��� ��� ��� ���  ��  ��  ��  ��   �   �   �   �*� �� �� 
� 
� 
� 
� 
� �� �� *� �� �� 
� 
� 
� UUUU��ZUUY` Y�Y� Y� Y�
Y�*U�*�V���Z"*V
�TEUY��ZUUU                                 ?  �� ��? ��� ��� ��� � ��  UUUU���ZUUY  Y
Y*Y�
Y�Y�Y(HY
Y@YUUY���ZYUUYUUUUUUUU���ZYUUY  Y�Y(*Y**Y*�Y�Y��Y�"Y�*YY�YYUUY���ZUUUUUUUU���ZYUUY  Y(
Y�*Y�*Y�*Y�*Y�
Y�Y� YYUUY���ZYUUYUUUUUUUU�Z�Z�
Y�*Y��Y��Y��Y��Y�*Y�
Y)
Y�
Y�YUUY���ZUUUU������ ���������0������� ��� ��� ��� ��� �������0���������������� �0��0�� ��3  �  ���������������������������������      ?   �   �  �  �?  ��  �� �� ��? �� ������?�������� ��0 ��� �� � � 0� ���  �  �  0�  ��   �   �   �   �   �   �   �   �  ��  ��  ��  �� ��� ��� ��� �����?����������������� 0�� �� ��� ?�0 � �� �  0      �   3         ���� �����0������� ��3 �� ��3 ��� ������0��������� �   �   �   ?   ?   ?   ?                              ���� ���  ��   �                                                ������? �?  ?                                                   �������������������������� �� �� ��  �?  �?  �  �  �  �     �   �   �   �  ��  0�  �  � ��� 0� � �� ��0 �� ������������?������ ��? �� �� ��  �?  �  �  �   ?               3   �       0  �  �� � ?�0 ��� �� �� �� 0����������������?� ��� ��� ��� ���  ��  ��  ��  ��   �   �   �   �                                �  �  �  � �� �� �� �� ������������������������������������������������������������������* ��* ��* ��* ��* ��* ��* ��* ��* ��* ��* ��* ��* ��* ��* ��*                     �( �

 �� ��  �*  �
  �  �   *   
      ����������������������������������������      �                                    W                                  <Tw                                  ��V�                                  ���?                                  @h��                                    ���  ������?                           ���=  0 <?0                           h��?  ��??�?                           ��=�  ��??3�?    <                       ��� ��???<                             �/ ��???�?                             �'  ��???�?    <                        �'  ��<?0                             h)  ������?                        ����������������������������������������                                        ��������        @UUUUUUU                <� � �        @      @����            ��������        @���3C����            ��������        @�333C����            <� � ��        @���� C����            ��������        @�33� @����            ��������        @��33� C����            ��� �        @UUUUUUU����            ��������                                ���������������������������������������� �   \  �  t  �   �  w5 �����������?_����s���s�_����?�� � < v��?����|W��P���P]��P��?��� ��? �� <� �  �  _  �   �?  �� �s� ��� ��� ��?0�� ���w�W���|U�? ��� �� �s� ���  �?�?  ��  p�  p�  �� �� ���?������������}���_�?�U> wW� V��   ��?_�����������������?����������? \�  �W   W  �  �7  �5     �?  ��  p�  ��0 ��< �� �� ��__�u������=_�����Ý < � @/��  _� �� �� ��_ �U=�_W������7? ?7�� _� �� w� _�  ��     ;��� �� �U���O_�}��w��w�����? ��� ���  �  �  _  � �   \  �  t  �   �  w5 �����������*
����#���#�

����*�� � < vÏ*����|W��P��P]ϠP��*��� ��? �� <� �  �  

  �   �*  �� �#� �� ��� ��*0�� ���w�W���|U�/ ��� �/� �#� ���  �* �  

  � � <� �� ��? ��� P��*P]ϠP��|W������vÏ*� < �� ��*

�����������������*����������? \�  �W   W  �  �7  �5     �*  ��   �  ��0 ��< �� �� ��_
�u������=
��ר�Ý < � @/��  
� �� �� ��_ �U=�_W������7? ?7�� 
� �� 2� 
�  ��     ;��� �� �U���O
�}��w��w�����? ��� ���  �  �  

  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �   �� �<�??���������                                      <   �   � P�  W? �� _�3                              �  p  p?  � @� ��  @�  t  ��         <   �   �  �   7   7   �     �   7   7   7   7   ?           �  p  p?  �  �  p  �3  �?  �  p  |7  �<  ?<  �                                      �   \    �  �W �<|0��                            �   \    �  �W  ��  �M  @ ��         �   \    �  p  p  \  �  �  p  p  p  p  �          �  p  �  p  �  �  �7  ��  ��  �  �=  <�  <�  �  ????333333333333 3333  333    3     33333 33333 3333  333    3     3333  3333  3333  333    3     333    333    333    333    3     3     3     3     3     3        �  (  "  ������?���l�� <) q q q qqq q q  q$q () q q q q q q qq q$q&i	&Y	$I IIY	i	() qqqqqqqq q$q i() qqqqqqiqq q$q6�() qqqqqqiiqq q$q() qqiq iq q iqiqq  q $q6�() qqiq iq q iqiqq  q $qi�() qqq q q qqq  q $q$i iiiii6�() q q q qqq q q  q $q  iiYEE55%%  $$�$� � �������%%5 5�() q q q qqqqq q$q iiYYI%%  �$�$�$� � ���������% %Ս() q q q qqq q q  q $q  iiYEE55%%  $$�$� � �������%%5 5$= =�() qqqqqqqq q$qii ==��� � �$�$�$� � ������������� ��() q q q q q q qq q$q iiYYIIYYii))) )$)9	I	Y	i	() qqqqqqqq q$q ))))))9	I	Y	i	iiYYI I 9"9$9() 999999 AAQQa a q q qqqqqq q$q() q q q qqq q q  q$q iiKL() qqqqqqqq q$qiiKL() qqqqqqqq q$q iiYYI5 5  5 $5  -$-$-�() qqqqqqqq q$qii      EE55%� �  � $� $��() qqqqqqqq q$q �        --() 1 1 1 1 1 )iiYYII9)		� � �$�  qqqqqqqq q$q ٌ() qqqqqqqq q$q � � � 
�� � �  � ь() qqqqqqqq q$q ]]MM==5 5 5 5 5  5 $5  -$-$()        ����� � �$�$ qqqqqqqq q$q& () qqqqqqqq q$q       �،() qqqqqqqq q$q iYY YY$Ii	() qqqqqqqq q$q IIIII)) )$)i	Y	9	I	Y	i	$!�() qqqqqqqq q$q ))i	Y	I	9	)	)	�() qqq q q qqq q$q iiYYII99))99IIY Y i$i  () qqq q q qqq q$qii     MM="="-""��� "� $� "�() qqqqqqqq q$q �  ��         "�() qqq q q qqq q$qi!11AAQQ ! 11QQAA1!	  	 $	  �() qqqqqqqq q$q 	  !!11QQAA11!!"�() qqq q q qqq q$qi  
  QQAA1!	  	 $	  �() qqq q q qqq q$q11!999 91 1 !QQAA1!	  	 $	 aaqq ii �() qqq q q qqq q$q  
  QQAA1!	  	 $	  iiYYYYY �() qqq q q qqq q$q ]]MM=  $$�() qqqqqqqq q$q%%%%$�() qqq q q qqq q$qYYI
I
99)iiYYI9))!  ! $!  � !� � � ���  �() qqq q q qqq q$q !  !!���� � � � � ��$� $�&��() qqqqqqqq q$q � ������55%%$�() qqqqqqqq q$qEEEEii5�() qqqqqqqq q$q111111!!�!�!�����������Ս() qqq q q qqq q$q!11AAQQ ! 11aaqqQQAA1!	  	 $	  �() qqq q q qqq q$q iiYYII99))99AA A$A() qqq q q qqq q$q A AA%%����QQUUUUUUU U$U%�%��() qqqqqqqq q$q U M�	�	����EEE=!! ! )$)$9�M() qqqqqqqq q$q 9 Q Q Q Q II99)    %$% )J() qqqqqqqq q$qii i ]]MMEEEEE"E$E=="=$=i	Y	I	i	Y	I	 -�() qqqqqqqq q$qii i===55"5$5i	Y	I	i	Y	I	A	 -�() q q q qqq q q  q $q  iiYYII99))99IIY Y i$i�() qqqqqqqq q$qiii"i	KL() q q q qqq q q  q $q  iiYYii==--�������� �   --�L() q q q qqq q q  q $q  iiYYii==--���������M() q q q qqq q q  q $q  iiYYii==--���������M() q q q qqq q q  q $q  iiYEE55%%  $$�$� � �������%%5 5$= =�() qqqqqqqq q$qii ===-
-
�������
�������

--
�J() qqqqqqqq q$q 	  !!11QQAA11!!$�() qqqqqqqq q$q iiYYii55- - 5$5$= �() qqqqqqqq q$q =======5$  i
iQL() qqqqqqqq q$q      ]]MM==MMUUUU U"U--  �$� $�() qqqqqqqq q$q � � � 
� 9 9 9 9 11!!�  � $�  �() qqqqqqqq q$q � � �  ��	�M))99Q Q  Q $Q $Q() qqqqqqqq q$q
))	���
���� � 	
�LQ Q Q Q Q  Q�() qqqqqqqq q$qiKLiM M =$=$-$    $ !11999 91 1 !$��$�  � () qqqqqqqq q$q�  � 
����� � � ����� � $$$�$� � �ƍ() qqqqqqqq q$q  --==E E E E E ==- -   �����  � $�  � () qqqqqqqq q$q � � � � � ��� � �$�$ �() qqqqqqqq q$q  � $$�() qqqqqqqq q$q  ���5 5 %$%$]]UUU U$U M$M��() qqqqqqqq q$qAQQYYYYYI I 9() qqqqqqqq q$q iiQQQ$A() qqqqqqqq q$q AAAEEE1"1$1$!�i() qqqqqqqq q$q 1 )%�(                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���*      �?�?      ���  i�  ��� ����  L��  ��`����� ������� � �� ��� ��� �����  L��ˢ ���  ������� ��� � ��`���  �4�� �@�� ���" �(��!   �`		




2Px(( ( X(*(JLbd(-:-�� ��U� �	 
 �� � �`�U� � �� �	 
 �`�
    �
    �
    �
 
�  � �  � �  � � 
 � �  � �  � � � 
  �
    �
    �
    
                   
     PP            
   PUpp  P       �  
 P �ppPUp          
 p p pp�p         
 p ppqp p         
 p ��]pp         
 p p ��p         
 p pU p pU         
 pU�  pU�      �  
 �    �          
                   
                    �
    �
    �
    ��  �  � �  � �  � �   � �  � �  � �      �
    �
    �
     �
    �
    �
    � � �  � �  � �  �� 
  � �  � �  � �  
   �
    �
    �
  
                   
     PP          �  
 P   ppPU           
 p PUpp�P         
 p �ppp p         
 p p pqpp         
 p p�]�p         
 p ��p p          
 pUp  pUp       �  
 �pU  �pU        
   �    �        
                    
                  � 
�
    �
    �
    � � �  � �  � �  �    � �  � �  � �      �
    �
    �
     �
    �
    �
      � �  � �  � �  � �  � �  � �  � �� 
    �
    �
    �
  
 P                 
 p     PU          
 p   PP�P       �  
 p PUppp p          
 p �pppp         
 p p pp�p         
 pUppqp p         
 ���]pUp         
   p ��pU         
   pU   �      �  
   �              
                   
                    
 �
    �
    �
   � 
� �  � �  � �  � �  � �  � �  � � 
    �
    �
    �
     �
    �
    �
      � �  � �  � �    �  � �  � �  � � �
    �
    �
    �� 
                    
 P     PU          
 p PU  �P         
 p �  p p       �  
 p p PPpp          
 p ppp�p         
 p �ppp p         
 pUp pppUp         
 �pUpq�pU        
   ��]  �         
     �          �  
                  
                   
  �
    �
    �
    
 � �  � �  � � � 
�  � �  � �  � � �
    �
    �
    �
     �
    �
    �
     � �  � �  � �  � �  � �  � �  �  
�
    �
    �
    � 
         P        � 
   PU    p          
 P �  PUp         
 p p PP�p         
 p pppp p       �  
 p �pppp          
 p p pp�pU        
 p pUpqp �        
 pU��]pU          
 �  ��          
                   
                 �  
                   
   �
    �
    �
  
  � �  � �  � �  � �  � �  � �  ��  �
    �
    �
    � 
    �
    �
    �
  �  � �  � �  � � 
� �  � �  � �  � 
 �
    �
    �
   � 
                    
   PU    P         
   �PP  p         
 P p ppPUp       �  
 p ppp�p          
 p �ppp p         
 p p pqpp         
 p pU�]�pU        
 p ��p �        
 pU   pU           
 �    �        �  
                   
                   
    �
    �
    �
  �  � �  � �  � ��  � �  � �  � �  �   �
    �
    �
     ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WuU5 �_U pU�  �_� <�{5 ��k� W��� \WU� �WU? W�� �� ���? �_�      ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WuU5 �_U pU�  �_�  ܫ7  ��7  _��  W��  W��  ���  ��� �W�� ���      ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WUU5 �_U pU�  �_?   �?   ��   �_  �U  �U  ��  W�  �� �� ��� ���  ��� ���? ���? pw�� pU�� pW�� |W�� W��� WU�� WUU5 �_U pU�  �_?   �?   ��  �W <�U� <�U� ���� ���� ����  ���    �  � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \U]� �U�?  WU ��� \�7< W��� W��� �U�5 �U� W�� ��� �WW? ��       � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \U]� �U�?  WU ��� ��7  ܪ�  �W�  �_�  ?�  ?��  ?�?  _� ��       � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \UU� �U�?  WU  ��  �7   ��  ���  �U�  �U�  ���  ���  �W�  ��� ���  � ���? ��� ��� ��� ��U �_� �W�= W��� WWU� \UU� �U�?  WU  ��  �7   ��  ���0 �U�< �U�< ��?? ��?? ��?? ��      �?��?�����?�������?�?���ꬪ����:;쬯��Ϊ:��;��묮����:;�������?;�;�;��� ��:;��  ��: ;��;�;��� ��;��� ����:�;�;�����;������:;�;����:;� ���: ;�;�?�묯����:�������?;���:�ꬪ����:�꬯���:;��?�?�?�������?�� ���??��?������? ����?���쫳���:�� 찳Ϊ:;��쬳��?;� 찳��:;���쬳�� ;  찳�:?;�� ������? 쿳�: ��� ����;�� 쿳�:?����쬳� ; � 찳�:;;���쬳��;?� 찳��:;��쬳���:�� 찳Ϊ:;��?������? ����??��� \UW����<p �  7 � |�?WU���  �  �      �������������������\Wppppp|�W5��?<�?���<���?���<��<<���<��< � ��<��< ���<��<<�������?�?��?�������?��? ������?��� ����< �� �������� �������� ���� �? �������� ���?���� �?������<������?������<�����<<�< ��<��� <<�?���<��� �?����<������ ��<����<?������<����?<<��?���<���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ���  i驀� �
�4  �� ��� �� H� n� L� � K� $� r� �� �� � z��? �@ � �C  =� �� �� ��� �H  A����� ��  `� g� ��` �H ���W �����* ��������\�� ^������  ������ ������ 2������ �� � ꦀ���� ������Ч ݢ��� �� � �� $� ˬ �L:� i� ��  `� g�L© ��  `� g� =�:��`Hڢ
�; �0��0��0��0��0��0ʎ4 �h`H�Z� �  ��" ��! � �	 ���
 �
 � �	 �   ��
 �r� ���
 ��d� ��� �
 �
 � �	 � � �  ��!   �� � � � � � ��! ��    �� �D� ���� �� ���
 � ��! �	 � � �   ���	 i�	 �   �� � ��   ��� 8�� �   �� �T� ����z�h`xH�Z�  
����� ���� �! � �" � � ��� ��� � JJ��- �� i� � i � � � � �Ȁ�� � � �
�" � �LE�z�hX`H� �   ���� h`H�Z�/���� ���� ��z�h` ������ ͦ���� �� +� �� |� �` v�����e ͦ���^� �� +� �� |� ꦀK ڤ� �D� �� +��� V� ꦀ2 $�� �+� �� +��� V� ꦀ h�� � +��� V� ꦀ���H `�< � �>�< ��I�� �< m m i)�0im� mD mE ��  ^��� �ֈ� �� �`H��D � �E  |�h`H�; �� ��h`�Z�D ڮE ڮC ڭ@ �A  �� ި� �,mD � �,�(� ȱ,mE � ���  ����
Ș��̩��� ��C ��E ��D z�`H�Z�@ �A  ި� �,mD � ȱ,mE �  ^�����z�h`�Z�@ �A  ި� �,mD � ȱ,mE �  ����	������� z�`�Z�D ڮE ڮC ڭ@ �A  �� ި� �,mD � �+�'� ȱ,mE � ���  ����	���ͩ��� ��C ��E ��D z�`�Z�D ڮE ڭ@ �A  ި� �,mD �0:� ȱ,mE �  ����	���ܩ��� ��E ��D z�`�Z�D ڮE � ި� �,mD �� ȱ,mE �  ����	���ܩ��� ��E ��D z�`�Z�D ڮE � ި� �,mD � ȱ,mE ��  ����	���ܩ��� ��E ��D z�`�; �<  � ;� � ͦ������0��� � ;������ 4� ;������ �� ������� � ��© =�:�� ��`��� � � �B� � ��� �V� � ��
� �d� �;  ^�`��� �� �V� � ��� �d� �<  ^�`� �� �� �� �� �� �� �� �� �� �; �< �b�B `�5 �6 �7 �8 �9 �: �= �> �? �@ �C �H �# � � �K �� ��`H�  � �4 ��h`ڭ  � �4 ���`H ͦ���� �h`H� h`ڮ; ���� �`�Z� � �� ���z�`��� �� �D� �;  ^�`��� �� �� �7 )�  {��6  ^��5  ^�`��� �� �%� �� )�  {���  ^���  ^�`��� �� �_� �> )�  {��=  ^�`H ͦm? mD mE m5 m; m= )�0� �? h`H�Z�C H� �C �? 
����i� 轹�i�  짭? �A  ��h�C z�h`H�Z� H� H� � �
i� �


i� �a�  {���������h� h� z�h`H�Z�B H�F � �G � �a�B �@ �A  ��h�B z�h`H�Z +�����D �����D �����E  |�z�h`H�Z�D �E  E�� �F � �G �@ �A  ��z�h`H�Z� � � �  ި� �,
m � ȱ,


m � �B �  {�����z�h`H�Z�A 
�����* 轗��+ �C 
��*�, ȱ*�- z�h`�7 ͍ 0��6 ͌ 0��5 ͋ 0 '�`�5 �� �6 �� �7 �� `�W�N0��V�M0��U�L0 Z�`�U�L�V�M�W�N`H�Z��)	��& � �3��� ��0���h�2 �N�3 � � ���. ȹ��/ � � ���� �. ȹ� �/ �� F�� =�:� ���0�� �2 �2 �C�2 Z� �c��� ��0��z�:Ъ�ߍ& z�h`HZڭ2 i�0 �3 �1 � � �m2 �h�.�0������. i�. �/ i �/ �0 i0�0 �1 i �1 ����zh`HZڭ2 �0 �3 �1 � � �m2 �h�.�0������. i�. �/ i �/ �0 i0�0 �1 i �1 ����zh`HZک�� �� �2 i�0 �3 8�@�1 �1 � �	�0 0�00�0 8�0�0 �1 � �1 � �ڭ0 i� �$�; )�JJJJ�  {��; )�  {��zh`H�Z�9 �0f� ��  `� g� �� �� � m��� � ��� ��8 )�8 �9 �: �C �� �K �K ʈ� ��K �L �M �N  � � $� K� r�� n�z�h`H�Z�I �J � � �
��K ���ȹK )��	H� =� H�h���ܭI � ��J � � �� r�z�h`H�Z� �� +����� z������Z�
��K � �K � �
�� �k ȭ �k z�� �ψZ�
�� �k șk z� �� �k �K �� �� � ��z�h`H�Z� ڢ� z�����b�  m�� �� =�� z�����a�  m�� �� =������z�h`H�Z���  E� {�����z�h`�C ��� �C `�C ��:�C `H�Z�@ 

mC �����m5 �5 �6 i �6 �7 i )�7 �z�h`H�Z�@ 

mC �����m8 �8 �9 i �9 �: i )�: �z�h`H��; i�; �h`H�; � ��8��; �h`H��< �0��< ��< i�< �h`H�< � ��8��< �(h`H��= i�= �> i �> �h`H�Z� �0�� � JJJ� � 
m � �� � �	� 
�� ��� � �K  �K z�h`H�Z� �0�� � JJJ� � 
m � �� � �	� 
�� ��� I�� �K - �K z�h`�Z� �0�� � JJJ� � 
m � �� � �	� 
�� ��� � �K - � ����� z�`H�Z� �0�� � JJJ� �� � �	� 
�� ��� � �I  �I z�h`�Z��0�� �JJJ� �� � �	� 
�� ��� � �I - � ����� z�`H�Z� ��  `� g� �� ��J� �c� �  m�ڊ�I�:� m�� =������ E���� �  ��( =�:��z�h`H�Z� � � �  �����B � ��a�  E� {���������z�h`H�Z�
i� �


i� z�h`H�Z `� g��)��&  ��� �� ��� � �� ����� �� $��ߍ&  W� ��z�h`H�Z� � H� H�
� �� �  ^�h� h� z�h`H�Z� � H� H�
� �2� �  ^�h� h� z�h`H�Z� � H� H�
� �F� �  ^�h� h� z�h`��� �� �� �  �驪� �� �
� � ���� � @��0��� ��C��0��`H�Z�)�JJJJ�  {��)�  {�z�h`xH�Z� �a��$��b��%��c��&��d��'��7� �`� �� � ��� ��� � �- �� Ȳ- �� �� ��� � z�hX`� � � � � � � � � � � �( �) �* ` ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              ��>�����i�"���>�����i�"���>�����i�"���>�����i�"�ۍۍˎˎS�S�ˎˎۍۍˎˎS�S�ˎˎۍۍˎˎS�S�ˎˎS�C�C�S�3�#�#�3�S�C�C�S�3�#�#�3�S�C�C�S�3�#�#�3�F8-$$      		      ; <         �      �    �   �  �  �   �      ��  � ��   �  �   � �   �   �  �  �� �   �      � �   �    �      �   �     ǳϳ׳߳����������'�/�'�/�7�?�7�?�G�O�G�O�W�W�W�W�_�g�o�w������
dnx                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       ���ة��  ��� � � � � � � �ߍ& ��"  갢 t ���� �� �� � ����� ��� i�XL �H�Z� � �P0� � � � �� �0� ��0� �� �� ��� � �� ��(z�h@H�$ �% hX@                                                                                                                                                                                                                                                                                                                                                               ���  :�� �� =�:��  � `� H�� � n� �� =� �� �� =� i�� ���  �� �� i� H� n� �� �� �� =� i�7��� ���Т  v� �� ��`�� �� � ��� �(� � ��� ��� �� 3� �� Z�` �� �� �� ��`�� �(� `�� �� `��� �  v�� L� �ʜ  i�ߍ&  :�`�6�L�M�N�O�P�Q�R�S�T`�U�V�W�# `� �
� �H� �I�
 � �	 � �
 ��� ��� � �- �	 ��	 �	 �(��	 � i(� � i � � � �J�� �Ŝ �H� �
 ��KФ`�H� �I� �J�! �K�" � � �
�  ��`� � �
� �W �V  �U  �`� � �� �N �M  �L  �`�d� �� � ��; ���d�
������ȩ� �W �V  �U  ���Ui
�U�Vi �V�Wi �W��� � =���`H�Z� � � � � � �	 � � ��� ��� �	 ��� �- ��	 �	 �(�� i(� � i � �	 � � �! �� ��� � � � ��" М� � � � z�h`H�Z� � � � � � �	 � � ��� ��� �	 �- �� �M��	 �	 �(�� i(� � i � �	 � � �! �� ��� � � � ��" М� � � � z�h`H�Z� � � � � � �	 � � ��� ��� �	 �- � ��	 �	 �(�� i(� � i � �	 � � �! �� �Ŝ � � � ��" Ф� � � � z�h`� �	 � � ��� ��� � �	 �I��� � �! ��	 �� �	 � ��" ��`�F� �� � ��R� �� � ��^� �� � ��6� �� � ���; �
� �F� �c�  ��  ��M������H�� �� �� =�
� �a�  ��; ���
� 8� �� �; ����; �
� �^� ��L;ǩ �� �� =�
� �a�  ��; ���
� � i� �; L�Ʃ�; �
� �F� L�Ʃ ��
� �a�  ��� � � �
� ��! �
�" �
� � �  	� =� =� =�� � � ��`�K� �� �
 ��_� �� � �� �7�
� �K� �c�  ��  ��������<�� �� =�
� �a�  ��7���
� �K� �7����7�
� �_� �� �� =�
� �a�  ��7���
� �_� ��7���7�
� �K� L�ǩ �� ��`H�Z `� g� �� ��  ��� �H�F� �I�
�J��K ,é ���)��&  ��  	��� =� �� v� W� ����� �� �  �� ��z�h`H�Z�  	���  �� �� KȀ i� � ��  `� g���Gz�h`� �G�:�5��F�4�(�E� ���� ��E�E�E���2� �D oҜ� ���	�8�9�&�'�)�*�+�-�,�A�B�C�� ` i� �� �� �� 0� �� �� �ȩ ��  ��`�(�� �� �Щ �"�#� ��i�� ����  ϭ�� =� =� �  ���٢�P� �  ��� � �<�0 5������� �� ��8� �� � ��<�0 5����� �� ��` ��i��(�����" � Q� �˭�(� =� =� ����� =�:��`�� �(� � ��` �� �� ��` � x� �� �� �� �í6��� ��` � _ɩ  n�
�����$ ȹ���% ��$�
�	�$����F�  �� k� kӭG����ߍ& L­:��a �� IЭ9��e ]� έ8��	 ���L�� � i� n�F� �� � �� �� ĩd�0 5����� i�  y� �� ��L�ʩ� �<� �	 ���� �<� � ��x�0 5����� i� n� �� �<� �  ��d�0 5����� i�`�
� �(� �
 ��` �Ω��0�  �� 5����� i�`H�Z�
����( ȹ�i@�) ��(�D �(�t�iȱ(�E )�ɀ��%�E mpR� ��� �H�D��% aͭ$��5 Z�ȱ(� )��@�ɀ�� )� ��)��� �3)�  �̀���L��z�h`H�Z�,mD 8�� �E m� z�h`H�Z�

����( ȹ�i@�) ��(�(���Ȁ���(� �)�~)�ɀ��@�#�'� �g� )� ��&��V� �3)� ��(�E )�ɀ��%�E mp4� ��� �*�&��% aͭ$����(�D i�0
 )� �̀���L��z�h`H�Z��D 08�D � �8� � ��D 8�i� �E m� z�h`H�Z�E I�i�E 8��� �$���$z�h`H�Z��! ��" � 
����� ȹ��i@�  �� g�z�h`H�Z�%���q� F��8� �" �;��E 0�8�E � �'� �E 8�� 

m � � i � �8� �" z�h`H�Z��)�8�&�(�&�)�'�)�����$�
�	�	�$��d�,��8�%� �!�(�&�	�	�$����$�
�(�z�h`H�Z������; ��
�; �����; �z�h`�
� �P� � ��� �P� �;  �
� �d� � ��� �d� � �`H�Z��" �(�! ��� �� � �,�� ȹ,�i@�  g�z�h`H�Z�"��+� ��+�"i���+�"
����� ȹ��i@� �� �� ��! ��"  g�z�h`H�Z�"
����� ȹ��i@� �� �� ��! ��"  ��z�h`�Z�"� ���� �(�� ȹ(�i@� �� � � �i
� ��! ��"  g�z�`H�Z��1�0�F� �; �����i� ��� �	�i� 
m ��<��=ȹ<��<ȹ<��;z�h`�0� �� ��1�0��`� � �d�F� �;� ��;�%�<� �
�<�	�;��=� ��=��<�	�; 0р��9�C�	��C��C�B���B��B�A ��`�� ��  ��`�A  �d�  ��B �C �`�<� �� � ��P� �� �=  �d�  ��< �; �}� �
� � ��d�0 5����� i�`H�Z�� ��� �=  �� �< �� �; �z�h`H�Z "�)�	�1 H�)�	�% n�)�	� ��U� ��U��Lkҩ ��3)�ɀ�
��'�)���&�3)����8��[��v�
�wLk� oҭ2i�2��UiP�U�Vi �V�Wi �W؀l��Vi�V�Wi �Wح<���<�M�=�<�E��Vi�V�Wi �WحF�0+�F�&�F�!��UiP�U�Vi�V�Wi �W��4 ��z�h`H�Z�2�	���	����
�������D ���� ���z�h`H�Z�2�� �  ���D��� z�h`H�Z��! ��" � �.�� ȹ.�i@� ��� �D�  ��z�h`H�Z�1�0����������
������  %�z�h`� 
��.�� ȹ.�i@� �� ��� ��! ��"  ��`H�Z� � ��  %ө�� z�h`H�Z�#� � ��L���� �Ԁ$�� jր �� ـ�� ؀��
 ?ڀ� ��z�z` ���2`H�Z R� IЭ9���L�ԭ6���b �ȭ  	�����  	����խ2� �� �� ��L�ԭ  	�����2� �	 �� ��L�ԭ  	���� ��L�� 5���Ж� �"� 5����� *��� ��� �׀#����&�6����"�� *�L�� �L�ԩ�"��#�C ���& O�%�0�-��#�  	�����-����-��1�1�1�1��#�	�F�1 a�z�h`H�Z R� IЭ9���L�խ6���_ �ȭ  	�����  	����խ2� �� r� r� �� ��L�խ  	�����2� �	 �� ��L�խ  	���� ��L�� 5���А� �" *��� ��� �׀#����,�6����"�� *�L�� �L�խF�1��"��#�+ ���� ���F�1� �#��F�1��#�-z�h`H�Z��"� *���e���R ������ �\ �� �H �� �� k� ]ѭ  	���� 5������� а�  	���� *��8�"�3��#��"�' ߀"��#�-���"� �� �� ����#z�h`H�Z R� IЭ9���Lj׭6���a�  	����$�  	�����2� � �ө
�/ $�Lj� w�Lj� IЭ9���Lj׭  	�����2� � �ө
�/ $�Lj� 5����� ���� �ש �� ���#��"Lj� ����: *���H�6���  	����� ���#�-�,� ���#���-���#� ���" �� �� �׭F�1 a�z�h`��i�$ O�%�� �<��1 �� �� �׀1 �� �� �� k� �� ���"�#���# �ל-`��(0�8���	�i�`�� ��i��	�8��`H�Z�6����  	���� ��  	���� �� ����& O���"���' ��� �� �׀)L��La�L'� �� ��5 �����'L'�L�حF�1�"� �����"��#Ld�LM� *������έF�1�"� ������ �"�#Ld�LR� ������L\�L�� *��������1�1�1�1�"� �����7� �"��#�=�F�1�"� ��� �� �ש�"��#� 9� K� �� h� �� a� 5�����z�h`H�1� ��1h`H�Z IЭ9���L8ڭ6����  	�����2� �� rـ�  	�����F�1���1 *�����#��"L1� ����� O�%� �.�� �"� � �"�#�+�1�1�1�1��#�"� �׀�F�1��#���- 5����� a�z�h`H�Z�,��6�  	�����  	������1��2� �� �ө�, r� rـ�F�1�"��3��]��������
��L=�L��L��L��Lk�L � �� ��L]� ���� O�%� �� ��L=� ����" �� ��L=� ����! *��� �� �� �׀W �� ��L=ܩ�" ��L=� ���� ��� �# �� �� ��L=ܩ�" �� ��L=� K�L=ܩ�#�- ��L=� ������ �� �� ��L=ܩ�" ��L=� ��� ��� � �� �� ��L=� ����"L=�L]� O��� ��� ��� �׀Q��" ���D O�%� �
��#�-�0 *��� �׀!� �� �� �� x� �� =��� ���# a� 5�����z�h`H�Z�6���	�  ��t�3 �ȭ,��)�  	���� �� �� k� =�-��# �׀C��� IЭ9��3�6���
 �ȭG���" �� �� �� k� =���М,��#�U�-�F�1z�h`H�Z� �� r� r� �ҩ
�/ �ȭG��� IЭ9���Lޭ  	������"� 5����М"� 5����� *���~���	 �� $�L� �� ����#��#���-�,�#��%�1�1 �ҩ�#��#� � r� r� �ҩ �# έ8��L� ��� k� ]� ���/��ML�ܭ"��/��*� ��G���K ����>�/��*��#���-�- �� � �� *�� *�����#��"� ��*�F�1z�h`H�Z��* �� r� �ҩ�"�6����  ���L�� ����L�� ����- ����7� ���/�� ���� ���� �ހ>� �� �ש�#� ��*��#��" �� �ש �� O�%� �LZ� ��*�F�1z�h` �� *��� O�%� ���#���-� ����#�� ���#�-`H�Z�F�1�  	����J��"� ��G���[��G���R IЭ9��H�i� έ8��5� �� k��� � S�ɩ�"� ����-��#��"�# �� k�z�h`�5�5��%�5�4���:�4�� �  ���Ei�E��� `�4��E�E�E���  ��`ک�� �E� ��.�� ȹ.�i@� ��! �
�"  ���` x� �� �� �� ��`H�Z�  �� �� R� �� � �� 9�LG� �� ����" k� =� =� =� �� �� ����" kʭ8�����" � =� g� � IЭ9���LG���� � �ȭG���� =� g� ��� �ͩ ���" � =� =� g� ��" � =� =� =� g� ��"� IЭ9��5� ��� � �ȭG���  =� =� =� g� ��� �͜" � =� =�z�h`H�Z�  �� �� R� �� ����" � ϭ8�����" � =� g� � IЭ9���L5���� � �ȭG���� =� g� ��� �ͩ ���" � =� =� g� ��" � =� =� =� g� ��"�� �� IЭ9��0� � �ȭG���  =� =� =� g� ��� �͜" � =� =�z�h`H�Z�  �� R� ��i��" k� �ȭG���^� �� � IЭ9��L O�%� � ��1���i� �� =� =� �� �� k�LV��� *��#����"�#�F�1z�h`H�Z�  �� R� �� �� ����" k� �ȭG���� �� IЭ9��L^� O�%� � ��F��: *���" ���i�& �� =� =� �� �� k�L��8�� 9� K�#��#�F�1z�h`H�Z O�%� ������ ��-��#�) ��$�6����" �׭-����U� �� ��z�h`H�Z�  �� R� �� ����" k� �ȭG���f � IЭ9��Y��i�B �� =� �� k� O�%��,�������%��L����L5���L5� K�#� 9� ��F�1z�h`H�ڜ% �����%����%����%����%����%����%����%����%����%����%����%����%����%����%����%����%z�h`H�Z�"� ��"���"z�h`H�Z�"���"��"z�h` |� 1�`H�Z�����)�����)����� )�����!)����z�h`H�i
� �i�  ��h`H�Z� ��� ��� � ���� � ��� ��� � ��� � ��� ��� � �� � � ��� ��� � ��!z�h`HZ�i���� ��� � B�zh`H�Z�i���� ��� �i B�z�h`H�Z��������)�����	� ����)�����	� ����)0�0����	� ����)�������	� ���z�h`H�Z�i���� ��� ���ȱ�ȱ� ȱ�!�����������������)�����)�����)0�0����)�������)�����)�����)0�0����)������� )����� )����� )0�0���� )�������!)�����!)�����!)0�0����!)������z�h` 
� 1�`H�i� �i�  ��h`H�Z�8����� ��� �i���z�h`H�Z�i���� ��� �i���z�h`HZ�i���� ��� �i���zh`HZ����� ��� �i B�zh` �� 1�`Hڭ8�� �ʎ  ���h` �� 1�`H�� �i�  ��h`H�Z��6���
 �ȭG���9 IЭ9��/ �� �� έ8��� k� ]ѭ*� � �� 5������� жz�h`H�Z�P���� ���� ��z�h`H�Z� ���� ���� ��z�h`H�Z� �@� � � � ����� ���z�h`H�Z�� �@� � � � ���(������� � i0� � i � ��z�h`H�  ����h`H�  	���h`H�Z
����� ���� � ��$��a��b��c��d�8�7�  ��Ȁ�z�h`H�Z)�  ��z�h`H�Z�)�JJJJ�  ��)�  ��z�h`xH�Z� �a��$��b��%��c��&��d��'��b��(��7� �`�i@� �� � ��� ��� � �� � - �� i� � i � Ȳ� � - �� i� � i � �� Ъ� � z�hX`xH�Z� �a��$��b��%��c��&��d��'��b��(��7� �`� �� � ��� ��� � �- �� i� � i � Ȳ- �� i� � i � �� к� � z�hX`H�




� ��) �& �h`� v����( ����) � �& �@�' � � �(�&��(���& i0�& �' i �' �( i(�( �) i �) ���Ωߍ& ` 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p�����������������������������������������H�� �� ���� h`H�Z�� ���F�� 
����� ���� �� 

����'�* ȱ�



�� �� ȱ��� �) ȱ�� �( �� � ��z�h`�� �* `����'�0�9�>�C�kw � % 10 ��
 11      � �� ��  `� g� � � � � � � � �� �� �� �� �* �� �� �ߍ& `H�Z�� ���Q�� ���.�� � `�� �� � �  W�� � g�� �� � �  ���� �� �� � ��� �� �� � ��� ���.�� � `� g�� �� � � � �  ��� �� �� � ��z�h`�� �̍� ȱ̍� ȱ̍� ȱ̍� ȱ̍� )
��|��� �|��� Ȍ� �� �� �� � �'�� �ō� ȱō� � ��� � ��� ��Ȍ� �� ��`�� ��� ȱ�� ȱ�� ȱ�� ȱ�� )
��|��� �|��� Ȍ� �� �� �� � �#� ��  `� g�� �� � � �� �� � � `�� �ٍ� ȱٍ� ȱٍ� ȱٍ� ȱٍ� )
��|��� �|��� Ȍ� �� �� �� � �'�� �Ǎ� ȱǍ� � ��� � ��� ��Ȍ� �� ��`H�Z�� )?	@�� �� 4��-� �� �� �Ӫ�� )@��J��� �� Ȍ� ������� �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� �ભ� )@��J��� �� Ȍ� ������� �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ��� )@��J��� �� Ȍ� ������� �� �� �� � � �� �� z�h`� �� `� �� `H�Z

��D��� ȹD��� ȹD��� ȹD��� � �ō� �Ǎ� ȱō� �Ǎ� �� �� ��� ��  � �� W� ����� z�h`�ZH
��h��� ȹh��� �� ���  �� ���� hz�` �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��    �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��    �� �� �� �� �� �� �� �� �� ��   ��:�\�������\�:���\���\���\�\�}�    �� � �� � �� � �� �� �� �� �� �� �� �� � q� �� �� �� �� �� �� �� ��T�.�� �� � ?� ?� �    �� � �� � �� � �� �� �� �� �� �� q� � �� �� �� �� �� �� �� �� �� �� �� �� �� �� �    ���.����� �.�T�}����� ���}���������:��� 0�    ���.����� �.�T�}����� ���}���}��.�}�T�}� �    ��.� �.� �� ��.� � �� �
� �
� �
�T� �}�T�.�� �T�.� �
�.
� �
� �
� �
� �
� �
� �
� �
� ��    � �� �� _� T� �� � �
� �
� �
� ��   ��\�\�\�\�\�\�����\�\�\�\�\����
��
��
���������\�\�\�\�����\�\�\�\�\�   \���\��
�\
��
��
��
��
��
��
��
�\�\�\�\���\�\�\�\�\�\�}�T�\� ����
�\
��
���    ��    K�    �� �� � �� � _� K� ?� /�    �� �� �� �� �� �� �� � w� q� j� d� _� d� j� q� w� � �� �� �� �� �� �� ��    �� �� �� �� �    �� /2�   
	�

		�
�	
	 �				�

		���T�  ��6�  P�X�\�b�8�>�����  O�  ��E�  ��E�  ���������������f�  ���������������� �� �� ��    _� T� K� ?� ?� � ?� K� T� _� _� T� K� K� T� _� T � � _� T� K� ?� ?� � ?� K� T� _� _� T� K� K� T� T� _� � � _� @�    _� 2� 8� ?� G� K� T� _� � � _�   
	�

		�GAMEaaOVER$PAUSE$SELECTaaLEVEL$BEGINNER$aNOVICE$aEXPERT$TIMEaaaOVER$BEGIN$YOURaMOTORaDAMAGE$CONTINUE$TIMEaLIMITd$GOODaaLUCK$YOURaTIMEaa$SCOREd$END$ITaISaAaNEW$RECORD$PLEASEaSIGN$YOURaNAME$LEVEL$HEIGHT$GaTaC$SCORES$HIaSCORE$PUSHaaSTART$PUSHaSLKEYaRESELECT$RACE$REACHaGOAL$�����������	�	���-�6�B�M�Y�`�d�p�w���������������������c2cgc�c�c�cd4did�die�erf�f$ghg�g�gh�hichJi�i�i%jZj�j�jPk�klml�lm�m�m3nnn�nAo+p�p�prqr�rTq sOs�s"t�tu�u�o�o�q�u$vhv�v5w�w�wUx�x=y�y�y6zwz�z�z�B�B0CpC�C�C0DpD�D�D0EpE�E�E0FpF�F�F0GpG�G�G0HpHqH�H�H1IqI�I�I1JqJ�J�J1K�OPQP�P�PQQQ�Q�QRQR�R�RSQS�S `@`�`�` a@a�a�a b�B�BqK@bEbhb�b�b�b�b                       ���������@�i����� 	 1	451	45d 23 
23 
d d $% 3"6
$% 3"6
 d ! &'(78 " ! &'(78 " d ) *+/9) *+/9 d ,-.:;<=>?00,-.:;<=>?00d GHI.@ABCDEF2GHI.@ABCDEF2d������]�������	�a� � �                                                                                                                                                                                                                                                                   R� ���