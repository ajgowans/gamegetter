                            !! !" ! !" !!!! !!" !!!" ! "   !" ! !"!!"  !!"!!!" !!" !!"  !!" ! "  !" !!!" !!"  !!" ! !" !!"  )++++++++, )++++++++,  )++, )+*+, )+++, )*+,  )++, )+++, )+*+, )++,  )+*,)+++, )+++, )++,  )++, )+*+,)++*, )++,  )++, )+++, )+++,)++, )++, )+++, )+*+, )++,  )+*, )+*+, )+++, )*+, #$$%#$$$%#$$$%#$$%                               #$$%#$$$%#$$$%#$$% !!!!" !!!!!!" !!!!"  !!!"  !!! !" !!!!"  !! !" !"!!" !! !"  !!!!" !!!!!!" !!!!"  "!"!!!!! "!!!!" !!!!" !!"!"  !!!" !! !" !!!!!!" !!!"   !!!"  !!! !" ! !!" -..../-....../-..../ )++++, )++++++, )+++++ )+*++, )*+++++, )++++,  )++++,)+,)++, )+*++,)++++, )+, )*+, )++++,  )++++, )+, )++, )++++,  )++++, )+, )++, )*+*+++++++*+, )*, )++, )++++,  )+*++, )+*++*+, )*+++, -..../-....../-..../                      )++*+++, !!!! )+*,!!!!! "      )++,  !!"!!!!!!!!!" !!!!!!!! +++++++++, )++++++++   !!" )+*+++*, ! " )++,)++++++,)++, )++*+*+++, )++++++++,  )++++++++,)++*+*+++, )++++**++, )+**+++++, +++, )++++, )++++, )+++++, )++++, )++++, )++++++, )+++++++++++,)++++++, )+++++++++++, )+++ )+,)++*+, )++*++*++, )*+*+*+++, )+++*+*++, )++++++++,)++++++++, b�b���������r�r���88Z00���  688Z\H�H�0x  688Z\`xz`�0x�H�x0�   688ZZ\`xzH��H`�0x�xH�    <<VT\rx�0�H��00�x��H   <>BTVttx�0��0��`���H�    &$6>PZ`nlH���`Hب�0�   68>NNbhll��0�H�0ؐ�0�   ***06Z```flrr��H�H�H0H��0��,,BBB```0H�`xHx  B,NNNr�`�0x`�H�		***8B`x���H�`x��x  ,8TTbbxx�H�0HH�x		BBBBBHTTTT�����H`x�� 0���xH��H�x� 	 	 
bb � � D D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �� �����?����?����?����              W�W=\UU�WUUP�WTU�W�\U=              W�W�\UU�WUT�WUU�W�\U�              W�W�\U�WUU�WAUU�_A?\U�              W���_U�WUAU�WPUU�_P?WU�              _���WUA�WUPU�TUU�?T�WU�              \U�A�WUP�WTU�UUU�3U�W�?              \U�P�W�?T��U���_U���U�U�?              \U�T�U�?U��OU���_U���U�U�?              \U?U�U�U��_U���_U���WuU�              |UU�U�U�\U�  \U�  WUU�              pU\UUU�U�\U�  \U�  WUU�              pTUUU�U�\U�  \U�  _UU�              pUUUU�U�\U�  \U�  \UU�              pAUUUU�sU�\U�  \U�  |U�               �PUUU�sU�\U�  \U�  pU�               �TUuU�sU�\U�  \U�  �UA�               �UUuUA�pU�\�  \�  �UP?               �UU�UP�p�\�  \�  ��?               �UU�T�p�\A�  \A�  ��?               �WU��?pA�\P�  \P�  pA�                WU�C�?pP�T�  T�  pP�                W��S�?0T�U�  U�  <T�                W��_�0U�LU�  LU�  U�                �����������  ���  ���                �����������  ���  ���                ��?�� �����  ���  ���                 ��?�� �� ��   ��   ��                  � �  �� ��                                                                                                                                                                                                                                                                                                                           ��   ���? ����?                         T �UU� WUT�                        �U� �AUU�WUU�                       \AUU�PUU�WUAU�                       WPUU=�TUU�WUPU�                      �TUU��UUU�WTU�                     �UUU��U�U�WUU�              ;   �   �AU�W�pU�W��OU��              �   �  pP��_�pU���_U��              ���?�  0T����pU���_U��              ����  0U���pUUA� \U�                ����  pU���pUUP� \U�                ��jU�  pU�  pUT� \U�                cUUU�  pU�  |UU�? \U�               �ZUUU�  pU�  \UAUU? \U�               �Z�U}U  pU��\UPUU? \U�               �VUUUU:  pU�\=\�UU? \U�             � �VUUUU: <�UU�W�\�W? \�             ��VUUUU:�;�UUAU�\A�W? \�             �>�U�WU�:�UUPU�\P�WA? \A�             ��U��Ε���WTU�T�WP? \P�             ���V�å�� _UU�U�T� T�             ���j�W	�� AU��CU�U� U�             ��
�ZU� �� �SU��SU�OU� LU�             �� �}*  �� ����������� ���             ��  � P�� ����?������ ���             ��  �@ �: ���������� ���             ��U?  �  ��? ��?���  ��             �� ��U�                              �
     �                               �*P�@ �:                               �  �: �                              �_�
 p9�>                               �U�+ p�                               _UU��|�                             �zUU���WU�                            ��UUU��VUU=                            ��UU�UV�UUU�                         �? �WUW�jUUUU                        p�|��WUU��UU                        _U�W��pUUU��VU              ?�     ��UUU�W� \UUU��jU5             ��30     pW�_UUU��WUUU� ��?             0 0     pW}UUUU5pUUUU� ��            0(0<     ���WU��\UUUU9  \}5            0�0�     �UU5  WUUUU9 �W5            0�  <      ��U �UU��W���W5            �( ��        � |U���WpU_?            �� <           W� ����pU��             ?  �         ���?����7pW��             0  �         p}������7�W�=             � ��         �WU����> ���             � �           \UUU�z�� W]�              � <        \UUUU鮪 �]�              �����       \UUUU��� ��?              0 ? �       \UUUU��>  �                 ��       \UUUU��                   �         \UUUU�                   �?          pUUUU�    0                ��        pUUUU�    0                0�?   ���� �UUU�j    �              �  0�?   <�� _]��o                  �
 ��   ��� �_��l                  _��     ��*� �W�l �              �����    ���*� � l �:  0            pU���    �ꯪ��z� l ��  �            \U���    ������^�  l5 k�             \UU��   ����>W_9  �5 [�  <           WUUUU   � ��:�u:  �5�Z�  �           WUUUU   ��?�:|u  �տ��   �         �UUUUU     ?�����  �V�5     ?         �UUUUU     ������  �ZU5     �        �UUUUU     ��Ϫ��   �U     ��        �UUUUU     �����    ��      ��      ��UUUU�     ��?���   ?�?        ��?  ���WUUU�       �;��7 ���           ������? |U�W=       ���? \�E           ���  �����     ���� �h�                 ��? ��?     �:�� |���                 ���  ��     �:��?PW�?                 ��   ��      �������?                                                                                                                                                                                                                                            ��                                     0                                      <0                                     �0                                     0                                     0                                     �0                                     <0                                     0                                      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��������������������������������^UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�nUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������������������������������������������������������������������������������������������������������������������������������������e                            ���e                            ���e                            ���e      � ���?  �?�       ���e      �<���?  ����       ���e      �<��� ����       ���e      �<��� ����       ���e      �<���  ����       ���e      �����  ����       ���e      �����   ����       ���e      �����   ����       ���e                            ���e �������������������������
 ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e �������������������������
 ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���e                            ���%UUUUUUUUUUUUUUUUUUUUUUUUUUUU�����������������������������������QUUUUUUUUUUUUUUUUUUUUUUUUUUUU���TUUUUUUUUUUUUUUUUUUUUUUUUUUUU����������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 E    D   Q   @                                                                                                                               EDDDDDQ                                                                                                                                    �    �"" "� ����    "                                                                                                                          ������"""""�                                                                                                                                    �    �33 3� ����   03                                                                                                                          ������#""""�������                                                                                                                              �    �33 3� ����   03                                                                                                                          ������������������                                  p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    ��    |�    ��    ��    ��    |�    ��    ��    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p�    ��    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:    p5    �:    �:    �:                                                                                                    �?    �:    �:    �:    p5    �:    �:    �:\    �    �    �    \    �    �    �    \    �    �    �    \    �    �    �    �?    �=    �?    w7    �?    �=    �?    �?    \    �    �    �    \    �    �    �    \    �    �    �    \    �    �    �    _    �    �    �    \    �    �    �    \    �    �    �    \    �    �    �    \    �    �    �    \    �    �    �    \    �    �    �    \    �    �    �                                                                                                    �    �    �    �    \    �    �    �                                                                                                    ������WUUUUU     WUUUUU������W�    �>    �                                                                                                    ������UUUUUU      UUUUUU������  W�    �>    �                                                                                                  ������UUUUUU      UUUUUU������                                                                                                                  ������UUUUU�     �UUUUU�������    W�    �>    �                                                                                                ������WUUUUU��������j�����Z�f���V���������������                                                                                                ������UUUUUU��������j�����Z�f���V���������������                                                                                                ������UUUUUժ����ꪪj��ꪙZ�fꪪV��ꪪ����������                                                                                                ������CU@USUPUWU TU W�����W�    \0    �                                                                                                    ������@U@UPUPUTU TU �����  C�    \5    �                                                                                                  ������@U@UPUPUTU TU ������                                                                                                                  ������@U@U�PUPU�TU TU������   ��    0    �                                                                                                ����������������f���Z�f���Z�f�����f�������������                                                                                                ����������������f���Z�f���Z�f�����f�������������                                                                                                �����������ꪙ��fꪙZ�fꪙZ�fꪙ��fꪪ����������                                                                                                ������CUPUT   CUPUC�������    0    �                                                                                                    ������@UPU T   @UPU�����  ��    0    �                                                                                                  ������@UPU T   @UPU������                                                                                                                  ������@UPU� T  �@UPU�����U�   ���    0    �                                                                                                �������������������������������zUU��������������                                                                                                �������������������������������^UU��������������                                                                                                ����������������몮���ꪮ����^UU�몪������������ p�Wp]]pWu�w�  w7  \  \ �z�  �5  W5 �U� �V�  [9  �? ���� p�Wp]]pWu�w�  w7  \  \ �z�  �5  W5 �U� �V��[����    �?� p�_pU�5�uu5�wu5�UU5 Wu \� �  \ \60 \�0 pY pU ��  �? �< \��pUw�]]�]]pUU�U] W�  �   \0 �5� \�0 pU pU �_ �� ���W\wU\]]\]�\UUp]� �s5  � 0p5 �5 �5 �e �U  �  �  <���_5p�UpuupuupUU�uU ��   ; �5 \6 �5 �U �U ��; �� �  p  p  p  p  p  p�  p�  p�  p  p  p  p  p  p  �  ���pUUpUUpUUpUUpUUp]UpwUp]UpUUpUUpUUpUUpUUpUU����?  �:  0  �:  �:  ��  �� �: �: �� ��  �:  �:  0  �:  �?    �  p  p  p  p  p    w    p  p  p  p  p  p  �����UU�UU�UU�UU�UU�Uu�U��Uu�UU�UU�UU�UU�UU�UU���  �?  �:  0  �:  �:  �: ��: ��: ��: ��:  �:  �:  �:  0  �:  �? � 7p �_ WU �] �] �] \�  �� �?  _��UW�UW��_���     � 7p �_ WU �] �] �] \� ���
 �?  _��UU�UW��_p�x5��?    � 7p �_0WU��]����?���WWWը�U��U5�U�7 _�� �(� �*� �
�� 7p �_ WU��]��� ����?WW5��U��U��UU5�U�7 _�7�~��ré��ã     �� ������U��u��w7W�w7W���WU+*\U��WU��� 7(� 7�� ?�>  �� �� ����U��u� w7�w7\���WU**WU�\UU�WU��� ���jÍ�Ã�� �� ��� �U� �u�  w7 �w7 ���0 +*� �� p�� pU5 p�7 p}5 �]5 ��? � 7p �_ WU �] ��  ��WW�� �? �_ \U �_ \} \u ��                  00  ��  \�  ��  ��  \�  �� �?  \�  \�  \�  ��                  00  ��  \�  ��  ��  ^� ��  �?  \�  \�  �_ ?�                 �  �} pU pw pw �Y ��  � �U5 �U��u  �                  �  �} pU pw pw �Y ��  � �U5�U�p�� ��?                   �  �} pU p� p� �e ��
 p�  \U�_U p] ��                   �  �} pU p� p� �e ��
 p� 0\U�_U � �� �  �  �� ����:������뫪�ꫪ�ꫪ������0;�3�:������ �? ���? �  �� ����:��;��;�3��뫯�ꫪ����:�3�:������ �?                                      �? S���TT����EE�S�� �?  �  ,  �2  +8  �2  +8 ��2 \+�W�rw=|��W�� g5 [5 \9  � � ��  ��  � �W� pUU\UU\PU\@U\AUpUUpUU�U�  W5  \  �             �� |U� WUW�VWUUWUUWUUWUUWUU\UU\UUpU� ��?     ����  �  ����UU�UU W�  \5  �  �  �  �  �  �?  ��  �   �  S5  W5  �  S5  W5  �  S5  W5  �  S5  W5  �  �   �   �  �  � ���p}}\]u5\]u5p}}����UU�UU ��  |=  \5  \5  �         �  ��  |� �WUpUUpUU\UU\UU\UU\UU\UUp�U��  �?                             ����SUU�SVV�CUU�Lee�UU10TU0�  ��      ��  ���00000000����\UU��UU= _� �?  �  �  �  �=  �����pUU\  5�*4B�ԇAAҫ�«AA�AA҇҇҇AAҫAA�«�     �e  pY \  � �e pY  \V pY  �e  �  \  pY �e              Y @e  �5  P�  TY  e P�5  e TY P�  �5 @e  Y             ��?�?�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �<<<<�    ������    � �� �    ����    ������    �< � �    �0 �<<�    ���� � �     �<�<<�    �<<� �  ��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                    ��  ��  �*V�V�V�V�V���*      �?�?                      ���  ��� � �6� � �7� �ύ& ��" � t ���d���� � �������� �ƩP�4d/��0�Z���# XL �H�Z�4�P��4��4�/�0�0z�(h@H�Z�' )������ Z� 8楝�# �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                                                                       � �� �Ʃ
 ��:�� � 7� � �̩ �� �� !� W� � �ƍC�C���HL­C	��[�C	�����C	�����C	�ɿ�$�C����/ �� �� �ƭC	�����C	�����b� ���	��E �ɀ � -րx � � �˩��KX � !� W� K� PǭL���L�� x� � �D��� PǭL���L��L*� Fɥ1� ��HL�LH�O�P��Q`�L�M�N�R�S�T�I�J�K��^���& G� � 9� s� �� t� *�`�H�G��U�P��V�Y��W��d?d@�N�O�P�Q� �Ui�� ��8�+�:� �Vi�� ��8頍;� �ƭH
�����轆�	�)��� ��U��W������ �UȀ� �íH������AdB���A��B���A��B� ��`�H
��t��8�t��9`� �ƭH
�����轘�	�)��� ��_�����E�D� ��`� �ƭH
��������	�)��� ������������������ ��`�H
���������� ��e�����y�z�{�|�}�~�������������������������������������`� �ƮH�b��X�
�����轪�	�)��� �����X����� ��Ȁ��mX��i �� �����X����� ��Ȁ��mX��i �� �����X����� ��Ȁ�������������`� �ƮH�k��[�H
�����轼�	�)��� �����[����� ��Ȁ��m[��i �� �����[����� ��Ȁ��m[��i �� ����[����� �Ȁ��m[��i �� ��"��[����� �"Ȁ�� ��`� �ƭH
��������	�)��� ��R����� ��`H�Z���H
�������������i������I�i������i����H���z�h`H�Z




���)�& z�h`H�Zd�@�� � � ��������z�h`�Z�/���� ���� ��z�`H�  �4�
��h`ڭ  �4�P���`H ������ �h`H ������h`Hd4h`�8�6�9�7dd�(�,`dd�(�,���A�8�6�9�7`� �L�b�� ?ҭb��Z���� � � ��a !� Wͩ0 ��:� ���^�^� ����L��� �� �� ��L� �� G� � s� 9ĩ �� ��LȠ �"� �Q��[���b !� Wͩ�� ��P ��:� ���H�H�	��H �� G� � s� �� t� 9� !� Wͩ �� ��`�C	�����C	����*�P�b� ����_�6�`�7 �ӥ"� ���bLȭb� ����_�6�`�7 �ӥ"� ���bL�`H�Z����& �ȭ��6���7 �ӥ"� ��I͘��H��z�h`H�Z�>����l��hL7ɭ`͘�1���I�_͗�
���HL+ɥ/)��L+ɍHL+ɩ�HL+ɭ`�I��H���6���7�7 �Ӧ'�U��L��LBɥ?�B�L�ȥ/)��L��z�h` � � ��d1���<��
 ����Z�� ��1���<���Z���d!d"�� �#��$d%���&� ��"��E�"��F �ѩ ��:� �� �ƍC� ��:� ���C	���C	�����C	�������1�1)�1LQɥ1� ��H �`�b����a�����a�	����a`H�Z� �Ʃ��&� �'��=��>� �������� �ʤ�r� ��������� �������� �'��> ����������>��' �ʤ�D� ��LY� �� �ƥ���>��� �' )���� �ʥ���' )����� �ʥ�� ��L�ʩ��� �2 ��:� ��� ��z�h`xH�Z�'
��?��E�?�	�)��Fd%d!d"�=� �#�>�$��8��$��$ ��z�hX`H� �& �ʩ��&h`��� �� �Ʃ 
��C��E�C�	�)��Fd%ddd!d"�(� �#���$ �ѩ �Ʃ
�����	 �� ��������� �`� ��:� ��� �Ʃ
��C��E�C�	�)��Fd%���'�d!d"� � �#�P�$ �ѩ �Ʃ��>�� ����H� 6���H�� ����^� 6���R�� ����Q� 6�P� 6�O� 6���\�� ����N� 6�M� 6�L� 6�L������g�� ���
��g��  �� �������  	��� �` �Ʃ��F�� ��P ��:� ��` � � �Ʃ��F�� ��H�)�� ��a��JJJJ� U�)� U�0 ��:� ��`�O� �1�O�N� �'�P�8�8�8� ���Q�9�8�9ə�� #�`H�Z��%�N�)�� ��a�JJJJ� U�)� U� � U� U�z�h`d'd(�������8���'���6e����8���'���*�8��+�7����8���'mU�'������"�8��$�'�(�8e�6�9e�7L"Υ$�A��@ n� �� �ϭb��	 �� -� �� �έA�$�@��e$��7e$�7��$d"���*�!�+�,��+�#��,�#�ɟ�QɈ���8��$ ��d!�e#�8��,�&�'�i8��,��,e��8��#LKΩ�#LKΥ(mU�(�'L��`H�Z�� d%�'�U
�����E轏��F ��z�h`H�Z�_��`� $Э<����a
�����E����F��% ��z�h`H�Z� �e��j��t��� �<� $Э<����o
����E���F��% ������z�h`H�Z�������?�A�� �<� $Э<�����)
��7��E�7��F��% ��z�h`H�Z� ������ $Э<�����
�����E����F ����X��z�h`H�Z� �������"� �� �<� $Э<����
����E���F��% ������z�h`H�Z��� �+������ $Э<�����
��;��E�;��F��% ��z�h`H�Z�� �#��$��6��68���L�Ѕ!���8�!�#LwХ8�6�,�L��e�d!�,e8����#��7�*�78���L�Ѕ"�78�9��8�"�A��A�$L�Х8�7�A�L��m78�9�d"�Am78����$���<�� �<z�h`H�Z�� �#��$��6��68���L�х!���8�!�#L5ѥ8�6�,�L��e�d!�,e8����#��7�*�78���L�х"�78�9��8�"�A��A�$L�ѥ8�7�A�L��m78�9�d"�Am78����$���<�� �<z�h`H�Z�"� ��Ee �E�Fi �F���Ee!�E�Fi �F� �C�@�D�� ��Ci0�C�Di �D���Ce�C�Di �D� � ڱE%&�%� ���1C�
��C�QC�C��#�����$��Ci0�C�Di �D�Ee �E�Fi �F��z�h`H�Z�`�;�8�;ɐ���bLӭD��L�ҭb����L�Ҡ ��>� ����>�t�����.�j�`�&�e�_�	�_8�e�8�_����b��aL����Ltҥ?�A�Lӭ��_�
8�_��4��_8���'���`�
8�`����`8���
��b��az�h`� ��>� ����>�t���e���j���o���y�����H���M���7��78���d�8�7��Z�����6͗�K8���C����6�98�6��1��M���U��
������U U��d�K�����>�K���t���e���j���o���y�H���M�����L�`d'�6����8���'����!�7����8���'mU�'�����"`� �=� ���7�L�Խ�� ���L������9��L����.L�ԭ]���6ݪ�X8����P�;���6�F8�6��>�)�]���6ݪ�-8����%����6�8�6���J� � �����=�	��X�L>�`� �?� �"� ��7����6�����\���?���[��`�_�6�`�7 �ԭ?���&�\�"�S�N�P�O���P���Q� �"`���� �C�d� �<�K����Smd�S�Ti �T�d��dmdmS�S�Ti �T�d� �K�LmR�L�MmS�M�NmT�N�ImR�I�JmS�J�KmT�K�R�S�T�Q�N��$�P�M�
��O�L��L�O�M�P�N�Q�K��	�^�K�K�`�?�A���@i�@�?i �?�`�b�]��c�D��V��M�_�6�6�6�`�7 �Ӧ'�U����#�6 �Ӧ'�U��
��E 3؀��E�D���E�D ـ ��Lq���l�D��_��V�_�6�6�6�6�6�6�`�7 �Ӧ'�U����#�6 �Ӧ'�U��
��E �؀��E�D���E�D ـ ��Lq���6�`��
� �b�]�% r׭_�6�`�7�c�) 9�)�c�]�bLq�� �) �׭b���_�6�`�7�c�) 9�)�c�]�b`�`��B� �b�`�`�`�`�`8�9�P��9���9�9�9�9�a� ���a�� �a`�`�;�8�;ɏ�f��b�`�`�`�`�`8�9�P��9�;��9�9�9�9�a� ���a�� �a�_�6�`�7 �Ӧ'�U�������b`�_��^��b�b�]� �=�_�6�`�7�J 7ԭ=���5�_�_8�8���8���8�P�E���a����a���a�E`�_�:�8�:�"�_��b�b�]� �=�_�6�`�7�J 7ԭ=���6�_�_8�8���8�:��8�P�E���a����a���a�E`�]��+�E���`���`�` 3؀;�`���`�` �؀)�E���`���`�` �؀�`���`�` 3حE� �C�D�_�6�`�7 �Ӧ'�U��������U� �b��'�c��U !� Wͩ�b`�]��.�E���`���` 3؀D�`���`�`�`�` 3؀,�E���`���` �؀�`���`�`�`�` �حE� �Z�D�_�6�`�7 �Ӧ'�U�������&�U� �b�+�'�c��U !� Wͩ�b�c�U��c�U����U`� ��>� ����>�t���e���j���o���y���~�F���G���H���I���M �ۭ��t���e���j���o���y�F�~�G���H���I���M�����Lz�`�?�A�L�۩�>�����������������������F���G���H���I���M �ۭ��������������������F���G���H���I���M��`H�Z �ȭ��]��'�M���>����������ML�ۭH��L
���c�F��V��M���6�6�6���7 �Ӧ'�U����#�6 �Ӧ'�U��
��G �݀��G�F���G�F �ހ c�L
���l�F��_��V���6�6�6�6�6�6���7 �Ӧ'�U����#�6 �Ӧ'�U��
��G >ހ��G�F���G�F �ހ c�L
���6����
� ���]�% ݭ��6���7���) ��)���]��L
�� �) Vݭ������6���7���) ��)���]��z�h`����@� ��ΘΘΘΘ�>��������	���������� ������ ��`���;�8�;ɏ�f��������>��������	���������� ������ �����6���7 �Ӧ'�U����
�����M`����f������]���6���7��J 7ԭ=���@Η�>����G�������
���!�����G��������������G`���:�8�:�"�f������]���6���7��J 7ԭ=���@��>����G����������!�����G��������������G`�]��+�G������ΘΘ �݀;������ >ހ)�G������ΘΘ >ހ������ �ݭG� �H�F���I���H���6���7 �Ӧ'�U����	�� ����'����U������U`�]��1�G������Θ �݀G���������� �݀,�G������Θ >ހ�������� >ޭG� �j�F���I���H���6���7 �Ӧ'�U����	� � ���6�'����U�U������U����U�����������U`H�Z �ӭ]� �/�"��&�'�U��� �]��)�U��
������UL��"� ��'�U���������]�U�'�)z�h`H�Z �ӭ]� �/�"��&�'�U��� �]��)�U��
������UL�"� �/�'�U��!��������
������U�'�)��]z�h`��� �L�᭩��2�������_Φ���6���7 �Φ���6���7 Ӏ9���:�8�:�#����$����6���7 �����6���7 �`H�Z�_�6�`�7�b�]��B�X�Y�Z�Y�Z�]��J�6�6�6�6� ���7� �6ݪ��Y�68���B�	�B�Y�Z��X���6�6�6�6�O��L���6�6�6�6� ���7� ���6��Y��8�6�B�	�B�Y�Z��X���6�6�6�6�X�Z�L�� �� � �ƮZ��� ����n�����e��(�������������������� � �� �ƀ9�����0�����'��#�������������� ������ � ��z�h`H�Z������� �Y��L��]���L��ΚL��]��3ΗΗΗ !� W�ΗΗ�4)����H���H��M������?�]��3��� !� W����4)����H���H��M������ z�h`�Z�]��6��� ���������B���_�����B���_:��L������
������B���_�����B���_:��� `� ��>� ����>�t���e���j���o�����H���M u䭚�t���e���j���o�H���M�����L�`H�Z�Z��͘�v��͗�8��8����+���H�����M�>�������� �������6��8���+���H�����M�>�������� ��Η���z�h`H�Z
����2���3d%� �2�$��a��b��c��d�8�7� U�Ȁ�z�h`H�Zd%��)�JJJJ� U�)� U�z�h`xH�Z� �C�@�D�� ��Ci0�C�Di �D����a��$��b��%��c��&��d��'�� � ��ȹ �����i��i �ʀ���%� ��QC�C���C�ȥ%� ��QC�C���C��Ci0�C�Di �D�� ����z�hX`� �K�L�M �� �� � � � � � � � �* d�d�� ����d�`�L����t� ��m� �n�  3��t�t�o� A�M������ ��z� �{�  ��恥��|� ��K���J�L����X� ��Q� �R�  ��M����f� ��_� �`�  ���X�X�S� ���f�f�a� �祜��� �� Z�`�N�O�QȱO�RȱO�SȱO�TȱO�U)
����V���W�U)0�[ȱO�����ȄNdXdY�S� �L��Z [�� �
�O� �dZ��ȄZdN���j�k�mȱk�nȱk�oȱk�pȱk�q)
����r���s�q)0�vȱk�����Ȅjdtdu�o� �� �L� ��)��	���Mdw ��`�w�x�zȱx�{ȱx�|ȱx�}ȱx�~)
������녀�~)0��ȱx�����Ȅwd�d��|� к� �M� ��)��@Ы���Ldj A瀠�\�]�_ȱ]�`ȱ]�aȱ]�bȱ]�c)
����d���e�c)0�iȱ]�����Ȅ\dfdg�a� й�h t�� �
�]� �dh��Ȅhd\����
��u녔�u녕���Oȱ��P`��
��}녔�}녕���]ȱ��^`H�Z�T)?	@���T;��%����Y�V��U)@��J������[�8��[��U)0�[ȄY�V����Y�UdY��� z�h`H�Z�b)?	@���b;��%����g�d��c)@��J������i�8��i��c)0�iȄg�d����g�cdg��� z�h`H�Z�p)?	@���p;��%����u�r��q)@��J������v�8��v��q)0�vȄu�r����u�qdu��� z�h`H�Z�})?	@���};��%��������~)@��J��������8�����~)0��Ȅ�����Ƃ�~d���� z�h`� `� `H�Z���������������)?
���녚��녛d� �z�h`� �K� � `d��* d�`������ȱ���ȱ���ȱ���)
���녉��녊��)0��Ȅ�d�d���� �d�`H�Z�����L�ꥆ����;��)����������)@��J��������8������)0��Ȅ������Ƌ��d���)����)����
�@����������( ��Ő��* ��戥�Ň� �z�h`H�Z�  [�  t�dNd\��Z�h �� �� �� �� ����Kz�h`H�Z�L� ��M� �d���)?ŗ�D�� �>��
����k���x载�l���ydjdw� �L�M��)�����M �祖���L A� ��z�h`�����������V���p�  ��2���^���� �  ��  ��  
�  
�  v���  v���  B�T���B�T����E�P�_�d�{��������������V� �   �G� �   �f� �    ��V� ��G� �   

		�
	�
	�
�	
	�	

�	
	��	���� <�� K��  �� K��  �� K��  �� Ki�#� T�� _��  Z�� _��  �� _��  �� _��  �� _��  �� Yx�#� T<��  <��     � <�� T��  �� T��  �� T��  �� Gi�#� K�� T��  Z�� ���  �� ��� ��� ��� <�� �<�� �<��  x�� �<�� q��  ��     � ���  �� _��  �� q��  �� �x�� ��  �� �<�� q��  �� _��  �� G�#�  �� q��  �� �x�� ��  Z�� ���     �  �� q��  �� T��  �� C��  �� 8<�� ?��  �� T��  �� d��  �� T<�� _��  �� q��  �� ���  �� <��  x��  <��     �}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�     �}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"���"��"� ��"���"��"� ��"���"��"� ��"���"��"� ��"�     ���"��"� ��"���"��"� ��"���"��"� ��"���"��"� ��"���"�T�"� ��"���"�T�"� ��"���"�T�"� ��"���"�T�"� ��"�     ���"�T�"� ��"���"�T�"� ��"���"�T�"� ��"���"�T�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�}�"�.�"� ��"�     �}�"��"� ��"�}�"��"� ��"�}�"��"� ��"�}�"��"� ��"�}�"�@�"��"�}�"�@�"��"�}�"�.�"� ��"�}�"�.�"� ��"�     �}�"��"� ��"�}�"��"� ��"�}�"��"� ��"�}�"��"� ��"�}�"�@�"��"�}�"�@�"��"�}�"�.�"� ��"�}�"�.�"� ��"�     �T�"� ��"� ��"�T�"� ��"� ��"�T�"� ��"� ��"�T�"� ��"� ��"�T�"� ��"� ��"�T�"� ��"� ��"�T�"� ��"� ��"�T�"� ��"� ��"�     �T�"��"� ��"�T�"��"� ��"�T�"� ��"� ��"�T�"� ��"� ��"� ��"� ��"� ��"� ��"� ��"� ��"� ��"�  Z�"�     � ��� ��� ��� ��� �� ��� ��� ��� ��� ��� ��� ��� �� ��� ��� ��� �Z��     �}(�"�.(�"� �(�"� �(�"� �(�"� (�"� _(�"� K(�"� ?(�"� /(�"� %(�"� (�"� /(�"� /�"� %�"� �"� /�"�     � K�� C�� ?(�"� K�� C�� ?(�"� C�� ?�� ?�"� ?�"� C(�"� ?�"� ?�"� K�"� T�"� _(�"�     � K�C� C�C� ?(��� K�C� C�C� ?(��� C�C� ?�C� ?��� ?��� C(��� ?��� ?��� K��� T��� _(���     � �
�� /d��     � �
�� ���  �� ���  �� ���  �� ���  �� ���  �� ���  �� ���  ��     � �� �� �� �� ?� � ?� � ?� � ?� � ?� � ?� � ?� � ?� � ?� �     �$�/�:�C�L�U�^�e�k�q�~���p���GAMEaaOVER$PUSHaSTART$STAGEaba$NUMBERba$HSCOREba$SCOREaba$STAGEa$PAUSE$READY$BONaTREASURE$aaCONTINUE$aaEND$ ��� ���@�Ђ`����������0���P���p� ������� ���@�Ћ`��������������0���P���p�p�p�p� ��� ���@�Д`����� �`����� �`����� �`����� �`����� �`���`����� �`����� �`����� �`����� � �`� @�@�A�Z				


���������








D D h8h8n8n8VPVPhP  � 0����~x|�����������)Mq�����		C	C	k	����,�,�@�@�T��	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	BV`     



BV`     



BV`     



BV`     



BV`     



                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  W� �r�