�Ń�`����	 I� &� � Â ��� |�L���������d���h�� �l��LW����p���t�� �x���������`    �������p����������l��)�D��������0�  ) ��  )����$��d�L̀�  ) ��  )������������������
��Ą��ń�� � ��`�	��`����� *���)��������
�������� � �ߊH�e�� e������h�`�o��`�  )���8������  )���e�� ����  )���8儐���  )���e�ɇ���`���⁍����܁�������������
��������� ����`	  ���ɠ������ ��o������������`�  )�`����G�����`���0��`ڮ���}]����}a����������������`�   ���o����o����o����o����o�`��i������������i����������������������`�������	��i����`�����������}������`�� ����������d�
�ڽb���c����d <���j���k����dL<��� ����������L@�ZH ;�h ��z�L@�`�r�ƃn�D���������*+,-*+,-*+,-*+,-*+,-�./01./01./01./01./01�	
	
	
	
	
��"#$%"#$%"#$%"#$%"#$%�&'()&'()&'()&'()&'()���� ! ! ! ! !�                    �                    �                    �                    �``҄ބ؄�؄؄؄	�  ��  ��  �*+�45�
�� ���
����
�  �  �L�M�N�O�P�Q���@�9�                                                                @� ��� ���A���� ��� ���  �������������� �������������@���    � ��?���?���� ?� ?� ??��??��??��?? ?? ?? ?? ??     ��� ��� ��������������������<��� �� �� �� ��� ��� ���    � �������  �  �   � � � � � � �   �   �   �������� �    ��?�������������������?������������� ��� �?? �      ?���?���?���?�  ?�  ?�  ?��??��??��?�  �   �   ��� ��� ���    �� ��� ����������������� ��? ��? �� �� ����            �P �� ��� @��.����j�y��                             �  OZ �  �� P��j� �                                                            @  ��  ��  �u  �y  ��  �  ��  �n                T   �  �  G+  �  �  �  t  m�� �� J�  �j                                        ��       �  ��~  '� �
�                                             @  �  @* �
 ��                                                  �� mi  �                                   �j  Y�   ����@F `@� X�� ع�                                       i  '
  g  	      �*          �P �� ��� @�  (�  U� @�9   �   �   �   �   @            �  OZ �  �� P��j� ��  ��� jW j)  j  �  �          @�   �   m   �  @  �  �  p@   �   �   �   �   �   �   @    �  �  Z  �=  y=  X<  i>  �>  �>  i?  �  �               `VZ�����9 `�M �� @�� � 8@f   �                            �  [� �� �� �  ܪ ߤ
 u@*  �   @                        �V� U��  �.  �
  �
� V��@i��� �  l  �                                                 
   (   �?  �  (  8   �   �   �    (�� ��� ��  � �� @�* �K^ ��� ��� �	� হ �[> @�  �         ��  ��  @�   �   ��  �  
�  ��  ��  �  ��  ��  ��   �   �   �        �P �� ��� @�  ��  �  �X ��� p�� |�� �)p �  �          �  OZ �  �� P��j� �                                         P  U ����� ��Y ��b @Ub ��i��� ��  �  �                �   +   �R �� ���
Z�j�Y ��Z ��R ��X �� �j  V         
   8   �  �
 (�o� ��J�Z n*V �)e 8�Y (� �% �� �Z �    �  �  �    (  
�  n� n��k���I�J��^���a �j  P  0     0     .�     .�  n� �{��b��b��{���v@*� �V  P       V  �j �� ��X ��R ��Z�j�Y��
Z � �� �R +  �           �  �j �� �% (� 8�Y �)e n*V�J�Z� �(�o�
  �   8   
      P  �j ��a�^��J���I�k� n� n� 
�  (   � �  �      P  �Z @*���v
P��
P��
@��@�� ��  .�     .�     0     0       �     @  @
 �@
�*����	]@ͤ���@
�* �  @
  @     �              �   
 �@	�%T��*9�A3Tj�* � i �@�                               P   $  @ �*��Z���PU��  �*                                       @ �@� � )Tj�*9�A3T��*@	�% �   
  �                                  �*PU���͐�Z�@�*  @   $   P                                           �   �   �   �   �   �  @�  �                 �   * ��� �G��������_/[ �F: �
 9]. {}�                              �?  �?                                                     T  �?   �                                                     T   �  �   /                                             P   P  �  �      /                                         @  @  �  �  �  �  �                                         �  �  �  �   �                                                P   T     �  �  �                                                P   W  �  �                       �                                                            ����Fk Z � { ��+ �%* �O �� ��; ��<   �                                          �  `  P	  �                                              �  p  �9  X%  P  �                                      �  �:  [�  W�  W�  U�  X9  �                                  �   �  \  �+  �  �  �                                       �
  X=  �  �  �   �   $  @                  h)  � ����������F��ê�����*�����
�������� �  h)  h)  � ����������F��ê�����*�����
�������� �  h)  h)  � ������������F����3����*�����
�������� �  h)  h)  � ����������F��Ϫ���?�*������
������� �  h)                              �  �                                                     �   �  �                                                     �   �  �                                                �   �   �  �  �                                         �  �  �  �  �  @  @                                             �  �  �  �                                                  /  �  �  T                                                     �/  �  �                                                                    �   �  �  �C   �               �   (   
  ��  �  �n���N|��n���V��E	�E��Z|��n                � kU+�
  &  P�@kUP �                                  0  ;�  *�  &�  &�  T                                           �   �   p  Z)  p  �   �                                       �   �  [  [  �  �                                              8  �  p  �  8                                        �   `  |  �	  �/   �                               �  ��  �7  `~ |��� w�  �}  �  � �          
 ��8�#���*�	�f�hB�3�4F>�J���b
�R��ME>��`���I���*(
  H����N  �n  �  ��   
   (   �                                    ���0����?�������      �  ��������?0�����                �  �  �            �  �  �              ��� �� �?  �  �  � �? �� ��? �  �  �  ��? 0�� ���    ��� �� �?  �  �  � �? ��  �?  �  �  � �? �����        0  �  ��������? ��  �?  �  �  �              ���0�� ��? �  �  �  ��?  ��  �?  �  �  � �? �����    ���0�� ��? �  �  �  ��?  �� ��?��������?0�����    ��� �� �?  �  �  �            �  �  �              ���0����?��������? �� ��?��������?0�����    ���0����?��������? ��  �?  �  �  � �? �����                                                                     ��D(\� ͰcfeY�}� �Z��Yp9 ���!�� (]�Ͱc�feY}� �Y��Yp9 ��� ��0\� B�c�eY"إ 3X�H@p9�� ��\��@�c�eY� 0X�@@s9 ��  $R  L� @1`  !I @�$  P    ��     �  �@  `Y  !  � @@	  ��           �   �   `          H   F   �  ��  ��  `�  `�  ��  ��i   �   �   �   �   �   �  ��  `��?X�_�k�@� ?��Է���P���� (   � �Q
 `�* �. F� Q�
 �� �� ��  �  �/  �+  �  �
  �                                 �   �   �   �   \      |   �   \  ~�  P �  �T�U�CuU��U�^���~��mp�j{r�j�}�j�}�k{n�m�W���Aݶ]@����@���U����Wj�[~U����������������\��\�����u��_��� ��� �  �   �   /   +      
                �   �  w  3  3                                                                ��   �   �                 ��� pt�����빪���@ǥ��ǔ���P��@]�����z�Gۯ��n�Х�0n��psk�pn�W���A��9?�z���ސm�^W��F�.��Ӯ���n��[n[��_���u�Z�Z�k@���Uz����E����Ѫ���V[�ZV��UV�VV�XVx `W� ��w  �  �             	   /   �   �
  ��  �� ��5 �k� �[U�VU ����uհy�e,u�\�eYkYe�G]�SWmYW[�G��QWk�U[lՖ�ey԰u��[�e �Zey�eu�Y�eYeYe�G]�YVmYGY�GV�QWY�U[�Q��U�Q�e�U�e�e�y�eYu�eY�G�eYW��GY�YV��GY��V�Q�Y�U��Q��U�Q�e�U��e��y�e�u���eY�Yem����
��W)�UU�jAU�j �n �nA��U�������������W���V5��]��]���V��Z��k�:鯿:���鿪�鿪������������꫿��Z���V��?�k�:�Z��V�  ��                                                            �����@]��P�ǔ��ǥ����@빪����� pt� ���                   �   ����.��n�Ӯ�F�.���l�^W��ސ?�z�A��9���pn�Wpsk�0n���Х����nz�G�} ��y �W��V��V���V[�UV��_V���������F�U��k@��Z麪Z����u[��_�VU�_U�~� ��5 �� ��  �
  �   /   	             �   �  w     \   �   |      \   �   �   �   �                            �Aݶ�W��n�m}�k{}�j�r�j�p�j{~��m^����U�CuU��U� �T �   P  ~���� ��� ��_���u�������������������[~U��Wj�U���@������]@�3  3  w  �  �                
      +   /   �   �   �    ��  ��  `�  ��  ��  ��   F   J      (   `   �   �   �        ���P�����Է ?��@��_�k��?h�  `�  ��   �   �   �   �   i   �  �
  �  �+  �/  ��  �  �� �� ��
 F� �+ `�. ��
  �  (                                                              	
	
	
	
	
                                                             ! ! ! ! !                    "#$%"#$%"#$%"#$%"#$%&'()&'()&'()&'()&'()                    *+,-*+,-*+,-*+,-*+,-./01./01./01./01./01                ��������������������������������������������������������������ﯪ�ꖪU�U�U�� ������Z�ZiVUTQP@�����������UQU 믫������V�UeU��E�fwV3Fwe����R����wW3wW����U��ݪ�U� vUު���Tuݥ�a�owm�o�eݩwJUK�-�UUUUUUUU��U�U��� �U�U�Uժ*tUDU��  tUDUTU���R�t?E@UUUUUUU���fo��V�z�~A목k�k����꪿Un���A� �E������UoA��U���Z��n�����������?�������k�����?�A�������m��cA�����n�z�o�����?��к���m��cA�������?���ᑻ����A�?���꾑k����cA�m䯿����?����o�z���n���~Ay���U�o�f��n��Uꪥ����k�k��oA�U����E� �A�������nZ���U���  UUUUUUյ-UK�* �U�U�U��� �Uժ�  tUDUTU��  tU��  UUUUUU?u�D�R�R�wDwfwV3Fwew�wU�w�w�wW3wWw�w�Du�ݪ�U� vUު���wJݩ�%�owm�o�aݥ �U�U�U������P@TQVUZiZ������� QU�U����������eU�U�V������믪��������������������������������������������������������������                                                                  UU  UU  UU  UU  UU  �W  �W  �W   W   T   T   T   T   T   T   TUUU�U=U�U�U�U�U�U���UU��UU��UU��UU��UU��U���U���U���U���U���U�PUUP�UUP�UUS�UU_�UUU�U�U�UUU�UUU�UUU�UUZ�U�Z�UUZ�UUZ�UU[�UU_�UUU%  U�  U� U�
 U�* ���@U���U���U��U�������U���U���U��U���U��� UUU@WUU�WUU�WUU�WUU�W���WUU�WUU�WUU�WUU�W���WUU�WUU�WUU�WUU�WUUT@Wp�W|�WU�WU}�WUu�WUU�WUU�WUU�WUU�WuU�W�U�W�W�W�_�W��W��UWUUWUUUWUUUWUUUWUUUW�VUW�^UW�_UW�_UW�_UW�WUWUUUWUUUWUUUWUUUWU�                U   U   U   U   U   U                      �   �                                                        ������������� ��� ��� � � � �                                  ����������������������������                                ����j�㪪�㪪�⪪�⪪jb��������                                ��������������ꩪ�������������                                ���������������������*���
 ��                                ꪪ*���
������ ��* ��
 �� ��                                    @�  ��  ��  �  �   �   �   ��  ��  ��  �   �  ��  ��  @�     �� ���A����?������  � �� �������������� �� �� ��       �? �� �������?���?���??��??<�?? �?? �?? �?? �?? �?? �    ����������  �  �  ��� ��� ��� �  �  �  ���������     ��  �� ��? ��?�? ��? ��? ��? ��? ��? ��? � ��? ��? �� ��     �������������������������?���������� �?� �� �� � �    ��?���?���?�?  �?  �?  ����������?  �?  �?  ���?���?���?�    �  �?  �   �   �   �   �  �  �?  �  �  �?  �?   �   �                                                                  	
                     !"#$%&    '()*+,-./0123456        789:;<=>            ?@ABCDEF             GHIJKL                                                                                                                                                                                                                                        @ P T U     VPe�Z�ZjTU @UUUUQU  �DUDYPB U  �     UE%XU �`             U        @ @ � � hPET�dY�Je�e�Zj�
j��U�P�RTR�E@PhP�yIjD��Z�A�D�ET�A� � ��������@�-C|A�PEe��Z�i@           *  � �@���������k�������oVo�U��zVjJ@*��ښ�Z�V��URUE��f��@A��a��V�V�Z�j���*V&U�YEYQ�f`A�BfA��	�	zP~ � ����^�   � � � �������  �?�?�?��������           � ��  ����?�?�*��   � � � � � � �  �?�?��������"  �����������  ������
 
   ���������Ϩ���  ���/�?�?�*�*   <�?�?�?�?�*�*   � ����*�*  ����?��������  ��������O

*  ������?������  ������
pq����������?�?U*�*�?���������P�
���?�?�?�QU�������?�?�?� @  (�������U�
�*�?��������PU�������� ��� 
 
 ������TE��������������U�  ? � ��U�*�*�?�?�?�? <U�*�*����  @U�
�?������?U �����������Ǽ�PU����?����� � �����o   ������ � Z i T  f��ji e U U   �'�m�Z����@B�V  Q� V� Q @   D@F   `  � @P�@�  e�DE@Z�QP  �*�
v
����  � � @          eUVPZ���T�EPd@��j�j�jiE�V�� � QEF�R VQ      Q A�@� @@Y�VJDED@%�����eUU�  %         � P            ZUUPPP U P     E DUTU P@@APTTUUU�UiUYQDUUU   QEU          �Ŕ�`��敭��
������������������d� .� �� (� \� �� �� E�旭�	 "� P� �斥�)��� z� �� [�����4� ��	����ؐ��LK�������������������`������������������`��*��&��i8��� �����}��8��݌�����o��`   ��������� ����`������������ Ѷ��`�8��
��8��
��o�����������LX�`���o�`����m����#�m������� ˷`)#1Q.�� 
��:���;��l ~�N�B�B���)� ˷LN���0`���������� �復��ɥ�������ɥ�`�o������`��)�����8������`�o��`��0`��i1��������� 
��X���Y���� ��`��8����� � Jf���8����� � Jf���
&��
&��I�i����I�i����Ŝ&�)�����` ��#����yK�8������i<8������`0   ����������� m���`��i28�� �I��i88���<�o��������  �� X���
��ĸ��Ÿ�����8������ �����`̸ظظ�	
	
	
��iP���i ��@��,� >���iP���iP��0��$� >���iP���ip��@��,��8�����8�������LX�`��0`�������������L�߭�0`��͎����L���N�����iͥ����L�����0��������8���`��m��������8���`��m���`�.������ȱ��I���`����E���U�$�
��L;��8�����������m��`ɪ��L;��i]H�8��h��`��0,���բ� *֭��?��o���������`�N��L0�`� Z�)�i� Z�)/im�� Z�)/im�� Z�)������
����������� ��` %(CF#:+. %(&CF#.7(&CF#F#.7CF#7:+.!����������������Q�P��\��]��^L�� ֩ �"��#���������� Sŭ���'���	������ Sũ��	� ;��� |�L�����	�� ���� Sũ��	� ;��� |��H�de�� e������h�L�******************�*                *�*                *�*                *�******************�LEVEL : FINAL LEVEL :   abc� defg�hijkl�mnopq�rstuv� wxyz�  {|}�`�b�b�b�9�:�e, the string must be null-terminated and  have the DOS filename format. If  lpFilename  contains a handle, the handle must be in the low-order word; the high-order word must be zero.   *      �  *   '    � �&K!��!� ��   �   �   *   �   -   ,� �&KP!��~�!� � ��� Return Value  The return value specifies the outcome of the function. It is nonzero if the function is successful. Otherwise, it is zero.  *      �   *   '    � �&K!��!� ��   V    *   V  E   \� �&KP!��~�!� � ��_  � �� � �  � ��� Comments  Any application that adds or removes fonts from the Windows font table should notify other windows of the change by using the   SendMessage  function with the  hWnd  parameter set to -1 to send a   WM_FONTCHANGE  message to all top-level windows in the system.  A    V  M  9   D� �&K!��!� �� � ��  � �����  The  RemoveFontResource  function may not actually remove the font r�Ԣ� *֜��f���� zũ��������� Sũ��������� Sũ ��������� Sŭ  )�� ��`��������H�e�� e������h�LN��N�� � ��L �PLAY START   (C) 1992   Thin Chen Enterprise  ��6���� zŜ������ ��������� Sŭ  I��`���Ȑ�H�e�� e������h� ��L���)���� ��F�� JJ��P�^JJ�	 ?�����L�)����� ����� ��U��0��U����p���JJ�	� JJ�
 1ߊH�e�� e������h���L��
���������d��LSŰ�Łځ���.�                      In A.D. 2X00 alien  Saya Empire secretly built a .Time space. Frontier Post on the Moon. intentionally  intrude the earth... 
��X���Y��d��LS�h�}�������т��� In order to defeat  the alien's intrusi- on. the Earth Defen- se Arms has launched an unprecedented ou- ter space war with   the alien Saya Empi- re.................. ���	�&�y�w���z�x������������F���n��������� zũf������� ��	������  I��`L���H�2e�� e������h�`��)���������}Y���F����}]�� ��n���������a������� �� W���
��� ����)�����)����柊H�e�� e������h�����Lk��)�L`���)����� C���� ��X��0��X��������JJ�	� JJ�
 1���L`�����������������������������������������������	
��  I���H�e�� e������h����  I���`
��c���d���� ����������L̈́ZH ;�h ��z�L̈́`���H�e�� e������h�� ��@�� JJ����PJJ�	 �ީ ��@��PJJ�����JJ�	 ����`���H�e�� e������h�� ��@�� JJ����PJJ�	 �ީ ��@��PJJ�����JJ�	 ���г`�S�� ��O��0��O��P� ���JJ�	� JJ�
 �ީ0��O��`��O����Q���JJ�	� JJ�
 1��б`���� ��@��0��@��� ���JJ�	� JJ�
 1ߩ ��^��0��^��������JJ�	� JJ�
 ���б`�	�H��ȑ����h��i0��i ���L?�`                                                            	
                    !"#$%&'()*+,-./0123456789:;<=      >?@ABCDE            FGHIJKLM             NOPQRS                                                                                                                                                                                                                                        @ P T U     VPe�Z�ZjTU @UUUUQU  �DUDYPB U  �     UE%XU �`             U        @ @ � � hPET�dY�Je�e�Zj�
j��U�P�RTR�E@PhP�yIjD��Z�A�D�ET�A� � ��������@�-C|A�PXdXԙ�Z�iX           *  � �@���������k�������oVo�U��zVjJ@*��ښ�Z�V��URUE��f��@A��a��V�V�Z�j���*V&U�YEYQ�f`Y�RfQ��I�IzEPR^ � �nV�V�  ���?�?�?̪�  ������
�*   � � � � �  *  � � � ����
   �������������  ����      �?�?�?�?�?�*�*  �?������ � � �  �������
�   ?�?�?�?�?�*�*  ���������� � �  ?�?�?�?�?�*�*�   ? �����𪨪�  �<������������   ���?�?�����  ?�?�������*��  ?�?�?�?�?�(� �  ���?����ê
�*       
       � � � � � �W+�*�����������P�*��������?�?�  �������������U�
�*�?�?������UU������������ �  �
�
����� T�*�*�?�?�?�?�?PT����������?�?E*���� ����U�*�*�?�?�?�? ? P � �����������U*�*
???�?�?�?�T� � � �� ? UT�������������<U ��(?�?��� �UU��������?���@

???�?���UU����������?�           ������ � Z i T  f��ji e U U   �'�m�Z����@B�V  Q� V� Q @   D@F   `  � @P�@�  ei�eEXZ
�aP  �*�
v
����  � � @          eUVPZ���T�EPd@��j�j�jiE�V�� � QEF�R VQ      Q A�@� @@Y�VJXET@e�Y����eUU�  %         � P            ZUUPPP U P     E DUTU P@@APTTUUU�UiUYQDUUU   QEU                                                                                          	
 !"#$%&'()*+,-./0123456"#789:;<=>-.?@ABCDEFGHIJKLMNOPQR                                                                                                                                        ������������������������������������������������������������������������������������k���k��������������������������������_�W�U�����V_e�Z�ZjTU UUUUQU  �DU�DYPB U  �������U�E�XU �`��������������U�������{F���������������������k_EW�dY�Je�e�Zj�
j��U�P�RTR�E@PhP�yIjD��Z�A�D�ET�A� � ��������@�-C|A�P��E�e��Z�i@��������������������/鿞��/�����������A����������������������k�������oVo�U��zVjJ@*��ښ�Z�V��URUE��f��@A��a��V�V�Z�j���*V&U�YEYQ�f`A�BfA��	�	zP~�����������^��ۿ�������`�e������e�.��@n���Z��������������Aݯ����������������Z{�fk&kk��U����������d�!�A�V��~�J����!�	�fzfA%�A A� TVne��od�E�UY��@�BzN�A�q aUR��������g�v���w*����e`�����������A.�e�����������������������ꫪ�������^�����	gYUP*Q*F��@� � PAE�~eQVU U   P @� X@T@���$A(�EjnY!Q ��WZ�Z�f*`�$U]�������֯�o�k�믪���������Z�i�WIEf��ji e U U ���'�m�Z����@B�V Q� V� Q @AQ D@F  ``  � @P�@�%Qe�DE@Z�QP�����v�����������[~����ށ��-/v�������������j��������������T����������������eUVPZ���W�E_d��j�j�jiE�V�� � QEF�R VQ      Q A�@� @@Y�VJDED@%�����eUUU��Y�e�����������o~��������[~�ߪ���������������������������������_������������ZUUP_P�U�_���� E DUWU�_@@APTTUUUU�UiUYQDUUU�U���Q�E�U�����������                                                                                	
 !"#$%&'()*+,-./012345 6789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVW X)YZ[\]^_`abcdefg   hijZklmnopqrstuvw  xyyz{|}~����������                                                                                ����������������                       �    B�U ��
j  TUP�
 � PTUTUUUUU  ��UZU�U�UEUE ��U�����j�YY��� Ui��������jU��     j ���jV�              �U`U`�X�XUXUXUZUPUTUUU��������UUUeUZ�Z�Z�Z�[�[ AAA@@@Q�PiTUP�� �UU��j������ifjjjjV��������j�V���U� j��+�/��                      ��        * � j��������������������������������[�k�k����������QUU�Z�j������UUUTVUV�j���j�����U��U�U�V�[���U�U�Uꕪ�������������������ﺿ    ? ? � � ��V���V���V��������������������������������������������������������������������j�������������o������������������������������ﾾ������������� � ���������V���V��                     �    @f������                    � � � � @        ����������@�    �����U�U�U�V V�WUU�o�����?�?e~U]��U�_U�UTVA������� @ @    ����������[�Y����������?�V���V���V�             P �    U0B                � � � 0 0 � 0 0�Z�f�frf2f:f�fr��	���]����������������	���           � ` ��W F F�AhPU TTUeUuU��jUUUUUUQ                  @ @ @ @ @�a���������Y������������������?�?�?�?�?�?�?�?��V���V���V@j@������������ٕ�0����Y�	�	�	�Y M d ] U � � 0 0 � 0 0 � 0f:f2f�fzf2f2f�fr���_��������������	����	�[�k��        %f                �       � �   @-UfUVUUUAU�U�[AVU         P P T � � �@�@������������������?�?�����������������������������	�	�	�Y�	�	�	�YTT����0�0!0!��9���f2f:f�frf:f2f�fz�]������_������������ۑK�+���ˑ+��j%�&�j��B�-��B�9  �j1���2P2��� @    
  ) & ZU^UVUVUVUVVV                     @ T � �@�P�P�T�U����������V������U�U�fm�����U�U�fm����������������� �UĪ��� �UĪ�� xUɪ�k �U�j��f2f2g�grg2������������ꪪ������������6�I�+���K�)�ۑ˓+)��CC))��BB9)��B2P2�r�rQr�����* ) & * ) & + . V V XXU�U �       @DUUUUUVU�Z �T�U�U�UUUUUUUUUU������������U�U����������������UlU�Y��lUlV�e�U���f�j۪ۦ�f�j۪��	�	�	�Y�	�	�	�	� �UĪ��� �UĪĪ Ui��� hU���z��������������������v���2r���2v����p��*ț�J�)ț�IB)-ԴBB))��BB+���W�W�W�W�W�W�* � ������VUVUXUXUXUXU`U`UUUUUUUU]U5UU@���eB��Z�T�T]U�����U��U�U_UUUUU�     U UUUU                                                                   �   @      �  ��  �7  m?  �+  t�  `x� ��  �  <       UU���oU���_U���U�?TV�?e~U]AUeQ Uu U� �j UU UU  U  U  UU��UAU�UQUUU��U�~YV�?�~��BUeQ Uu U� �j UU UU  U  U  UU��UUU�UUUUUUUU���V��n��EUU@UUEUUU UUU UU UU UU  U  U                    	
                                                                                                                                                                                                                                                                                                                                                                                                  UU�o�����?�?e~U]��U�_U�UTVAUUUAUQU�~�?�~����U�UU�UYVBUUUUUUUU������UU��U�UUUU�VnE@UeUuU��jUUUUUUQ           UUUUUUUUUUUUUUEU U         &KPтS~�!��� � �� � �� Parameter   Type/Description   L  �   W   L  U   |� �&KR�тS~�!��� � �� � �� � �� � �U  � �� � �� hDC   HDC   Identifies the device context.   nSavedDC   int   Specifies the device context to be restored. It can be a value returned by a previous   SaveDC  function call. If  nSavedDC  is -1, the most recent device context saved is restored.   *      L  *   '    � �&K!��!� ��   �   �   *   �   -   ,� �&KP!��~�!� � ��� Return Value  The return value specifies the outcome of the function. It is TRUE if the specified context was restored. Otherwise, it is FALSE.  ,      �   ,   (   "� �&K!��!� ���    2      ,   2   !   �  Q  S  RGB utility macro/      2   /   (   "� �&K �!� � �� RGB   z   5   /   z   E   \� �&KP!��~�!� � �� � � � � � � � �� Syntax   COLORREF  RGB( cRed ,  cGreen ,  cBlue )   �   t   z   �   (   "� �&K�!��!� �� This macro selects an RGB color based on the parameters supplied and the color capabilities of the output device.  *      �   *   '    � �&K!��!� ��   W       *   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description     �   W     T   z� �&KR�тS~�!��� � �� � �� � �� � �� � �� � �� cRed   BYTE   Specifies the intensity of the red color field.   cGreen   BYTE   Specifies the intensity of the green color field.   cBlue   BYTE   Specifies the intensity of the blue color field.   *        *   '    � �&K!��!� ��   q   D   *   q   -   ,� �&KP!��~�!� � ��� Return Value  The return value specifies the resultant RGB color.  *      q   *   '    � �&K!��!� ��   �   �   *     -   ,� �&KP!��~�!� � ��� Comments  The intensity for each argument can range from 0 to 255. If all three intensities are specified as 0, t7�5 a�5 ��5 he result is black. If all three intensities are specified as 255, the result is white.  �   �     �   <   J� �&K!��!� ��)  � ��*  � �����  For information on using color values in a color palette, see the descriptions of the   PALETTEINDEX  and   PALETTERGB  macros, earlier in this chapter.    3      �   3   !   �  R  U  RoundRect function5      3   5   (   "� �&K �!� � �� RoundRect   �   G   5   �   ]   �� �&KP!��~�!� � �� � � � � � � � � � � � � � � � �� Syntax   BOOL  RoundRect( hDC ,  X1 ,  Y1 ,  X2 ,  Y2 ,  X3 ,  Y3 )   �   �   �   �   (   "� �&K�!��!� �� This function draws a rectangle with rounded corners. The interior of the rectangle is filled by using the selected brush, and a border is drawn with the selected pen.  *      �   *   '    � �&K!��!� ��   W       *   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   ,  �  W   ,  �   � �&KR�тS~�!��� � �� � �� � �� � � � �� � �� � � � �� � �� � � � �� � �� � � � �� hDC   HDC   Identifies the device context.   X1   int   Specifies the logical  x -coordinate of the upper-left corner of the rectangle.   Y1   int   Specifies the logical  y -coordinate of the upper-left corner of the rectangle.   X2   int   Specifies the logical  x -coordinate of the lower-right corner of the rectangle.   Y2   int   Specifies the logical  y -coordinate of the lower-right corner of the rectangle.   �   �   ,  �   F   ^� �&KR�тS~�!��� � �� � �� � �� � �� X3   int   Specifies the width of the ellipse used to draw the rounded corners.   Y3   int   Specifies the height of the ellipse used to draw the rounded corners.   *      �   *   '    � �&K!��!� ��   �   �   *   �   -   ,� �&KP!��~�!� � ��� Return Value  The return value specifies whether the rectangle is drawn. It is nonzero if the rectangle is drawn. Otherwise, it is zero.  *      �   *   '    � �&K!��!� ��   �   �   *     E   \� �&KP!��~�!� � �� � � � � � ���5 5 ?�5  � �� Comments  The width of the rectangle specified by the  X1 ,  Y1 ,  X2 , and  Y2  parameters must not exceed 32,767 units. This limit applies to the height of the rectangle as well.  p   G     p   )   $� � !��!� ����  The current position is neither used nor updated by this function.   !       p   !   !   H   ��������'      !   '   $   � �&K ��� ��   0      '   0   !   �  S  V  SaveDC function2   
   0   2   (   "� �&K �!� � �� SaveDC   X      2   X   9   D� �&KP!��~�!� � �� � � � �� Syntax   int  SaveDC( hDC )   9    X   9  .   .� �&K�!��!� � � �� This function saves the current state of the device context specified by the  hDC  parameter by copying state information (such as clipping region, selected objects, and mapping mode) to a context stack. The saved device context can later be restored by using the   G      9  G   .   .� �&K!��!�Q  � ����  RestoreDC  function.   W       G   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   r   :   W   r   8   B� �&KR�тS~�!��� � �� � �� hDC   HDC   Identifies the device context to be saved.   *      r   *   '    � �&K!��!� ��   �   d   *   �   -   ,� �&KP!��~�!� � ��� Return Value  The return value specifies the saved device context. It is zero if an error occurs.  *      �   *   '    � �&K!��!� ��   �   `   *   �   3   8� �&KP!��~�!� � �� � �� Comments  The  SaveDC  function can be used any number of times to save any number of device-  =      �   =   )   $� �&K!��!� ���� context states.    :      =   :   !   k  U  W  ScaleViewportExt function<      :   <   (   "� �&K �!� � �� ScaleViewportExt   �   O   <   �   Q   t� �&KP!��~�!� � �� � � � � � � � � � � � �� Syntax   DWORD  ScaleViewportExt( hDC ,  Xnum ,  Xdenom ,  Ynum ,  Ydenom )   �   s   �   �   (   "� �&K�!��!� �� This function modifies the viewport extents relative to the current values. The formulas are written as follows:  XXXXXXXXXXXXXXXXXXXXXP�5 �5 :�5 �   �   �   �   ,   *� �&K!��!� �������  xNewVE = (xOldVE x Xnum)/  X  denom yNewVE = (yOldVE x Ynum) / Ydenom  The new extent is calculated by multiplying the current extents by the given numerator and then dividing by the given denominator.   W       �   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   �  r  W   �  �   � �&KR�тS~�!��� � �� � �� � �� � � � �� � �� � � � �� � �� � � � �� � �� � � � �� hDC   HDC   Identifies the device context.   Xnum   int   Specifies the amount by which to multiply the current  x -extent.   Xdenom   int   Specifies the amount by which to divide the current  x -extent.   Ynum   int   Specifies the amount by which to multiply the current  y -extent.   Ydenom   int   Specifies the amount by which to divide the current  y -extent.   *      �  *   '    � �&K!��!� ��   �   j   *   �   -   ,� �&KP!��~�!� � ��� Return Value  The return value specifies the previous viewport extents (in device units). The previous   �   [   �   �   2   6� �&K!��!� � � � ���� y -extent is in the high-order word; the previous  x -extent is in the low-order word.    8      �   8   !   M  V  X  ScaleWindowExt function:      8   :   (   "� �&K �!� � �� ScaleWindowExt   �   M   :   �   Q   t� �&KP!��~�!� � �� � � � � � � � � � � � �� Syntax   DWORD  ScaleWindowExt( hDC ,  Xnum ,  Xdenom ,  Ynum ,  Ydenom )   �   q   �   �   (   "� �&K�!��!� �� This function modifies the window extents relative to the current values. The formulas are written as follows:  �   �   �   �   ,   *� �&K!��!� �������  xNewWE = (xOldWE x Xnum) / Xdenom yNewWE = (yOldWE x Ynum) / Ydenom  The new extent is calculated by multiplying the current extents by the given numerator and then dividing by the given denominator.   W       �   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   �  r  W     �   � �&KR�тS~�!��� � �� � �� � �� � � � �� � �� � � � �� �F�5 ��5 ��5  �� � � � �� � �� � � � �� hDC   HDC   Identifies the device context.   Xnum   int   Specifies the amount by which to multiply the current  x -extent.   Xdenom   int   Specifies the amount by which to divide the current  x -extent.   Ynum   int   Specifies the amount by which to multiply the current  y -extent.   Ydenom   int   Specifies the amount by which to divide the current  y -extent.   *        *   '    � �&K!��!� ��   �   �   *   �   9   D� �&KP!��~�!� � �� � � � �� Return Value  The return value specifies the previous window extents (in logical units). The previous  y -extent is in the high-order word; the previous  x -extent is in the low-order word.  ,      �   ,   (   "� �&K!��!� ���    8      ,   8   !   �  W  Y  ScreenToClient function:      8   :   (   "� �&K �!� � �� ScreenToClient   s   4   :   s   ?   P� �&KP!��~�!� � �� � � � � � �� Syntax   void  ScreenToClient( hWnd ,  lpPoint )   S    s   S  C   X� �&K�!��!� � � � � ��  � �� � �� This function converts the screen coordinates of a given point on the display to client coordinates. The  ScreenToClient  function uses the window given by the  hWnd  parameter and the screen coordinates given in the   POINT  data structure pointed to by the  lpPoint    �   �   S  �   (   "� �&K!��!� ��� parameter to compute client coordinates, and then replaces the screen coordinates with the client coordinates. The new coordinates are relative to the upper-left corner of the given window's client area.   W       �   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description     �   W     O   p� �&KR�тS~�!��� � �� � �� � �� � ��  � ��� hWnd   HWND   Identifies the window whose client area will be used for the conversion.   lpPoint   LPPOINT   Points to a   POINT  data structure that contains the screen coordinates to be converted.   *        *   '    � �&K!��!� ��   C      *   Q   -   ,� �&KP!��~�!� � ��� Return Value  None.  XX��5 �5 �5 *      Q   *   '    � �&K!��!� ��   �   [   *   �   3   8� �&KP!��~�!� � �� � �� Comments  The  ScreenToClient  formula assumes the given point is in screen coordinates.  ,      �   ,   (   "� �&K!��!� ���    2      ,   2   !   P  X  Z  ScrollDC function4      2   4   (   "� �&K �!� � �� ScrollDC   �   d   4   �   ]   �� �&KP!��~�!� � �� � � � � � � � � � � � � � � � �� Syntax   BOOL  ScrollDC( hDC ,  dx ,  dy ,  lprcScroll ,  lprcClip ,  hrgnUpdate ,  lprcUpdate )   d  *  �   d  :   F� �&K�!��!� � � � � � � �� This function scrolls a rectangle of bits horizontally and vertically. The  lprcScroll  parameter points to the rectangle to be scrolled, the  dx  parameter specifies the number of units to be scrolled horizontally, and the  dy  parameter specifies the number of units to be scrolled vertically.  *      d  *   '    � �&K!��!� ��   W       *   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   �  6  W   �  �   � �&KR�тS~�!��� � �� � �� � �� � �� � �� � �� � �� � �   � ��� � �� � �   � �� � �� hDC   HDC   Identifies the device context that contains the bits to be scrolled.   dx   int   Specifies the number of horizontal scroll units.   dy   int   Specifies the number of vertical scroll units.   lprcScroll   LPRECT   Points to the   RECT  data structure that contains the coordinates of the scrolling rectangle.   lprcClip   LPRECT   Points to the   RECT  data structure that contains the coordinates of the clipping rectangle. When this rectangle is smaller than the original pointed to by  lprcScroll , scrolling occurs only in the smaller rectangle.   �  �  �  �  U   |� �&KR�тS~�!��� � �� � � � �� � �� � �   � ��� hrgnUpdate   HRGN   Identifies the region uncovered by the scrolling process. The  ScrollDC  function defines this region; it is not necessarily a rectangle.   lprcUpdate   LPRECT   Points to the   RECT  data structure that, upon return, co��5 ��5 �5 ntains the coordinates of the rectangle that bounds the scrolling update region. This is the largest rectangular area that requires repainting.   *      �  *   '    � �&K!��!� ��   �   �   *   �   -   ,� �&KP!��~�!� � ��� Return Value  This value specifies the outcome of the function. It is nonzero if scrolling is executed. Otherwise, it is zero.  *      �   *   '    � �&K!��!� ��   �  x  *   �  K   h� �&KP!��~�!� � �� � � � � � � � � � �� Comments  If the  lprcUpdate  parameter is NULL, Windows does not compute the update rectangle. If both the  hrgnUpdate  and  lprcUpdate  parameters are NULL, Windows does not compute the update region. If  hrgnUpdate  is not NULL, Windows assumes that it contains a valid region handle to the region uncovered by the scrolling process (defined by the  ScrollDC  function).  �   �   �  �   9   D� �&K!��!� ��Z  � �� � ����  An application should use the   ScrollWindow  function when it is necessary to scroll the entire client area of a window. Otherwise, it should use  ScrollDC .    6      �   6   !   �  Y  [  ScrollWindow function8      6   8   (   "� �&K �!� � �� ScrollWindow   �   U   8   �   Q   t� �&KP!��~�!� � �� � � � � � � � � � � � �� Syntax   void  ScrollWindow( hWnd ,  XAmount ,  YAmount ,  lpRect ,  lpClipRect )   �  �  �   �  L   j� �&K�!��!� � � � � � � � � � � � � �� This function scrolls a window by moving the contents of the window's client area the number of units specified by the  XAmount  parameter along the screen's  x -axis and the number of units specified by the  YAmount  parameter along the  y -axis. The scroll moves right if  XAmount  is positive and left if it is negative. The scroll moves down if  YAmount  is positive and up if it is negative.  *      �  *   '    � �&K!��!� ��   W       *   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   )  �  W   5  }   ̀ �&KR�тS~�!��� � �� � �� � �� � � � �� �Y�5 ��5 @�5  �� � � � �� � �� � �   � �� � �� hWnd   HWND   Identifies the window whose client area is to be scrolled.   XAmount   int   Specifies the amount (in device units) to scroll in the  x  direction.   YAmount   int   Specifies the amount (in device units) to scroll in the  y  direction.   lpRect   LPRECT   Points to a   RECT  data structure that specifies the portion of the client area to be scrolled. If  lpRect  is NULL, the entire client area is scrolled.     �   5    G   `� �&KR�тS~�!��� � �� � �   � �� � �� lpClipRect   LPRECT   Points to a   RECT  data structure that specifies the clipping rectangle to be scrolled. Only bits inside this rectangle are scrolled. If  lpClipRect  is NULL, the entire window is scrolled.   *        *   '    � �&K!��!� ��   C      *   C   -   ,� �&KP!��~�!� � ��� Return Value  None.  *      C   *   '    � �&K!��!� ��     �   *     3   8� �&KP!��~�!� � �� � �� Comments  If the caret is in the window being scrolled,  ScrollWindow  automatically hides the caret to prevent it from being erased, then restores the caret after the scroll is finished. The caret position is adjusted accordingly.  �  |    �  f   �� �&K!��!� �� � ��  � ���  � �� � ��� � � � � � � � � � ��  The area uncovered by the  ScrollWindow  function is not repainted, but is combined into the window's update region. The application will eventually receive a   WM_PAINT  message notifying it that the region needs repainting. To repaint the uncovered area at the same time the scrolling is done, call the   UpdateWindow  function immediately after calling  ScrollWindow .  If the  lpRect  parameter is NULL, the positions of any child windows in the window are offset by the amount specified by  XAmount  and  YAmount , and any invalid (unpainted) areas in the window are also offset.  ScrollWindow  is faster when  lpRect  is NULL.  p    �  |  Q   t� �&K!��!� �� � � � � � � � ��  � �� � ����  If the  lpRect  par��5 ��5 @�5 ameter is not NULL, the positions of child windows are  not  changed, and invalid areas in the window are  not  offset. To prevent updating problems when  lpRect  is not NULL, call the   UpdateWindow  function to repaint the window before calling  ScrollWindow .    7      |  7   !   �  Z  \  SelectClipRgn function9      7   9   (   "� �&K �!� � �� SelectClipRgn   m   .   9   m   ?   P� �&KP!��~�!� � �� � � � � � �� Syntax   int  SelectClipRgn( hDC ,  hRgn )     �   m     (   "� �&K�!��!� �� This function selects the given region as the current clipping region for the specified device context. Only a copy of the selected region is used. The region itself can be selected for any number of other device contexts, or it can be deleted.  *        *   '    � �&K!��!� ��   W       *   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   �   d   W   �   F   ^� �&KR�тS~�!��� � �� � �� � �� � �� hDC   HDC   Identifies the device context.   hRgn   HRGN   Identifies the region to be selected.   *      �   *   '    � �&K!��!� ��   �   i   *   �   -   ,� �&KP!��~�!� � ��� Return Value  The return value specifies the region's type. It can be any one of the following values:  *      �   *   '    � �&K!��!� ��   J      *   J   7   @� �&KPтS~�!��� � �� � �� Value   Meaning     �   J     5   <� �&KR�тS~�!��� ��������� COMPLEXREGION New clipping region has overlapping borders.   ERROR Device context or region handle is not valid.   NULLREGION New clipping region is empty.   SIMPLEREGION New clipping region has no overlapping borders.    *        *   '    � �&K!��!� ��   �   z   *   �   3   8� �&KP!��~�!� � �� � �� Comments  The  SelectClipRgn  function assumes that the coordinates for the given region are specified in device units.  Y  (  �   e  1   4� �&K!��!� ��
  � ���  Some printer devices support graphics at lower resolutions than text output to increase speed, but at the expense��5 \�5 �5  of quality. These devices scale coordinates for graphics so that one graphics device point corresponds to two or four true device points. This scaling factor affects clipping. If a region will be used to clip graphics, its coordinates must be divided down by the scaling factor. If the region will be used to clip text, no scaling adjustment is needed. The scaling factor is determined by using the   GETSCALINGFACTOR  printer escape.  ,      e  ,   (   "� �&K!��!� ���    6      ,   6   !   B  [  ]  SelectObject function8      6   8   (   "� �&K �!� � �� SelectObject   r   3   8   r   ?   P� �&KP!��~�!� � �� � � � � � �� Syntax   HANDLE  SelectObject( hDC ,  hObject )   �  [  r   �  @   R� �&K�!��!� � � � � � � � � �� This function selects the logical object specified by the  hObject  parameter as the selected object of the specified device context. The new object replaces the previous object of the same type. For example, if  hObject  is the handle to a logical pen, the  SelectObject  function replaces the selected pen with the pen specified by  hObject .    �  �    8   B� �&K!��!� ��� � �]  � ���  Selected objects are the default objects used by the GDI output functions to draw lines, fill interiors, write text, and clip output to specific areas of the device surface. Although a device context can have six selected objects (pen, brush, font, bitmap, region, and logical palette), no more than one object of any given type can be selected at one time.   Select-Object  does not select a logical palette; to select a logical palette, the application must use   SelectPalette .  *        *   '    � �&K!��!� ��   W       *   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description     �   W   #  F   ^� �&KR�тS~�!��� � �� � �� � �� � �� hDC   HDC   Identifies the device context.   hObject   HANDLE   Identifies the object to be selected. It may be any one of the following, and must have been created by using one o��5 �5 ��5 f the following functions:   �   �   #  �   C   X� �&KR���S~�!��� � �� � ���  � ��� Object   Function  Bitmap (Bitmaps can be selected for memory device contexts only, and for only one device context at a time.)   CreateBitmap    �   F   �   �   E   \� �&K���!���  � ���  � ���  � ���  CreateBitmapIndirect     CreateCompatibleBitmap    CreateDIBitmap   X       �   X   8   B� �&KR���S~�!��� ��  � ��� Brush   CreateBrushIndirect    �   @   X   �   E   \� �&K���!���  � ���  � ����  � ���  CreateHatchBrush     CreatePatternBrush    CreateSolidBrush   M      �   M   8   B� �&KR���S~�!��� ��  � ��� Font   CreateFont   H      M   H   1   4� �&K���!���  � ���  CreateFontIndirect   L      H   L   8   B� �&KR���S~�!��� ��  � ��� Pen   CreatePen    G      L   G   1   4� �&K���!���  � ���  CreatePenIndirect   P      G   P   8   B� �&KR���S~�!��� ��  � ��� Region   CombineRgn    �   u   P   �   Y   �� �&K���!���  � ���  � ���  � ���  � ���  � ���  CreateEllipticRgn     CreateEllipticRgnIndirect     CreatePolygonRgn     CreateRectRgn     CreateRectRgnIndirect   *      �   *   '    � �&K!��!� ��   �   �   *   �   3   8� �&KP!��~�!� � �� � �� Return Value  The return value identifies the object being replaced by the object specified by the  hObject  parameter. It is NULL if there is an error.    �   �     :   F� �&K!��!� �� � ���[  � ����  If the  hDC  parameter specifies a metafile, the return value is nonzero if the function is successful. Otherwise, it is zero.  If a region is being selected, the return is the same as for   SelectClipRgn .   W      c  <   J� �&KP!��~�!� � �� � ��  � ��� Comments  When you select a font, pen, or brush by using the  SelectObject  function, GDI allocates space for that object in its data segment. Because data-segment space is limited, you should use the   DeleteObject  function to delete each drawing object that you no longe��5 ��5 ��5 r need.    �   c    ,   *� �&K!��!� �������  Before deleting the last of the unneeded drawing objects, an application should select the original (default) object back into the device context.  An application cannot select a bitmap into more than one device context at any time.    7        7   !   W  \  ^  SelectPalette functionD      7   D   +   (� �&K �!� � � �� SelectPalette   [3.0]   �   K   D   �   E   \� �&KP!��~�!� � �� � � � � � � � �� Syntax   HPALETTE  SelectPalette( hDC ,  hPalette ,  bForceBackground )   j  6  �   j  4   :� �&K�!��!� � � � � �� This function selects the logical palette specified by the  hPalette  parameter as the selected palette object of the device context identified by the  hDC  parameter. The new palette becomes the palette object used by GDI to control colors displayed in the device context and replaces the previous palette.  *      j  *   '    � �&K!��!� ��   W       *   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   f  �  W   f  i   �� �&KR�тS~�!��� � �� � �� � �� � �  � ��� � �� � � � � � �� hDC   HDC   Identifies the device context.   hPalette   HPALETTE   Identifies the logical palette to be selected.   CreatePalette  creates a logical palette.   bForceBackground   BOOL   Specifies whether the logical palette is forced to be a background palette. If  bForceBackground  is nonzero, the selected palette is always a background palette, regardless of whether the window has input focus. If  bForceBackground  is zero, the logical palette is a foreground palette when the window has input focus.  *      f  *   '    � �&K!��!� ��   �   �   *   �   3   8� �&KP!��~�!� � �� � �� Return Value  The return value identifies the logical palette being replaced by the palette�ZHM�	��	�m�	��	��	��	 [� '����hz�@���+� ��� ������m������� � � � ��`
��
m��� �s����������`�,
� � 8� � 
�@@ 
�S�V}S�( �  �S����@d ��� �� ������ �󩠍  � � � � � � � � � � � �	�& ��"d#� ����/�O�o������멀� �`������_���`� ��@����'� ����0e�� e����`�


 Q��
e�� e�`d
&
&
&
&��
&e��e��@e�`H� |�hHJJJJ ��h)	0�:���H�Z�Z�Z ��z�z�z�h`8� d
&
&
&iN���e�� Z��
 ���� ��� ��0e�� e�z����8��~����`�"�NŅ�#�NŅ	F
�	F	*F	*L�F*F*F
�	F	*F	*L'�F*F*F
�	F	*F	*L:�F*F*F
�	F	*F	*LM�F*F*`        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l���  �U�`LX�� ;�� ��������������� ��L[�`dd� Z��� ��z���Z����� ��z�����`H ;���I���hdi��
&
&
&
&e��e�� �� ��������0����1����`����a�����������������	�����
����������� ����!����P����Q��`����`������`�$�%� 8�$H� �%�h`H�$E$�$�I�i�hI�i ��$$� 8�,H� �-�h`H���,
�-hJH��e-�-hf-f,��,�-`�%E)H$%� 8�$�$� �%�%$)� 8�(�(� �)�) 	�h� 8�,�,� �-�-� �.�.� �/�/`� �/�.�,���-F%f$��.e(�.�/e)�/f/f.f-f,��`````��8��
��i
�$�



$`�$�%��$�tǥ%�uǐ
�%�$�tǅ$8&,&-���,�-`    
  ( P d � � ���@�E�$��ǥ%��ǥ&��ǐ�&�$��ǅ$�%��ǅ%8&,&-&.����`        
    (  P  d  �  �   � � � @ '  N @� �8��@� 5```I�8i@�@�!���"

JJ(�I�i )?��C�(�I�i � `�� `����` 	"%(+.0369<?ADGILNQSUXZ\^`bdfhjlmoprsuvwxyz{||}~~`�)�(�JJJJ�)�
)


8�(�$�
)�J8�)�%�)


�&�)�J�'�e$f,8��jE,.�$e&8�(�,�,� �	e%f,8��jE,�%e'8�)�,�,�8``�|�$�5ɥ%�6ɥ&�7ɥ'�8ɐ�'�$�5Ʌ$�%�6Ʌ%�&�7Ʌ&8&,&-&.&/�����`            
      (   P   d   �   �     �  �  �  @  '   N  @�  �8 �� @ �  5 @B ��  	=  z ���  -1 Zb ������� ��8���I�i���8�	��I�i������������LZʰ0�Z� ��� y��e�8�����e��e � z���`Z� ��� y��e � 8�����e��e�z���`Z� ��� y��e � �e�z���`�"���H� Q��)��JJ����1�h=���` U��0����?```� �H�@�I��H����I�I�`�����[������d��������� � �˭����������i<���`

�� �˙ � �����`� �/ ������`������@�]�<��8�� !եHi0�J�Ii �K�������J�H���J�Hi0�J�K�Ii �K�������  �̭��a�1�]�-�D !բ���HȑH�� ��� �H�Hi0�H�Ii �I��ߩ��� ���_��a�Ș �ʭ��a�����`��`�����`���M�]�I��8�� !եHi�H�Ii �I�Hi0�J�Ii �K�������J�H���J�Hi0�J�K�Ii �K������� �̭��a�1�]�-�D !բ�ȱH��H��'��� �H�Hi0�H�Ii �I��ߩ�����a�����`��`



}�̅J���i �K�J��� !չ��eH�H�Ii �I��J�H��`�̽� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �ɍ& ���  ��� � � � � � �� � �( ����]�F�ЅG թ@�KdJ�� �J����K�K�`���� ��� �ӥ)������)�S� ��L�`ύ������gϘ �Ϭ �nύ�� ���uϘi ��� L|�@@@@@@8  0@P`8@@@@@@p�����Т ��	�8�������p���	�i������������i����ɀ�L�d�ɴ��  ����  ����`

��%Н�&Н�'Н�(Н����i������i��� ����`	
+,)*78'(56%&34#$12!"/0 -.                   P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������)��
�`�
�����0'� ���������Z v�z�����۠ ����������Z ^�z�����ة �`����������� !խJJeH�H�Ii �I��



eF�J�Gi �K�JJJJeK�K�)�	���J���J�	�
..
..���QH�HȭQH�HȭQH�H�Hi0�H�Ii �I�Ji�J�Ki �K��L��`e���`� ����`H)��<ՅHhJJJJ�I
eIi@}LՅI` 0`��� P���@p��      Hژ��\
�h�Ph�O`�k�l� �kH
���Ս�	��Ս�	� ����(	`l�	�բհբ �k� �����`� �k� �����`� �k�( ��������k`� �N�:	� �N��)�� �	�c	� �	��"�� � � �( ����`dN �բ!�c	�	���(�:	�N��` *֥N��`�(tN���!�	��L�՜	�W�X� � �W�O��������\� �Y�(	�	��_�`�a�N`�N�`�_��Lf����`��`�`� �_�am	�`�\�
�Y�	�Y�� LVؽ�ت�O�U�P�V�_� �U0L����L����L1����� �\����� �رU�am	�` ��L����� �رU�,	�U8�,	�U�V� �VL�����L8�����	�	�	}�ب�	�U�	�V ��L�����- �رUH �رUH�	}�ب�U�	�V�	�	�	h�Vh�UL�����' �ؤ_��ؠ �U�.	������Ui�U� eV�V�_L����� �رUHȱU�Vh�UL�����2��ع0	)��0	:�0	� �1	� ��U���٦_�YLJ� �� ��L������_���)��0	)�0	�0	�0	 �ئ_L��ɀ�(逼��

���ٙ.	��ٙ/	��ٙ0	��ٙ1	 �ئ_L�֤_�(	���ب�ٝ �Cٝ �0	� �1	�  �ؠ �U���٦_�Y �إ_
��U�O�V�P�_��(	��(	��`�^��[��[�LVؠ �S���� �^Lr���� �رS�8	�S8�8	�S�T� �TLu�

� �رS���م[ �ؽwٍ( �xٍ) �y�)�* 	�* LV�   �U��V`�S��T`H���,	
�-	hJH��m-	�-	hn-	n,	��-	�,	`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   �٨�1���  <�m�0((� 0 ('(0((� 0 (&(0((� 0 ('(0((� 0 (&0000 0 0�((((0((((0��  $0 �m�0 00#000!00	0!00	00#000#000#000!00	00!0	0!000#0�                              ���x����  60000000000000000000000000000000000��  "00000000000    	000    0 	  	 0 	  	 0	  	  
0	  	  00    0  00� ��^ݒ���  80 0 00*00000 0 00*0��  $	000%0	00	000%�            ����#���  :
�  �  0 0 ���  &			0	 0 	������	m�	��	M�	��	��	��	.�	M�	��	m  M  e`�	���ȑ����� ��i0��i ���L��`��ȱ����	��� ��i0��i ���L��`��Hȱ����	��h��i0��i ���L��`�	����
0�������8�0��� ����L�ޤ
� ���	����`�	����
0�������i0��i ����L1ߤ
� ���	����`��	���
�������	`��'�����0e�� e��0e�� e���` PAUSE  `

����	� �
��7����BɎ��d

&$
0%��	���	���	���	����i�f
L��Ȟ�	��	��	��	L�ߥ	��m�	�f
L��``H)��4��uhJJJJ�v
evi@}D��v` 0`��� P���@p��      ```����`��� � �Z��ٝ	���ٞ	���ٟ	���٠	�L��)������	����	����	����	Z ��z��	����	����	����	����	)�	� ��z������Љ`��	��	��	��	��	��	��	��	��	)i��	��	)Ji��	�0�~d��	��	m�	:H���E~�~h ଡ଼	JJeu�u�vi �v��	�



ey�m�zi �n��	J�jJJJen�n��	)��	��	� ��	,�	p��m��	��0�� �mڪ������	��	�!�	.�	.�	.�	.�	�	.�	.�	.�	.�	��߬�	��	Qu�u���ue~�u�ve�v�mm�	�m�ni �nΓ	�Lg�` @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��d�������� ������o�����������������������������������������o������d���������d�d�d����[�\�]�^�Y�Z� ������	`����P���_��� 鹩c�
�P�������������������O������������2������o��M� ��)���5������d��������`�	���	���"� �#�	��� ;��  ��`�	��&� �"��#�	��� ;��  ���	������"� �#` 7Ǎ)��
���� ��NNNN���������� ��
��������� ��`
����������������������S�T�U�V�W�X�Y�Z�[�\���ȝp���4�H�\�� ���`� ڎ � Z������`��! ��]�!��5�H�d	
&	
&	
&	
&	��	�

&
e��
e		@�	hH F�hHJJ�h)��V�Q�`0���qd	
&	
&	��I8��I�5�	�5�  Z�)�p�)?i �]���5 Z�)i�q`���p�4�\�� ���`� ڎ �� -������`��! ���]�!��5�H�d	
&	
&	
&	
&	��	�

&
e��
e		@�	hHJJ�h)��)�Q��0e���	�)�Q�`8��q}]�]ɠ� Z�)i�5�] Z�)�q`�	�& ��"� �#�J�y�w���z�x���	��� ��	�������������0�������ɠ� �L��H�e�� e������h��J���� zũP�� �2 �� �歆�L��)�& L�Ά� ��@�� JJ����PJJ�	 �ީ ��@��PJJ�����JJ�	 ��`��  B筇����� 5�LW੩���� L��
��[��\���ȱ��I���`_�q��	
 ���	�& �J�y�w���z�x���	��� ��	����� ��������8�V�H�e�� e������h� @��� ��@�� JJ����OJJ�	 �ީ ��@��PJJ�����JJ�	 ����`Ί������
��[��\�� � �� W��H�e�� e������h�L��^�' �]�& �\�% �[�$  �ȩ�"� �#���	������ Sũ��� ;��/ �.  v����� ;��- �,  v��� ��`******************  TOTAL SCORE  **_______________**               ****************** �  I���H�e�� e������h����  I���`�ŉ�`��� �饈)�	 �� D�L��`��h��d��i8�� �W��i8���J�o������� X������
�������l    ����饅�
��`��`L䥄���`���o` Z��d�)?i!��)����������`���ƋƋ`�o��`���o�	�

���	`��������
������� ��`#�'�)�#�)�#�'�)�%�'�<�=�>�?� iߥŠ�`��汥�Ţ�d� iꥨ |� �� � �� �� s� �� �� 2� ���`�����������������)�����`����������������������)`�����`����o�������� Z�)��8���d�Lm�` ��L-��1��-����������	��
���������  �Ȑ��d�`"""""""����������� I���`�8��� �8����o��������d�� X�Lc�`��

i�����������
��������� ��`�o�`����7����}����}��������
��E���F���� ���`�o��`                        ��ɭ���� ����"�`権���`pppp���������������W��`��Ţ��`��9b���������`          
��������)�*�+�,�-�.�/l ������������7�b������d�d��������`��������`��������`��������`��������`���������������������`(<Pdx��������������2����������`�������������]����������`��������������������������`Fn(Z����   �������	����������������`������ v v v�������
�������������`������ v v v�����`��
��!��"�l      L�L�L�L�L�L�L�7�L�g�L�d�`���F`����榐ƦƦ����槐ƧƧ`���n�`���v`��
�������l `�������)�W�����索


 �ɀjɀjiF��ƦƦƦ�`檥�

 �ɀjɀje�i2����


 �ɀjiP��`檥�

 � �ɀjiK����i!��`檥�

 �ɀjɀje�i#����

 �ɀjiS��`檥�
e� � �ɀjiP����
 � �ɀjɀje�i!��`��!�)�/���������8���`��i��`��8���`�����}���}�` ���  ��� �檥�


 �ɀjɀjix8媅���
 �ɀjɀjiP��`������`�)�`桥�)i��`        �!�'�-�3�5�7�9�;�=�?�A�;�A�C�=��� ����HI� R��&�(�(�&�'�(�)�*�]�S�U�W�Y�[�]�7�8�9�:�;�  �  ��% �) ������$ ����(  	ǭ, m[�[�- m\�\�. m]�]�/ m^�^�^�' �]�& �\�% �[�$  �ȩ�"� �#��� � ;��/ �.  v��
�� � ;��- �,  v�`
 �� E� �� c�L񦥽M�A���L&�C������i&��5��A���L��9� ����M�58���5`�o�M���5`���M0`�5��A���������� ����`�8����8����������o�����M`����#�M��8�5����8�A�����o�M`��0` Z�)ť�� ��M�o�`���M���5���A`xآ�� ����� ��	����� � �ʩ��	 � � �Ω)�& ��"� �#  � ���  m� ֩	�&  ���y�w���z�x t㍽� ��	����� �䭋� 0����� ;�����	��  ���L���"� �#� �� ����� S� �� ����� *֭�0�o����� V�憥���d�LK��0*�	�� 퀥N� z�N��L0� ���������  X��
�(�A���3�)�"I�#���
������ Sť����� � �� �� ���d� ��L��毥�)�2�0��C�� JJ����JJ�	 �ީ ��[�� JJ����JJ�	 �ީ�� +����������  )��v �թ` Q������� Q� |ߩ �"��#��������߅ Sŭ  )����H�e�� e������h��  )����  )��� �թ� Q������` Q� |� ]� ��  � @� &� W� ��L��Ŭ�`��步�)?��
��
LQ�`�`�`�a)�`�� ��΄ ���ƅ���
�����`�`��a��b��c`� ��C����0� ����0e�� e����`� � ��	����(���0� ��	�������` DANGER           SCORE:        POWER: ��������  X��
�(�A���3�)�"I�#���
������ Sť����� � �� �� ���d� ��L��毥�)�2�0��C�� JJ����JJ�	 �ީ ��[�� JJ����JJ�	 �ީ�� +����������  )��v �թ` Q������� Q� |ߩ �"��#��������߅ Sŭ  )����H�e�� e������ by the  wMSeconds  parameter. The caret flashes on or off each  wMSeconds  milliseconds. This means one complete flash (on-off-on) takes 2 x  wMSeconds  milliseconds.   W       �   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   ~   F   W   ~   8   B� �&KR�тS~�!��� � �� � �� wMSeconds   WORD   Specifies the new blink rate (in milliseconds).   *      ~   *   '    � �&K!��!� ��   C      *   C   -   ,� �&KP!��~�!� � ��� Return Value  None.  *      C   *   '    � �&K!��!� ��   �   �   *     -   ,� �&KP!��~�!� � ��� Comments  The caret is a shared resource. A window should set the caret blink rate only if it owns the caret. It should 0'6 Z'6 �#6 restore the previous rate before it loses the input focus or becomes inactive.  ,        ,   (   "� �&K!��!� ���    5      ,   5   !   �  g  i  SetCaretPos function7      5   7   (   "� �&K �!� � �� SetCaretPos   g   (   7   g   ?   P� �&KP!��~�!� � �� � � � � � �� Syntax   void  SetCaretPos( X ,  Y )   h  4  g   h  4   :� �&K�!��!� � � � � �� This function moves the caret to the position given by logical coordinates specified by the  X  and  Y  parameters. Logical coordinates are relative to the client area of the window that owns them and are affected by the window's mapping mode, so the exact position in pixels depends on this mapping mode.  �   �   h  �   5   <� �&K!��!� �� � � � ���  The  SetCaretPos  function moves the caret only if it is owned by a window in the current task.  SetCaretPos  moves the caret whether or not the caret is hidden.   W       �   W   7   @� �&KPтS~�!��� � �� � �� Parameter   Type/Description   �   �   W   �   R   v� �&KR�тS~�!��� � �� � � � �� � �� � � � �� X   int   Specifies the new  x -coordinate (in logical coordinates) of the caret.   Y   int   Specifies the new  y -coordinate (in logical coordinates) of the caret.   *      �   *   '    � �&K!��!� ��   C      *   C   -   ,� �&KP!��~�!� �  TP     BAT           �K�Ma�    TP     BAT           �K�Ma�    TP     BAT           �K�Ma�                                                                                                                                                                                                                                                                                                                                                                                                                              ���