wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwxww�wx�w�w�w�x�wwww�w�wx�w�wx�ww�w��w�wxwx�wxww�x�x�w�wx�x�x�w�wwww�w�wx�w�wwxwwww�ww�w�w�w�w�wxwx�wx�x�wx�x�w�wx�w��x�x�w�x�w��x�xwxwx�wx�w�w��wx�w��x�h��h�f�w�ww�wx�w�w�vx�w�w�wx�w��w�w�ww�w�x��wxw�x�wwwwxw�w��x�w�x�h�w�w��g�wx�w�wwxww�wx��w��g��w��w��wx�xwx�w��xw��w�w�x�w�v��x�w�w�w���x�wx�g��h�g�g�v�w�w�g�w��h�fx�h��g�g�f�wx��x�f��w��w�fwx�x��x�h�vx�g�g�g�xw�vx��xw�w��vy�w�w�w�h�g�f�g�W�x�g�g�h���wx�w�xwx�w�g�v��h�ww�h�g�w�f��h�g�g�vx�f�vx�v�vx�w�vh�uy�h�h�h�x�h�f�w�wxxw�g�w�w�ww�ww�w�vx�x�g�v�xwwx�g�f��f�g�vx�e��h�h�x�hw�h�h�hv�f�f��wx�w��h�V�uh�V��Y�W�vx�x�xw��g�f�v��h�h�xw��w�g�w�w�g�g�g�g�g��w�f�v�x�g�w�w�vy�w�vx�h�v�wg�v�uywwwx�g�fx�wx��g�g�g��h�x��w�x�x�X�fx�f�w��x�wx�g�vx��h�xx��g��h�e�v�vh�V�ui�Y�G�F�vx�vy�X�W�g�v��w�xwxw��g�f�f�g�wx�wx�v�v���wwx�g��wx�wx�w���w�w�w��x�w�wx�x�ww�w�w�ww�wx�ww�wx�w��ww�wwwwwx�����x��wvgeVwwx������wfeDUUfx���˩��vUDD35Vg����˩�vTCC"4Vx�˼�̺�vT""Ex�ݽ��˩�U0 Fy�����ʘvC! Eg������eT225x�������d4B2 5CDW������ɆB4#1eEUx�����ڇS#3CfUfg�����ۇSCD"WffV�����̗d4EBGvvex��﷭�u!$ESFvgeW���ƌ�u1$Fd6�weVz���|�v1FuF�xuEh���j�wAE�E�x�DW���YɈQ5�V�x�DE���W��s $�fwh�d4|��e���z��g�u2I���y��AI��fx�C5���X��c ���gxd3j��v�y� j��UgvCF���wV�R &�܆UVd4k���dhu i��uEUDF��ږEwS%�ݨdDTD{���dVe2X�ۖC4DW���EeT"5zݺt24E{���tEUC#W�ܨC"4W����DTD25i�˅25{����EDC#V�ܹS#X���DTD3Ez�˄!F����dED34h�ܦ1 %����tEDC3W�ܷA ����c5UD3F�ݸA ����B5UTDF�ݷ0 '����4geDG�˕[���P5�vTX��c ���� X��Vw�uCG����  &���eUUV����sF���eD4h����1 W��uTDX����RFx�vUUh����cFx�vUUh����d!EgwfVg�����uC#DVffgx���˩vTDEVgww������wwwwwwwwwwwwww����wwwwwwwx������wwwwwwwwx����wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwvffwwffgeVx�������������fg����������wwwwwwwwwwwwwwwwwwwwwwwwwwx����������x�wwww�������wwfffffw�������vUTEUVfw����˨vC"#Eg�������u1  F��������u! #W��������S 4h��������B#Eg��������  4Vx�������R 4Vg��������  Efx�������Q  5gx���x����  h���������@ G�����w���� x�xx�vx����  7��ww�fx����  7��wgwfx����  7���fveW����  ���vwfUy���` X���gveV����  ���vwfTF����  %���v�eCF����  6���w�eC6����  %���w�uB$���� z�����C#Y���P X�����S!&����  %��x��u1Z���P X�����S����  %��x���BH���� G��x��d |���  h�w���B6����  5��g���2j���` W�vwx�e26���� x�gfxvUEz���r F��vVwfUh����! W�vefffh����c!EwveUfgx���ܦT3EgwfUUfw�����wfw���vUffgwx���ww����wwwwwwwwwwwx����wwwwwwwwww����wwwwwwwww������wwwwwwww�����wwwwwwww�����wwwwwwww�����wwwwwwwwx����wwwwwwwwx����wwwwwwwwx����wwwwwwwwx����wwwwwwwwx����wwwwwwww����wwwwwwwwwx���wwwwwwwwww���wwwwwwwww���wwwwwwwwwx���wwwwwwwwwwx�wwwwwwwwwx���wwwwwwwwwx��wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww�wx��x�wwww���wwwwwwwwwwwwwwwwwwwww�www���wwwwwwwwwx��wwwwwwwwx����wwx�wwwx����ww��wwww����wwx��wwfffh���wx���wvfTVh���x���vg�eT4Vy�ܘ���vTWvT24W�������C"UDC#Vg������s U4TE�w������b v3VW�e[��g��r &�"Gw�Dk��W��RFuX�eE���i�BDSi�Ef���y��C"DCztFx�����C#3CydVw���z��C#C3$�SWw���|�uC$22%�Chx����TC4"27t5�������D3A#gSX������TC3"6d6����y��4304fDy������4C1#VSH������CDB#ETF����l�s4C5T5����z��ED4TE�������5D 4TDy������4T04TDh������4T04D4h������4TA4D4h������4TA4C4h������DUA4C4g������ET0325g������EU03"4W������VT2Eh������fB Ex�����fe0 3F������fS  4h������u    F�����ɇB   $j������d   X������u1   G������A   G������t!   X������S   F������e1  6������vd!3F���̻�weDDUg������fefw����wfeUW������DT"Fx������TC4Vx�����vUDUg������vUfg�����vfUVy�����fUDV������eUDW������feVx�����ffUg�����wfUVx�����wfUgx�����vffw�����wvfw�����wvwfwx����wwwwx����wwwwx�����www�����w�wwx�x��x�w�w�w��x��������x�w��x���w�ww�wx�x��x�������w�ww��x��w�g�wgwww�wvxvg�f�wx�f�vg�g�vy�y�y�xx�W��w�f��gwwxuhu�fxvxvh�g�h�vx��W��x����X�g���vy�Z�7�W�v��X�X�X�F�Ux�f�v�vx�g�vx�h�x�h��f�X�i���z�Y�x�vz�{�I�Y�Y�X�Y�W�ti�W�e�ez�I�G�uj�i�h�f�e�uyw�w�uz�h�f�u�uyv�d��g�g�W�E�u��{�i�v�vy�x��vx��w��xw�h�G�D��Y�8�G�wx�W�e�tk�y�y�i�i�i�Y�X�i�xxvx�g�V�w�i�[�m�k�i�g�f�e�wg�f�g��x��vy�g�T�E�V��g�vx�g�gx�X�F�E�uy�h�e�uz�J�X�X�i�j�i�w�i�X�vi�y�i�fx�F�U�v��f�e��X�8�X�W�d�e�v�e�C�E�V�ez�i�k�{�x�wx�f�U�tj�h�ty�xv��v�V�X�h�e�u�w�x��uxfh�Y�H�H�i�x�u�d�e�tz�ze�e�V�W�w�W�g�u�d��w�hu{�Z�k�[�F�f��z�j�x�x��W�g�Y�j�y�Z�9�Y�hwxy��wxw��w�u�uy�k�I�Y�8�g�h�V�G�W�u�vyv�f���wx�f�vx�xx�xv�ui�f�w�X�w��X�X�w�f��X�vxx�wx�g�x�h��y�i�i�wx�h�x�w�vxw�ww�g�h�h�xv��xw�w�x�x��w�wwvx�h�h�w��w�vxvgvh�x�����vVUUUx������eT2#4Vh����˗e2#5y����ܩt!  $h������u    W������v0   F������uB  #Y������!!  T5������s  Fwv����I�C@dW��wx���%�et�Ug�uD4g����ȇ6S4W�DUW���V�vr WUV{�r5T4j��lۙ0fTE��S4TE������ fei��14\���� EUX���"  ����ʀ Vf���P   ����P W����@   	���ޔ   Y����P   ����   :�����   ����a   �����   �����    >����    ������    ����@   �����   ����    
�����   U����    ,�����   �#����    �����@  �R���    ������  M�[���    ������  �X���    ��ڿ��  �v����   [������  ��|���   G������  
�����@  V��ʜ��P  �ɜ���   Gz�ܙ���  	�����@  ������  n����   Y��˘���   �ڽ���  ��ܩ����  �����`  ��ʘ����  
�����   )�ܹ�����  �����   )�ܹ�z���  �����  9�ܨw����  	�����   �ݹ�y���  �����p  ��ʇg����  \�����   Z�˘vz���  �����p  �ܹ�V����  �����   8�˘vg����  �����  I�ʈvh����  �����  Y��x�g����  �����P  8��vff����   ~�����  �ܖffh����  �����@  9��eff����`  L�����   �ݧUgw����0  n�����  ��Dgx����@  n�����  ��EWw�����  *�����   |��TVwx����  �����P  ��dV�w����   �����  ��Ex�x����  �����@  ;��TExwy���P  L�����   ���DX�fz���  ������  ���4W�f����  ������  ���EgfV����  ������  ���Ex�U{���  ������  ��Egvez���0  L�����   }�Tg�eh����  �����0  :��dVfeV����  ������  ���DhvUi���@  ;�����  [ݸfh�TV����  ������  �ۆVxvUi���p  �����0  )޸vg�TE����  J�����   j̨w��DF����   l�����  �̗wxuDG����  {�����  �ˈ���CG����  ������  �����u3W����  z�����  y����u3G����  Z�����   X�����C5����0  �����   &�����C$j����  �����`  h�y��t3X���� h�����  Fwh���26����b  �����P  Ww�̹d#W����0  'h����  Vg�ݸS$h����  Vi����  #Di�ۖCEy����  ej����  4X��CEy����0 TX����    i��TEx����@ U6����   5��eUg����S 53z���Q   {�ʆffh���� %Q&����    &�۩vwfi���T E7���t2#  J̺���U|���B DR X���TDT  j�����U����BUPX���ffd  X�����V����TU@ X�����u  FVh�˗f����VBEB &��ʙ��@  3F���������s$Ch�몫��   X���������RE3 Xͺ����!   V���������cD2 G������C! 5h�x�����˦fT5��w���UC33"4Vwwx�����ډ�R"FeUWy�wffUC4DUUVx�����˻�eTDT33DVfffwwwfffffw���˫�̺���weTDDDDDEUUUUVfgx�������ܻ��vTDC3333DDDUVfwx�������ܻ��vTD33233DDDUVfgw��������˻��eDD33#3DDDEUffgx��������˺��eDD33#DDEDUUffgx��������˺��eDD333DDEDUUffgw��������˺��eDD333DDEUUUffgw��������̻��vTDD334DEUUUVffwx�������̻���eTDDC4DEUUUVfffwx�������̻��veUDDC4DUUUUVffww��������˻��vUUDDCDDUUUUVffww��������˺��veUDDCDDUUUUVfffww�������̻���eUTDC4DUeUUffffwwx������̻���fUTDD4DUfUUffffgww���̼��˺��veUUTDDEVeUVffffwwx������̻���fUUUTDEUfVUffffgww���̻̼˺���fUUUDDUVfVfffffwww���̻̼˪���eUUUDDUVeVfffffwww���̻̻�����fUUUDDUVeVffvfwwww������˻����fUUUDDUVeVffffwwww������˻����veUUTDUUfVffffwwww����˼̻����veUUTDUUfUffffwwwwx���̻̻����wfUUTDEUVUffffgwwwx������˻���wfUUEDDUUeVfffgwwww����˻˻����veUTDDUUUUffffwwww������̻����wfUUEDEUVeffffgwwwx����˻˻����vfUTTDUUfVffffwwwwx�����������wveUUTDUUfVffwwwwww������������wvfUUTDUUffffwwwwww�������������vfUUUDUUffffwwwwwwx������������wfeUUTEUVfffgwwwwww�������������vfUUUDUUffffwwwwwwx������������wveUUUEUUffffwwwwww�������������wfeUUUUUVfffgwwwwww�������������wfeUUUUUVfffgwwwwww�������������wfeUUUUUffffgwwwwwx�������������wfeUUUUUffffgwwwwwx�������������wfeUUUUUffffgwwwwwx�������������wffeUUUUffffgwwwwwx�������������wffeUUUUffffwwwwwwx�������������wvffUUUUfffggwwwwww��������������wffUUUUUffffwwwwwwx�������������wvffUUUVffffgwwwwww��������������wvffUUUffffwwwwww�x��������������wvfffeUffffwwwwww�x��������������wffffeVfffgwwwwww�x��������������wvfffeVfffgwwwwww�x��������������wwfffffffffwwwwwwx����������������wvfffffffwwwwwwww�x���������������wvfffffffwwwwwww��x���������������wvffffffgwwwwwww��x���������������wvfffffffwwwwwww��x���������������wwfffffffwwwwwww�������������������wvfffffffwwwwww�x�x���������������wwvffffffgwwwwwx�������������������wwvfffffgwwwwwx��������������������wwffffffgwwwwwx��������������������wwvfffffgwwwwwx��������������������wwwfffffwwwwwwx���������������������wwvfffffwwwwww���������������������wwwwffffwwwwwww���������������������wwwvffffwwwwwww���������������������wwwwffffwwwwwww���������������������wwwwvffgwwwwwww����������������������wwwwffgwwwwwww����������������������wwwwwwgwwwwwwwx���������������������wwwwwwwwwwwwwwx����������������������wwwwwwwwwwwwww����������������������wwwwwwwwwwwwwww����������������������wwwwwwwwwwwwwwx����������������������wwwwwwwwwwwwwwx����������������������wwwwwwwwwwwwww�����������������������wwwwwwwwwwwwww�����������������������wwwwwwwwwwwwwwx�����������������������wwwwwwwwwwwwww������������������������wwwwwwwwwwwwwx������������������������wwwwwwwwwwwwwx����������www�����������wwwwwwwwwwwwww����������wwww�����������wwwwwwwwwwwwww����������wwwwwx����������wwwwwwwwwwwwww����������wwwwww�����������wwwwwwwwwwwwwx����������wwwwww�����������wwwwwwwwwwwwww�����������wwwwwx�����������wwwwwwwwwwwwwx�����������wwwwwx�����������wwwwwwwwwwwwwx�����������wwwwwx�����������wwwwwwwwwwwww������������wwwww������������wwwwwwwwwwwww������������wwwwww�����������wwwwwwwwwwwwwx�����������wwwwww������������wwwwwwwwwwwwx������������wwwwwx������������wwwwwwwwwwww�������������wwww�������������wwwwwwwwwwww��������������www��������������wwwwwwwwwwx�������������������������������wwwwwwwwwwx������������������������������wwwwwwwwwwx�������������������������������wwwwwwwwwwx�������������������������������wwwwwwwwwwx��������������������������������wwwwwwwwwx���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU=|UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�\�����������������������������������\�����������������������������������VUUU�����_=   |����_VUUU�   p   �   ������������        �:        �:        �:        �:        �:        �:        �:        ��        �����������ZYYY����������������ݶݪ����ݶ������ݶ������ݶ������ݶږ����ݶڶ����ݶݖ����۶��z�y�~�zww�����zww�����zww����yw�w����yw�w����yw�w������~���*X%X%Z�V�X%`	�P��V��@�V��u��}��u��v��v��v��v��u�����U��U�j��jW�je��Z��֥�u�j]�jW�j��jU��U�j��jW�je��U�����U�je�jW�j���U��Z��֩�������ݩjݩjשjץj��jե�Z�  ��         0         ��        ��#     ���>�Z  h�����Oݪ�U[PUU ЫVU�T)@��@�S� %�eU}��S� ��~��ݼ�S�  @�U����S�   h�����S�  @�W����S�  @����?S�   d @��P� U   �?TU�UU    PUD��U       �W        `�~        @���<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�                   �    0   ��  pu  \}5  \U�  U�  T�  WU�  [U�  l�:  ��  ��                                      �   p?   ��   ��  p�  _� ��_�p�~���W� �_�:  ��  ��                                  �    0    �   �u  �U  �A  pU:  pE:  \Q�  \Q�  lU�  lU�  ��:  ��:   �                           �   �=   �� �Zo ���? �u�� �����^����� ���  ��?  ��� ���  �   �                                �   �}   �   �   �   \   �  ��  p�  p�  ��?  ��   �   �   �                            T    �    �    �<  �?�  ��  � |W ��� �� 嵧�鹯����  ?                                      ��  ��: ���� ���� ���� ���� ����  ��:  ��:  ��  ��  ��    ?                                  3   ��  <3  <3   <3   <3   ��   3   3   3  <3  ��   3                              �    0   ,   +  �.  �+  �.  �
 ���  ���  ���  ��2 ���0 �* � �?�   �                                      ��  �P?  K�� �`������fЪ�������  ��>  ��                          ������������\�\�����P���{� 0�?��.\  �,��pppppp?z;z;�4 0d6�:�:�?�?�:�:d6 0�4z;z;?pppppp�,��UwUuUuU]UWUUUuUuU]UuUuUUUWUWUUuUuUUUuUuU]U]U]U]U�_�]�]�]�]�]�_�_�]W]W]WW�U�_�]�]�]�]�_W]W]�_�U�U�_�]�]�_��������u�]�����������u�]�����]�]�����������������������  W�����������������������������������   ������������������������������������V  p媪�������������������������ZUU����[  \�����������������������������������n5  W����������������������������  ������ ��������������������������������������Vp嫪����������������������������������[\�������������������������������������o5W�������������������������������������j�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�[UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����������������������������������������>�������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU �������������������������������������� ������������������������������������������������������������������������������������������������������������UUUUUUUUUU]UuU�UUU��U�W�_UU���V^[yUUu�ו^WzUU���f^�yUU��ת^�zUU��U�W�_UUUUUUUUUUUUUUUUUUUU�U�U�WUUu�սW�^UU]�w��UzUU]�w�ޕzUUu�թW�^UU�U�U�WUUUUUUUUUUUUUUUUUUUUUVUYUeUUU�_UU�UUU�y��U�WUU}����w_UU}�����~UU���w_�}UU��U�W�_UUUW�]�wUUU�UUWU]UUU�U�W�_UUU�UuW�]UUU�U�W�_UU�{U�U�WUU�vU�UmWUU�}����WUU�_u��UUU�U�W�_UUUUUUUUUUUUU]UuU�UUWUU�U�W�_�yU�U�Wu^��U�W�_u~u�ՕWW^]y���VW[]muu�եW�^]z�U�U�W�_UUUUUUUUUUUUUUUUUU�}��U�W}_�굪ת^�z�굪ת^�z�굪ת^�z�z��U�W�^�^U{U�U�WUWU]UuU�UUUUUUUUUUUU�U�W�_U�U�W�^U{UgW�]uv���y��]�w}�]�wy��y����՟W^�y]yu�ՕWW^�_�U�U�WUUUUUUUUUUU]U]U]U]UU_U_U_U_U�^�^�^�^U�^�^�^�^U�W�W�W�WUkWkWkWkW��������U����UUUUUUUUUUUUUUUUUUUUUUUUUUUU����uUUuwwuw]wUUuuwuw]WUUuuwuw]WUUu��ww]UUuuwuw]uUUuwwuw]u]Uuwwuw]wUU�w��u]]UUUUUUUUUUUUUUUUUUUU]���]UUUU]]�]]UUUU]]�]]UUUU]]�]]UUUU]���]UUUU]]�]]UUUU]]�]]uUUU]]�]]UUUU��u��uUUUUUUUUUUUUUUUUUUUUUUUUUU]UUU��UUU��WUUu�WUU��WUU��WUU��UUUUUUUUUYUUUUUUU��UUU��WUU��_UU�w_UUU�WUUU�]UUUUWUUU�WUUUuWUUU�WUUU�UUUU�UUU��UUUuUUU�WUUUUUUUUUUUUUU]UuU��U�W���V^u�ו^���f^��ת^��U�WUUUUUU�WUUUuWUUU�WUUU�UUUU�UUU��UUUuUUU�WUUUUUUUUUuUUUU�UUUU�UUUU�WUUՕWUU�VWUUեWUUU�UUUUUUUUU�UUUU�WUUU�]UU��]UUuy^UU՟WUUu�UUU�UUUUUUUUUUUUUU]UuU��U�W���V^u�ו^���f^��ת^��U�WUUUUUUYUUUUUUU��UUU��WUU��_UU�w_UUU�WUUU�]UUUUWUUUUUUUUuUUUU�WUUUwUUUU�WUUUuWUUU�WUUUuUUUUUUUUUuU�UU�U�WU�U�WU�W�_ՕWW^�VW[]եW�^U�U�WUUUUUU�U�UU�W�WU�]�]����]uy~y^՟ןWu�u�U��UUUUUUUUUU��z��z������������wz�zwwwwzw�zzww�zw�zzwwzw�zzwwzzw�zwwwwzw���wwzw��?��? � ��  � ��  ��� � ��  � ��  ��?0�?�       < <��?<����� < <�<�<<0030 < <�< <0030 < <�< ��3030 < <�< � 3030 < <�< �3030 < <�< <3030 < <�<�<<���� ���?�?<�                                                                                                                                                                                                                                 �    ��        �      ��0<� �0��   �0�0��?�0  30?�� �0<  �00�� �<�  ��� 3?                 �3  � 0� �?  0   �3� 0   �3����0 3??�0� �3� �3� � 30���3� 0 3� 300� 3� 0 30���3���00 ���               �     �� �   �  �   �0  �   � �� ����   � � ��3�   �� ���0�   � � 0�0�0�   � �� ����0�   �0      0     3����3��0�03�0����3�0� 3 03���           �3  0      0  0      0���     �0�0     0��0     0� 3     0��0                �3  � 0�   0   �3�   �3����  �0� �3�    30���3�    300� 3�   ��3���0  �  <   3           �      � �  303�    0�? 0 0�    0 ? 30�   0�0 �0�   �� ? 3��                   �  �?          �   ��          ���<�<       ���0�?��       ���0� ��        ���0� ��        �0� ��                        � 0     � ��   �  0     ��   ����?�������� 30� 0��0��0���3�0� ����� �3000� 3��0� <��3��� ����       ?   ? ?       ?   ��  ����   ?   ��   �� ���� ��   ��  �� ���� ��  ��  �� ����? ��  ��?  �� ����? ��? ����  �� ����?���� ������������?���������?�����?��������?�??�?����������������?��������?��������?��������?���� ����?���� ����? ��? �??� ��? ����? �� �?� �� �??� ��   ?   �� �?� ��   ��   ��  ����  ?   ��   ?   ��       ��?      ��  0  0  �  �� 0  0  �  �  �  � � ��? �  � �0< � � ��0<��� � ��3����� � �3�������������?��?�0<��������?��?����������3��3���������������?��?����0<��?��������?�����3� � ���������� � ��0< � �����3� � �  �  �  � � ��?�0< �  0  0  � �  0 � �  0    ��<   ��� ����<��?�?0303���?�?�������������������?�?0303�?�����?�� ����<��  �  �<  ����������������������������MQEQ�  �3��5��WQEU� O�GQ�  �<3��� _@�� \A5� �  ;�̬�� |QE� � �UUU5� ���?�^� ����? � ����7�0���~� �   �    �� �: ��z�  ��� �  ���U�0�> 0�z�  7 �  �  pU�������?�z�  7?�  � �pU��0���z�  7 �  � ��pU?� ������  7�  � <0�U �0� ���  7 �  �  �U ��� ��� ?7��  � ��U��� �< ��� �7 �  � � �Us�� �  ;�� W5��  � �?�U����?����� W5 �  � � �UU����� ��� ���� � � wUU��������O������ � �����������_������� ��������L������?� �����������\��������� ��������ë��� \�|����>������� ���30� O�\=�����������> ����<<<�\�\�ë�������������0\�\U��������������?0L�\U��������*�������?p������_=�������>���ëì�0������\����Wլ«������0�����������W��#����:������:������_���������<00���?����>����������� <��𺺺���������� ��� ���?������������< ���� ��������� �� ���� ����������������� WUu ��������������<�� WU} ��߫> ���������� �W�� �������  pU�� 7W=  ��� ��� pU�� ?W= � �|����� �  p��  W= � �\�� ����� p���  W=0� �\����:0� p ���W5�< �|����: � <�s ��|W5  �|���0� p ��_W5  �̵������ ��s ��W���� ���0 �0�  p ���    ��:� � � ��� ��p���� ��:���0��   ���sUUU= ������ ������? �� \p�� �\��� � |QE� � ES��|�3� � _@���EQ��p��3� ��WQEU����������������������������0 ��������������    ((((�*�*((((�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������?� � �?� ��? ��� 0<�� ? �00000�00��? 00 � 0 00� 00  000000� <�3 �000�00�0000000  0 ��?�0 0 00  0000000 0�3 � 00030 300�? 0  � 0�0 00 ��?�  ���?�0�3 � 0000�  <0000 �  0 �?� 0�?00 0�  0000 0000�3 � 03000 3�?00 0 00�  �00 000 � � 0000 000��0� 0000�00000� 00��? � ��?��� �?�����<�0���3�000000��?��
�
����
�
�*� �  
(�(����
((�� �  
((����� 
((�� � ��
(����* �
(�� � �
(������ �(�� �  
((������
(�� � ��
(�����

*�*��������*�
��� ��  �� ��  �� �
�*� �� �   ���   �� ��� �����
  *"   "   
�   ""    "�"    " �
� �*"������������?�  �  �  �  00    <0    <0    300� 0� 0� 0�000� 0� 0� 0�00�0 �0 �0 �000       00       00       00�0 �0 �0 �000�0 �0 �0 �0000� 0� 0� 0�00    30    30    <�  �  �  �  0�  �  �  �  00    <0    <0    300� 0� 0� 0�000� 0� 0� 0�00�0 �0 �0 �000       00       00       00�0 �0 �0 �000�0 �0 �0 �0000� 0� 0� 0�00    30    30    <�  �  �  �  0�  �  �  �  00    <0    <0    300� 0� 0� 0�000� 0� 0� 0�00�0 �0 �0 �000       00       00       00�0 �0 �0 �000�0 �0 �0 �0000� 0� 0� 0�00    30    30    <�  �  �  �  0�  �  �  �  00    <0    <0    300� 0� 0� 0�000� 0� 0� 0�00�0 �0 �0 �000       00       00       00�0 �0 �0 �000�0 �0 �0 �0000� 0� 0� 0�00    30    30    <�  �  �  �  0������������?  �? �? �? ?�? ?�?���?���? 0�? 0�?���?  �� �� ���������� 0�� 0�� <�� <��� ��  ��� �� ��� ��� ���� �� ��� 3�� 3����?��   �� ���  �� 0��� 0 �� 0��� 0 ���0����0 �� ����   �� <��  �� <��  �� �<�� � ����<���� �� �<��  �� �� �� �� ���������� 0�� 0������  �? ?�? ?�?���?���? ?�? ?�? 0�? 0�? ?�?                                                    �?  �?  �? �? �? �? ?� ? ? ? ?�?���?   ��  0��  �� �� �� �������������� �� 0��  ���  ��  ��  �� ��� �� ���� �0�� ���� ��   ��  ���  ���  ��  �� ��� 0��� 0�� 00�� 0���   ��  ��   �� ���  �� �� ��� ��� 0�� �<��  ��  ��   �� 0�� �� �� ���  �� 0������  �?  �?  � ? ?�? ?�? ?�?���?�� ?��0 ? ?�?                                                    � ?  �?  �?   ?  �?  �?  �?  �?  �? �?  ���  ��   ��  ���  ��  0��   ��  ��  �� ��  ���   ��  ���  0��  ���  ��  ���  ��  �� ��  ���   ��   ��  ��   ��  ���  0��  ���  ��� ���  ���  ���   ��  ���   ��  ��  0��  ��   �� <��  ���  0��  ��   ��  ��  ��  0��  ��   �� ��  �?  �?  �?   ?  �?  �?  0 ?  �?  � ? ?�?  ?� <�0�? ? ?�<�0�?�? ��� < �������� 0 < ���� ����  3� �0��0����  3� ���  ?��? �0 0��? �?��00 0��� �������� ������ ����0 �� �����0 0 �� ����00 ��  ?�?�0��� ? ?�?�00���?                               ��� ?����?����?��� ? ���? � ����� ���  �� � ����� �� �?�����? �� �?�����?0��0�?���  ����� � �� � �� ���� ��  ����� ����� � �� ������ �� ��������0��0������ �� ����  ?�?�?�?�?�?�? ? ?�?                                0  ?� ?� <�?�0�?�?�< ?  < ������ ��<�� �� ���  3 ��� ���  �� 3 ��� ��� 0�� �0  ?� 0��? �� �0 ? 0 �?�� �� ��� ������������  �����  0 ��� ���0��0 00���� ��  0  ?����?�?�0�?����? ? ��  <  ?� ?���� ?��0����?  0   ������� ���<0 ��   �  ��� ���?���  3 ���  0 �?  �� 0� �� ?  �0  ��  � ��  �� � ����� ����  �� �� ��  0� ������0 0 00 ��  ?  ?  ����?�?�?�0��?                                ?  0  <  ?� ?� ?� 0� <� ?�? ��  <   ��������� <� �����  �  3 �  ������ �� 3�� ��� ��  0 �0 �?  ?���� 0��0��?� ? ��   �� �� ������ ������������    0 �� ������ � 0������0�� ��  0  ?  ?�?����0�?�?�?                                  ? ��  0 ��  < ��  ?  ?� ?   ��  0  < �     0 �� �����    �    3 �? �    �� �����    0  0 �0  � �?    ?  ����      � ��  � ��   ��  ����     ��  0 �� ��   ��  0���  ? ��  ?  0  ?  ?    ?  �?������?� ���?� � ������3000   303 � ���� 00000   303 � ���� ��000 �  ���� � ���� 0000   3 0 3 � ���� 300   3 0 � � ���� �00��� �  �0 �?��������3030 ��?�0 ?��?�30��<�< 3 0 0 �� 330��0333 3 0 0 3� 300�0030 ��0 0 � �?��0030 3 0 0 � 30�0030 3 0 0 � 30�30�00 ��?0 �??�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ��������?��<<�����<<����?<<�����<<����<<����� �����          ����?<< �0<<�����? ��<<����<?���< ����<?���<<����<< ��<<����<<�������?<<�                                                                                                                                                                                                     UUUUUUUUUUUUUUUUU                                                                                                                                                                          UUUUUUUUUUUUUUUUU                                                                                                                                                                                           UUUUUUUUUUUUUUUUU                                                                                                                                                                                           UUUUUUUUUUUUUUUUU                                                                                                                                                                                           UUUUUUUUUUUUUUUUU                                                                                                                                                                          UUUUUUUUUUUUUUUUU                                                                                                                                                                          ���� ,  ���?�� ��� � ��p� �  � �� �  �  ���     �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���*      �?�?          � �   � �     ����  ��  �0 �  ��    � � � �    @        ��      � � 0 <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ������?��?��   ���������?��   ���������?��   ? �����  ?�   ? �����  ?�   ? �����  ?�   ����������   �����������   �����������    �����?�  ?�    ���� �  ?�    ���� �  ?�   ������ ��??�   ������ ��??�   ����� ��??�                                    ?������� ?    ?��������?�?    ?����������?    ?��� ����?    ?��� ����?    ?��� ����??    ?���������??    ?����������?    ?���������?    ?�� ������?    ?�� ������?��  ��� ������?��  ������������?��  ���������?��?��  �?������� ?��                  ��� �� ����0��������� � � ��� � ������� ������ �����?�?����� ����� ������� ������ ����������� � ����� ������� �� ���� ���0�0�0�0�<� ��� � ������� ������ � �����<��<���� � ����� ���� ��� �0��0��?������W��W��W��W��W��W�:W�:W�����?��:{{;_]={{;��:��:{{;_]={{;��:{{;_]={{;��:��?       ? ������6w7{7w7w_7��6���� ?       � � � �� 0� 0� 0� 0� 0� �������?     ���� � � � � � � � � ���     ��?�0� � � � �� �� �� � � � �0�0��?   ����� � � � � � �������   ���� �� �� �� �� �������� �� �� �� �� ��   ����������������?�   �? ���������������������������    ����������������� � � � � � �    ����������������� �? �� �������?     ��� � � � �? �� �� � � ����     ��?��0��0�� �� �� �������� �� �� �� �� ��   ������������������������������   �??������������?����                                                                                                                            ���?                                    �?�?                                   �?�?                                   �?�?                                    �?�?�������?�?                          �?�?���?�?�?�0                          �:�:��:�:�:�                           �:�:������:�                           p5�5�\pp�5�                           p5�5�\pp�5�                           p5�5�\pp�5�0                          ���?�������?�?                                                                                                         ����������������������������������������������������������������������������������������������������������������������������������������������������������������                                                ��                ��          ����������������������������������������2WUUUU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�UU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�UU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�UU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�UU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�UU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�UU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�VU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�ZU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU)ZU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU)ZU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�jU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�hU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�hU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2WU�jU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2W��jU�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2W�"�U�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2W�"�U�WUUUUUUUUUUUUUUUUդWUUUUUUUUU��2W���U�WUUUUUUUUUUUUUUUUդWUUU��WUUU��2W���V�WUUUUUUUUUUUUUUUUդWUU���_UUU��2[� �V�WUUUUUUUUUUUUUUUUդWUU���UUU��2k� �V�WUUUUUUUUUUUUUUUUդWUU����UUU��2����V�WUUUUUUUUUUUUUUUUդWUU����UUU��2����Z�WUUUUUUUUUUUUUUUU֤WUU? ��WUU��2��*�Z�WUUUUUUUUUUUUUUUU֤WUU ��WU���2����Z�WUUUUUUUUUUUVUUUU֤WUU ��WU���2����Z�WUUUUUUUUUUUVUUUU֤WUV?���WU���2��(�j�WUUUUUUUUUUUVUUUU֤WUV� ��WU���2������WUUUUUUUUUU�ZUUUU֤WUV����W����2������WUUUUUUUUUU�jUUUU֤WUV����U�"��2��*���WUUUUUUUUUU��UUUU֤WUV���U����2������WUUUUUUUUUU��VUU�ڤWUV��~U�"��2����*�WUYUU�UYUU���ZUU��WUV��_��"��2�"""��[UYUU�VjUU�""jUU��W�Z�?�W��"��2����*�kUYUU���UU���jUU�٤W�j5 �_�����2�"""���UYUU���UU���jUU�٤W��>�����"��2�"""*��VYUUi��UU����UU�٤W�������"��2�"""*��VjUUi��UU����VU��W����i���"��2����*����UUi��UU����ZU�ȤW���z������2�"""���VjUU���UU����j���[�|m�O�?��2�"""*��ZjUU���Ui���*���Ȥk�;=��Ԫ���2�"�**��jjUU���U��������꤫�9��?��j���2����*��jjUU)�������(���Ȥ�^4m����Z���2�������jjUU)�������*���Ȥ�m�o�[U��2����*���jUU)�����������Ȥ�Am�l�U��2����*����UU)�������(����� m�o�P��2����*����VU���"����*���Ȥ�@m��@��2��""�����ZU������������Ȥ� m0�5�@Y�2����*��*"jU)"������(���Ȥ3�m�5� Y�2��""*��������������(����;��1�5�T�2��""*������������������Ȥ3�5��9�P�2��""���*���*�������(�����;�4�1�>� �2����?��*���*�������(����������k@ �2�������*���*�������������?��?���^�2�������*���(�������(�����?�D�������2�������������j�����(��������6s�����2���o���������j����������������|0���2����������("b�����(��@���1P;s0|t��2�����������������(�� ����P�|0p��|�2��������������������� �����@;s��A�\�2������*"��(������(�������C;s��U�0�2�������*"��(������(�:����EN�|@�}�<�2������*"��(��������2�J���5M;s@����2����������*������x� ����5M�|@����2���������(������x�	����5u;s@�U��2������ޫ��������z����>�5u�|@���2�������ܣ���*�����|���T�6�M�;s@��>�2��������ޫ�*"b�����s��C����]��| �� �2����W���ܫ���^�����s��C���tS�6s ��@�2�������ޯ�( V������������| ��P�2�������������W�����Т�C������B�yP�2�������.��*"_�����Т���>�+�o��^@��2��/��������k骪�� ��������[�_T� ��2��z����[��( �鈈�� ���>��P�<D��2����?���[ ����戈�����?��j��@9�W��2���[����[ ������������������R����2��~�� l� ��9    ;� �O������P���2������ l0 p�:   �� ����6���P���2�����   �? \�:   ���0�V��:��P�@���2���������[�������������������R�����2���U��������������3��?W�����������2��jU� �[���<�;0  0���U���� ��������o�jU� �v��o3�;0  C�|U���j�� ���Ʋ�����VU �մ����??  �:oU���j�� ��Ʋ���z�jU������;  L��ZU���jW�����Ʋ���������j������>  CP�VU�����������Ʋ������ZU�j@������?  C]P�V����j�������Ʋ������jU�9�?���  S@UU�����������򾪮�UUP  ���  S]EU��j��jW�W����򾪮�i��Z�   ��  [zU������×�W�������������VU�    ��   �zU������_���������������ZU9 �������ꕪ����������������z���o��� ��ο�������jo��_��������2뫺���������������������������������2�������              �S��W�?���� ��2����� 3ê��������������P�_������ ��2��ꪻ[?��������������?�z������� ��2����W?     ����     Dz������: ��2��깮Ws9     ����     �]��j���: ��2����U0W:      ��      kP^������: ��2�����Y0��      ��      �����j���: ��2�����Uϧ�      ��      ���������: ��2�뻪�Uϫ�      ��      �����W���: ��2�뻪�VE�:      ��      ��嫾�W���: ��2�믪�VE�?      ��      �����j���: ��2����VA��     ��     ������ڪ��F�: ��2[����Z����?    ��    �����������V�: ��2�����������   ��  ���������ߪ���: ��2�����������?  ��  ����믪�۪��j�: ��2�����j髪ꯪ� �� ������ꫪ�������: ���?𫪮jꯪ����� �� ��������ꫪ�����: ���
𫪮�ꫪ������� ���������ꪮ����: ���
�����꿪��ꫪ>�������������������: �   �����ꫪ�����ꬪ�����ꪯ�����꿪�: �   �������������������ꯪ��������:      �몪ꪪ����ꪯ�𪪪�������������:      ����ꪪ�������������������������:      �������������������꪿�����꯺��:      ��������������������ꯪ���������:      �����������������������������:      �������������������������������:      �����������������������������:      ��������������������������������:      ��������?���ꮪ�����������������:       �   �: ���ꮪ������   �������:  ����������������������������������������    �                                      0 �������?�?���������� ����?�      � � �����s�777�������� p��<7p      0������s�777��������  p��<7p      0< �������?���������� ����;�      0��������;������  �� ;�      � � �������??�����<� ���<?�       0 �������?<���������� ����?�       �                                  ����������������������������������������                                              @  P �������������?�������������������������������?������_��        @  @  @                      @  P ������������������������������������������?������_��                                             @  P ������������� ��? ��? �� �� �� �������������?������_��                        ����                 ����>                �����                �� � ������ ��  ���  �: �:������ �?0  �� �꼪:�:�����0  ?� �_��U5�:���:�� �? �_��U5�:������� ��_��?���ο����  ��_�� ���ί�����  ������ ����������  �ʿ2 �?�� ?�;����?�  �0�0 ���� ���ί���?�? �����������ί��������������5_����� �����׼�:�:���:�� �������U5�:����� ���U��U5�:�� ���� ������?�?��� �������������������������������������������������������������������������������������������������������������������������������������?��������꿪�������������?���_��U�������������? ��_��U���������������_������������� �����_��������������������������������������ʿ�������?�;����?����0����������������?����������������������������������_����� ������׿����������� ��������U���������� ����U��U������������������������������                          ������             �������            ��������           ���������          �j������          ��Uՙ����?          �]e�������          �w��������        ��w��������        ��w[�������        ��w�w������?        �w_�������?        ��o��������        ��}���������        ������������       ������������       ������������       ������������       �?���������       � ���������       �  @UUUP���      ��      @���      ��      @���      ��    @ ����      ��      ����      ��      ����      ��      ����      ��     @U���      ��     @U���      �� �� ������      �����?�������      �����?@������:      �� U�:@�@��>      �� ��:@�����;      p� ��;@�?����:      p���?;@��󗪿:      p� ��;P���V��:      p�  ��*  P��:      p� �,���P��:      p�   �Z  T��:      p�   �j ���:      p�   �Z ��:      p�   �j@��      p�   �� ��      ��  ���V ��      ��  ?P����      �� �0P�����      �� 00P��j���       � �\U������        � �������        �����������        ����������          ��������          �����           �   ���           � �����           �������           @�������          0  �������         �    U����         �    ����         �    ���         ��    �����        ��   ������       �U  P�������       � �U��������?      � ���ꯪ������?    �� T�������jU��   �U P����z��jUUUU  ��U U�j��^��ZUUUU �_�U P����W��VUUUU U�U� @�j��U��UUUUU�UU�UU Uj�z��nUUUUUUUUUWU @UU]��kU UUUUUUWU5  UUW��Z �?UUUUUU]U�  U�U� ��<UUUUUUuUU U}U 0?<UUUU@�UU U ���?UUUU�UWU ����� UUUU�<U ��|��� OUUUU�<  ��������@UUUU�<���������OUUUU<<<��<�����@UUUU<<�<�?3��� PUUUU<O<�<�?3? TUUUUUUO<�3<�?3 UUUUUUUU���3��? PUUUUUUUUU���? ��VUUUUUUUUUU��@U��VUUUUUUUUUU� PUU��VUUUUUUUUUUU TUUUU��TUUUUUUUUUU�WUUUUU�?�WUUUUUUUUU��_�}���?|_�]U�WU��}�}���?|�������}_U��}�}���?|�������}_U��}�}_U�?|�������}_U��_����?�W������WUU�UU}UU�?TUUUUUUUUUUU�U�UU��VUUUUUUUUU                          ������             �������            �������           ���������          �Z�����          ��Wՙ����?          |Ze�������          �u��������        ��u��������        ��u[�������        ��u�w������?        �w_�������?        �_o��������        ��m���������        ������������       ������������       ������������       ������������       �?���������       � ���������       �  @UUUP���      ��      @���      ��      P���      ��    @ ����      ��      ����      ��      ����      ��   ����      ��  @U���      ��  0@����      �� ���M������      �������������      �������������:      �� U�:@����>      �� ��:@�����;      p� ��;P�?����:      p���?;P��󗪿:      p� ��;P���V��:      p�  ��* $P��:      p� �,���P��:      p�   �Z  ���:      p�   �j ���:      p�   �Z@��:      p�   �j@��      p�   ��P���      ��  ���VP��      ��  3P�U���      �� �0P������      �� 00��몪��       �  �\�������        �  �������        � ��������        �L��������         �������         ����������          �? @�����          ����ﮪ�          ��������            �������         0  ��U����         �    P����         �    ����         �    ���         ��    �����        ��   ������       �f  P�������       �V�U���������      ����ꯪ�������    ��P�������jU��   �U ��������VUUU  ��U U��������UUUU �_�U P��������UUUU U�U� @���ꪪ�jUUUU�UU�UU �������ZUUUUUUUUWU ��U]��kU UUUUUUWU5 ��UW��Z �?UUUUUU]U� ���U� ��<UUUUUUuUU��}U 0?<UUUU@�UU�� ���?UUUU�UWU ����� UUUU�<U ��|��� OUUUU�<  ��������@UUUU�<���������OUUUU<<<��<�����@UUUU<<�<�?3��� PUUUU<O<�<�?3? TUUUUUUO<�3<�?3 UUUUUUUU���3��? PUUUUUUUUU���? ��VUUUUUUUUUU��@U��VUUUUUUUUUU� PUU��VUUUUUUUUUUUUUUUUU�?UUUUUUUUUUU�WUUUUU�?�WUUUUUUUUU��_�}���?|_�]��WU��}�}���?|�������}_U��}�}���?|�������}_U��}�}_U�?|�������}_U��_����?�W������WUU�UU}UU�?TUUUUUUUUUUU�U�UU��VUUUUUUUUUH�Z�������C��(��a� J� Z��/ �ƥ������� ��� Z��/ �ƥ�C���d� ��� � �v� � �t� � ���  �����  ������ ��� � � ��z�h`�� ���0� j�`�1��� �� j�`�Zd��0� 08�(� ��0�8� � �8�0��N�0d �
����e�轞�i �����T�e ����i �� �%���00����e��i ���z�`Hک �� � �ȩP�d�(������ ��P��� �� �� �28�� �8���8���8���i��i� �Ʃ@ �ƀʩ� �M�����d%d�� �Ȣ ���� �i������d%d�� �ȩQ� �H�ࠐ�  �h��  ����� �����W�ـ�d ddd�(���������	 ���� �Ʃ� �Ʃ� ���	�	���� �Ʃ� �Ʃ� ���h`H�� �M�����d�����% �h`H������ ���ʽ��� �i�����%d�� ������� �i��d��d%�W� �h`H�Z� �� � � 4ũ� �� ���>��Z��	���  ��� �����n��	���  ��� �����?�����	���  ��� �����Z��� �8� ��� ����� �;� ��� �Ʃn��<���  ��� �����������	��� �=� ��� ������	�Y��� �� ��d# 4�H��� 1�hɿ�" ���#���Y� ��d#�ܥi� ���#���������# ���#���� ����#���8�� ���#L1������d	 ���� �Ʃ�	 ���� �����z�h`H���� ��h`H�V�� ��	�?� ��h`H�Z� H�H�H�H�H�H�H�H�H�H�H�	H�
Hd���� �F��$��P�d% �ȩ �� � � 4ũ� �� ���Z�� ����� ���� ��` �����
��n������ ���� ��` ��������	�䩂������ ���� ��` �����	���	�Y��� �� ��d$ 4� �Ȣ�� 1�ɿ�" ���$���Y� ��d$�ۥi� ���$���������# ���$���� ����$���8�� ���$L������d���� �F��$��P����% ��h�
h�	h�h�h�h�h�h�h�h�h�h�h� z�h`Hک �� Ʃ��d����
� dd���� ��&��Y��Z����	�� �ƀ� 4�������L��������L��H�Z ?ǥ	� �� ����U�
��������
� � �
 ����������i0��i ���z�h`H�����dd ��h`H�� ��h`d ��`H �ȥ�dd�� ���� ��h`�  ����� �ƭ  ����H�  ����h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               x���� � ة��  ��� � � � � �ύ& ��" � t ���d���� � �������� �� !� 4� � ũ ��XL���@H�Z�' )�
 X���# �d��$ �% (z�hX@H�Z� � � �����



	� ��� ��� ��� �d:� ��z�h`ڢ
L�����������:���`Zڢ��������:���z`H�Z� ���� � ȹ��� � ȹ����y�����t� �  ����� ��Ȝ � ��z�h`� ������ � Ŝ � � � � � � � �* d�d�� ����d�`�������� ť�� ���  [�朥�ń� e¥������� ť�� ���  ��来�Ņ� �¥����J�������� ť�� ���  �å������� ť�� ���  �暥�ł� ��曥�Ń�  å���� 	� w�`������ȱ���ȱ���ȱ��~ȱ���)
��U����U�����)0��ȥ���������Ȅ�d�d���� �L�¤� ��� �
��� �d���Ȅ�d���������ȱ���ȱ���ȱ���ȱ���)
��U����U�����)0��ȱ������Ȅ�d�d���� �� ��� ��)��	����d� ��`������ȱ���ȱ���ȱ���ȱ���)
��U����U�����)0��ȱ������Ȅ�d�d���� к� ��� ��)��@Ы����d� e�������ȱ���ȱ���ȱ��ȱ���)
��U����U�����)0��ȥ���������Ȅ�d�d���� е�� ��� �
��� �d���Ȅ�d�����
����������ֱՅ�ȱՅ�`��
����������ֱՅ�ȱՅ�`H�Z�~)?	@���~;��%����������)@��J��������8������)0��Ȅ������Ɔ��d���� z�h`H�Z�)?	@���;��%����������)@��J��������8������)0��Ȅ������Ƈ��d���� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������ƈ��d���� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ɖ��d���� z�h`� `� `H�Z������ͩ��̅���)?
��;����;���d� <�z�h`d��* d�`���΅�ȱ΅�ȱ΅�ȱ΅�)
��U����U��ť�)0��Ȅ�d�dƥ�� 4�d�`H�Z�����L�ť��ʥ�;��)��ʤƱĪ��)@��J��ʅʥ��8��ɀ��)0��ȄƱ�����ƥ�dƥ�)����)����
�@��������ʍ( ������* ���å���� <�z�h`H�Z�  �à  ��d�d������ ��  � �� � 	ũ���z�h`H�Z��� ���� �d���)?ź�D�� �>��
�����������轂��������d�d�� ������)������ �¥����� e� 	�z�h`�Z����� ���� ��z�`H�Z�� � ?Ǣ � ڱ �����������i0��i ��e��i ���z�h`ڦ� ���1�
���Q%��`H�Z�
�����轞���� ��e��i ����e��i �z�h`Hڦ�T�e ����i ��h`H�Z�)���!�� �JJJJ� �ǥ������!�)��!��"�� �� �ǥ������!z�h`xH�Z��a��$�F�b��%�>�c��&�6�-��'�.�:��(�&�f��)��?��*��,��+��.��,��e��-�������������T������� �%��Ȳ%������� � z�hX`H�Zɀ�8�
�������LW�
�����轺��� ��$�3�a�'�b�#�c��-��:��f��?��,��.��e�8�7� ��Ȁ�z�h`H�Z ?Ǧ� �%�������������i0��i ��e��i ���z�h`�  ���L�� ��`H ������h`Hd d����(� ��h`�  �����F �Ʈ  ���� �ƭ  ����`���&  9� �� �թ �� � @�d1d-d '� � ��d.�  ��� v��/�/��� G�d/��  ���L���� �ʀ����Щ�� 1� q� �� �ѩ�  � �� _� �� �ͥ-� �� :� :� :� �� *ͩ�� 1� � �� c̥&ɪ��ύ& �� I� I� S�L�  ���L����-�-�
�� �� �d1d-d '� � ���.�.��L`�d.LGɩύ&  շ���& �$�	� �� ƀ���L��L&ɠ ����� ��4��`H���� H� ������ H� ������ H���� h�� ��4��h`HZ���� H�� H� ��h�� ��4��zh`H�Z� �.�	� i
�����יB ������,z�h`�� �=��# 0� v�d.������-��  1� P�����`H� ��d  ���� c̥ �����-L˩�*L�������L˩�*L�����  c̥ ����U���-L˥��J��*�g�������8��*�q��$�ύ&  շ���& �$�	� �� ƀ*��L��L&�������L��� 1Ʃ�d- :� 1� :�L��  ����L���� 1� �� � �� 'ѥ��L�ʩ�� 1� ��L���h`H�  ɩ�� 1����	��� �̀ � Ѐ�����1�B I�B  Ѐ���$�ύ&  շ���& �$�	� �� ƀ���L��L&������жL���h`��� �̩� I� �� �� ��`��� �̩` I� �� I�`Hd ���� �&�������
����&� ��U� ���&h`��e*�8��*��� ��`�8��*��e*��i �� � �� '�`Hdd�	����-�	�� �#���=��� ��h`Hd Х ��	i� �1��� d1h`Hd Х ��	8�� �1��� ��1h`H�Z����
�-�d��+��e+��i ����e��e��z�h`H�Z�,� �B )���יB ��B )�B ����z�h`H �� Υ-�	�J >Υ-��A eΥ-��8 �Υ-��/ �ϥ-��& �Υ-�� �Υ-�� ϥ-�� Gϥ-��d-h`H�Z� ����B �*ȹB ��*���B ȥ*�B � �����z�h`H�d- �ϥ-�"�0�+ |ϥ-����B )������-��	�-�h`Hڥ-�� �ϥ-����0�+ �ϥ-����-�h`HZ� �B )��+ȹB )��+�ȹB )��+�����+ȹB )��+�����-zh`HZ� �B )��+ȹB )��+�$ȹB )��+�ȹB )��+ȹB )��+�����-zh`H�0�+ |ϥ-�� ��h`H�Z� ��B )��+������B )��+����-z�h`H�Z� � �B )��+����B )��+��+��������-z�h`HZ� �B )�ɰ��+����������B )��+��+�������-zh`HZ� �B )�i�+ȹB )�����+��+i�+����-zh`HZ�0�+� �B )��+�'ȥ+i�+�`��B )��+����ȹB )������-zh`HZ� �B )�+ȹB )�+�	�����-zh`H��� H� � �� ��h� h`H��d��dd����� �Ʃ��h`H��ddd dd�(���� �Ʃ� �Ʃm� �Ʃ�� ��dd �� b�����d��� �� b�������d�����d����  �Ʃ��� ����� �Ʃ� ���
�� �� �� �d�o�d��d�������  �Ʃ��d�� �����d ��dd�� ����� ��h`H�Z� �q���n�� �}����������d�����
��	�e���d��d ����пz�h`H�Z �ԩ�)� �_��(Z ��(�(JJ�( �� �ѩ�� 1Ʃ� �� ��z����z�h`H��ddd�)i��F���� ��h`H�Z �ԩ�)� �B �*�_��(Z ��(�(JJ�( �� � �ҩ� �� ��z����z�h`��������d�*)

��)i��(�  �ƥ)i9��(i� �� �ƥ*)�JJ8��d���4��)i��(�  �����)iB��(i�  ��`�*)��0� ӀT�@� "ӀK�P� kӀB�`� �Ӏ9�p� �Ӏ0ɀ� �Ӏ'ɐ� �Ӏɠ� Ԁ�� ?Ԁ��� \Ԁ ��`���� �ԥ)i��(i�  �ƥ)i6��i� ��` �� �ԥ)i!� ��`���� �ԥ)i��(i�  �ƥ(i�  �ƥ)i6��(i� �i� �ƥ(i�  ��` "� �ԥ)i!��(i�  ��` "� �ԥ)i!��(i�  �ƥ(i�  ��` �ӥ)i��(i�  ��` "� �ԥ)i��(i�  �ƥ(i�  �ƥ)i(��(i� �i� �ƥ(i�  ��` �� �ԥ)i!��(i�  ��` �� �ԥ)i��(i�  �ƥ)i/��i� ��`�5��	� �ԥ)i��(i�  ��`���������*)�

e��)i��(i�  ��`�����*)
�
e�`�����*)�8�J�JJJe�`H���K��)��(�  ��h`H������  ��h`H���M�����  ��h`H�#���� ���V� ��h`�)��(� �7 b�� ����)iL��(� �7 b�� ����)��(i6� �L b������)��(� �L b�����`H�Zdd� J��*��J��**���T�����������W�%��[�%�z�h`� ���dd` <�d"� Uǩ�"� U�`H�� �� ��h`H�� �� ��h` <�d"� Uǩ�"� U�`H�� �.� ��ddh`H�� �� ��ddh`H�� ��d!��"� U�h`H� � �F�d!��"� U�h` �� �� ��`���&  �� �� � E� j�La֥6����s��t�s� �` � �t����L�֩ �&�ύ&  S�`�ύ&  շ���& � �� ƥ$��hhLS���hhL��`� �5��6dsdtd7d8��9� tR��+����w`�� �n��# 0� v�dk���� 1� �� �� 8�� �m� ���k�k��� ��d7d8d9`�`���9�� v�d7d8`�9�� ��` '� �ȅR�� ����L���� �� ��`ɿ� �� ��`��� �� r�`��� �� ��`��� �`��� ��`��� �� ��`��� ��`�u��`�v�v���` �� �� ��dv`H�Z�� �יJ ���\��� �B�k� �� �k��L�׵J�� ��\�� ��B�� ���\��z�h`H� �� �d ddd�'�����P�d �� �� �� �� �� ��d �P����(�P�) ��� ��� 0ȩ� ��� 0� � I� \� 9ʩ� ��� 0ȩ� �s�� 0�h` �� ��`d �%�dd�&������d`d dd)���( ��`d dd(���) ��`d ������(���) ��`��� d���(���) ��`�D� d�D�(�P�) ��`�O� �P��O�(���) ��`�5��6��� �����d!d"� Uǩ�"� U�`���d!��"�`�S��� �� <� U�`�T��� �%� <� U� ��`H�Z�`�� ��L�� `ݥS� � K� R� � I� \� �� ��L�� �� �� �ߩ�`�d �� �� � ��z�h`�p�� ��`�B)��k�C)��k���b`�� �Z����<� �� ��du`�� d�s�d����
�d�)� ��`�;)����+ �� �٩�u �� ��������M��� �� �٥w�� ��`��w�� �s����
� ��� d�}�d����
�d�)� ��L)ک�w�� �}����
� �� ��L)ڥS����V`J�V` �ڥ6� �&�5�V�  
� �� L� zީ� �r�� 0ȩ�eda`��a�58��V�5�6� �6� �`Hڥ9��d9�9dx� t:������(�R�)�8�� �*�B i��\�8���� 1� +�G�(��)�8�� �: ���[�8���� 1� +��(�R�)�8�� �*�C i��\�8���� 1� +��(��) �� �� �Ʃ��� 1� +�S�(��)�8�� �*�; i��[�8���� 1ƩS�l��m�h`�� �Z�� 0ȩ� �d�� 0ȩ� �s�� 0ȩ� �}�� 0� �ة�u` 8�� �c���� �� ��`H�� �d��&����P���d% ��h`H�� �d�dd�(��&����d ��h`H�� �d����(�d�) ��� �d���(�|�) ��� �|����(�|�) �驛� �d����(�|�) ��h`�� �d��&��� ��` `� � I� \� �� ��`�`� ��S� �
 �� �� R�` T� R�`�d��$�e�� 
� �� L� ��� �r�� 0ȩ�e`�e��de *ܥS����SL#�FS�5�eS�5�6i �6� ٥S�W �� �� ��a�� � ;� ��`�� �#�� 0�` {�d �Q��(��N� �� �� ��`�� �����O� �� �� ��`d �G����	� �� ��`d �/����	� �� ��d �;����	� �� ��`H�� �G�( ��h`H�� �S�( ��h`H�Z� H �h� ��dd������F�d ��z�h`��) �`H�� �G��  0�h`H�� �=��	 0�h`�� �d�` Bީ 0�` Bީ 0�`H Bީ 0ȥS��� �d� <� U�h`�h��� � 0�` �ީ 0�` �ީ 0�`�n��� `�`� ��S� �
 �� K� R�` T� R�`db�c���r�� ��` ��`�e��de *�dd�c� ��miL�ޥmi�m�(�R�)�7�ׅ*�\�B i��\�7 �n�p�^� ��ni
���pL2ߥp��)�p��L?ߥ\���c� � ��`�r����i`��j`�c���r����g`��h`��z W� ��a� � �� ;� �� ��x�6� �`�5����s�t` �� �� k�i���g��` Z�` �ޥj���h��` ��`H� �^� ��ni
L�ߥn�p�h` �^���n�o`�ni
�o`dnd^� �B #���\��`dnd^� �: #���[��`JJJJ���^�ni�nLY���
�ni�nLY���en�nLY�ni
�n` �� v�Z�B��\ �ߩ�r � ��`�[�m�(�R�)�8�� �C�* i��8`�^�_�\�]�p�q� �B�J��\��`�_�^�]�\�q�p� �J�B��\��`�T�8�S�Tإh��	 �� ��L��a�� �� W� �� S�L��f�� v�L��� �� �� �L��� �� �� ٥g�� ��W�X ��X�W ��L;�a�� ��LA�f�� C�Ld��� Q� �� �Ld��� _� �� � ;� ��` ٩� �R����L� ��S�(�R�)�Z�* i�`�`� ��S� �
 �� K� R�` T� R�`�e��de *ܥc���r�� Z�` ��`LV� ��r�� W� �� S�a�� ��y� �Ln�o��ӥp��'�\��!�o���[�� #� �� �Ln� 4� ��Ln�o���[��	 G� �Ln�p�o� #�Ln� G�Ln� ?�Ln�p���\��	 4� ��Ln� ?�c� �2�f�� �L���� � �� ��L���� "� �� �� � ;� �� ٥6� �`�5����s�t`�o���[��dy �`��y �p���\��
 � �� L�` � s�`�
� ���� 0�`�� �(�� 0�` �� L� ��` �� L� ��`�T�eW�W� ���f` �� ]��f` ���f`��f` �� ]� �� ٩�f`��5eV�5�6i �6�WeV�W�` ����WeT�W� ]� �� ٩�f` �� ����TeTeW�W�`�5�eT�5�6i �6�`�p��/�\��*��% 2�k�����B)��`��C)��`�	�D)��`�` ��` �� �� ����WeT�W�d �1��" 0� ��dk���� 1� +� 8�d �0� ���k�k��� �� �dW`dk�B)��p��k�C)��p��k�D)��p��k`Hڥc���p��	�\���h`�g%h�� �^� �(�:)��`��;)��`� �� �^� � �ni
�� �n���oL��[����h`�li�l�(��)�7�צ[�:�* i� +� +��[�7` �� �ة1��%� ��`�W��� �1� <� U�`�� �G�� 0�`�� �G�� 0�`ڢ  ��������`ڢ  �������`���� �F�dd����	���`�� �G��z���Ll�! 0Ƞ  8� �Ʃ�� 1� � �����`�� �x�� 0Ƞ  8�� �w���� �Ʃ�� 1� � �����` {ݩ;�l� �li�l�(��)�:�* i驅�� 1� +���[�� �ةS�l +�`L��L��H�`���d���6� ��5�S��e�� 
� �� L� ���eL��p�
����e�� 
� �� L� ���eL��5�8�S�5�6� �6�TeS�T� � I� \� 2� �ޥx��) ��L��e�� 
� �� L� ��� �r�� 0ȩ�edxh` zީ� �r�� 0�`�� �n�� 0�`�� �h��
 0ȩ� �h��� <� U�`�`��`�b� �!�e�� 
� �� Lܩ� �n�� 0ȩ�e`�a�� y�6� �	�5�k�LA� ��Le�6� �*�5�S�$�e�� 
� �� L� zީ� �r�� 0ȩ�e`��cdbdd ��de �� ��`�S�eV�k�`�� �R����L� ��`�C�Z ���(�R�)�B�* i� k� +��(�m�R�)�8�� �*�C i��8��r ��5�8�S�5�6� �6�TeS�T�Ui �U� � \�`�
 �� �<�� 0�`� �<��� <�d" U�`�
 .�� �G�� 0�`� �G��� <�d"� U�`� � m� 0�`� � m� 0�`� � m� 0�`�� �<�`� .� �� 0�`� .� �� 0�`� .� �� 0�`�� �G�`Hڥ`��L�� � Rݥ6� ��5���d |�L���� 1ƥS�i�S�T�58��5�6� �6� � I� \٥S�� r��h` `� �� ��`Hڥ`��Lf� I� \٥S��	 �� ]�Lf� � RݥS� � K�Lf��� 1ƥS�8��S�T�5i�5�6i �6� � I� \��h`H�Z���0�� � ��(�(JJ�( �� � ��z�h`H�Z��� bե �(�
��)����� ��z�h`Hd �Ʃ��h` �ȩ �� Ʃ��&  �� �� s��2 �� ��� �� a� �� �� ��d 3֮  ������� �Ʈ  ����  ���� ��L�����-L$���� ����$� �頻 �� �� �� ����3�  ���� �� 1� ������$� ����� ��d3����������i��
��� �� 1� �� �� �� ���# D� c�� -� -� -� -��� 1� �� ��d 3� c̥&ɪ����L~�'����' ;�s� �� ;�L��L�����M c̥ ���
�������-L$��*LA��� 1Ʃ� :̩�� 1� :�d-L�� ~� �� 3� ��L����#�ύ&  շ���& �$�
��L��L��d� �L�����L��� I� I֩ύ&  S�L��H�Z��'�2� P�� �2� n�  ɩ�� 1���(����'���'�٩�'�����ڥ'���'�ũ�'��z�h`H�	������ �x�dd�"� �Ʃ�� P��  n�  ɩ�� 1���0��%�ύ&  շ���& �$�
��L��L�� �� �L����L��h`H������� d�M��� ��h`H���d!d"�' U�h` ����Y� ��` I� ��
��^� ��` I� ���� 1Ʃ@ I� ��`H��d������� �� ��h`Hddd������� �K��� ��h`H�Z�����d�	��� �':

�� �������� �������z�h`����� �̩� I� �� I�`Z���*����e*��i �����z`��e��e��`dd� ����$������ d �Ʃ�������� �� �ƢX�� ������$� ���� �ƢX�� ������
�� ����d����  �����^�����(�����^�d  �� ;�� ��d��������� ����P� ������2� �������� �������4�� ��������d�
������ �� �Ʃ,� �ƩD� �Ʃ�����
��� �� �Ʃ��
��"� �Ʃ��	��9��D� ��d��������� �0� �Ʃ���  �Ʃ��� ���d������S�d�� d �Ʃ� � �Ʃ� �� �Ʃ� �!� ��`�����(��d d���l� ����ɟ��`����dd��� �������� ���� ������	����� �������� ���� ������`����d�&� ����� ��`��  �Ʃ
�  �Ʃ�  �Ʃ�  ��`������
���d���� ��4`�2�:�J��;�K��<�L��=�M�ڢ �: r�
�

e� ��8� �� �:�'�� �:��:��4�ҩ� �i
������J�K�L�M�J�:�K�;�L�<�M�=`H�������dd���� ��h`HZ�� � � 8��  {�����zh`�:�'�� �:��:`�:�'�� �ȱ
�

e� �ƴ:`H�Zd�d�d�dک�0�  r� ��
�

e� �� ��8� �� ��4�ܩ� �i
��0�0���������ک�� �J��'�J��J�J�:��4�멀 �Ƣ ������3�
���4��L���4�4�L��z�h`Hڊ
����������h`H�Z� �J�'����%�� �i� r������ޥ'��0�`�����������`� ���D� �� �<����4��3��,�����������2� ������ ��������L��L������e���Q��� ����g���	�_���
�W����O� ���G����?����7����/�'�����L��������������
��� ��� r�d���i
�-z�h`����ύ&  ³����# �ύ&  � W��#���L��LS�L� �� ��� ��� ��� �� �� ��� ��� ��� �� ��� ��� ��� w�� w�� ��� ��� ��� �� ��� ��� ��� �� �� ��� ��� ��� ��� ��� ��� ��� �<�� T0��     ��0�  0�  0�  ����0�  0�  0�  ����0�  0�  0�  0� .�� �� �� �<��0�      � ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �$�� �$��T0��T��     �T��@��.$�� �$��0���� ��� ��� �$�� �$��     �T��@��.$�� �$��0���� ��� ��� �$�� �$�� �H��     � ��     � �0�� ���     �T0��T��     �T��T��T��T��.��T��}��}�������� �$� T$� �0� ��      �����}$�h$�T0�T�.�� �$�T$�     �����}$�h$�T0�T�.�� �$� �$� �H�     �T0�T��     �T0�T�     �?�J��� �   �� �   i�s�����������������	 �       � 
	��     


����������y�����y�!���  ���3����3�����)���   � � � � � � � � � � ~ �     � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �     �     � ��� ���     � ?��� ?���     � � � � �     � �	� �	� �	� �	�     � �	�� /��     �T��T���� �� �� �|� �|� �z� �z� �w� �w� �u� �u� �s� �s� �q� �q�     �&�������������������������$�����,�������������ص^��������� �Y�V�ƃB�J���Q�a�q�M���7���ʏX�֗����    �8���P�             �!�            B�r���҂�2�b����"�R�������B�r���҅�      2�2�r����2�r���j�"�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____ #AFEJDEKBCDLBKGHBIJ@HJ
	                                                     	
	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRRRQPONMLKJIHGFEDCBA@?>=<;:9876543210/.-,+*)('&%$#"! 
	    
������~vnnz��nz��nz��E<



���?0�3G[ 0P$o��P02 !�r3RA��qaS��B����b@`C󒠂��c�2��Qp��0���s����1��P�� �4�G�S�d�n�y������������������������#�(�1�:�C�L�W�b�f�j�}�������  aPUSHaaa$aPLEASEaPLACEaBETf$PRESSaA-KEYaTOaDEAL$YOUaLOSEaINSURANCE$MINaBETaISa$aNOaMOREaCREDITf$SURRENDER$GOODaLUCKf$YOUaCANeTaDOUBLE$DOUBLE$ONLYaFIRSTaaaCARDS$CANaBEaDOUBLEDfaaa$CANaBEaSURRENDERED$YOUaWINaINSURANCEf$BLACKaJACK$TEAM:$:WINaa$:LOSEa$aYOUaCANeTaSPLITf$:PUSHa$BANKER$PLAYER$BET:$aaSTANDa$BANKROLL$YOUaWINa$YOUaLOSE$aaaTAKEaaa$INSURANCE?$YES$NOa$INVALIDaINSURANCEa$FIVEaCARDS$YOUaBUST$BONUS:$SHUFFLE$8?FMT[bipw~�o{��o{��o{��$$$$ 	$-6?HQZcnz��nz��nz��f�>������ 
	 	  		 	
  	 
	
  		
 	
   P�   0@P`p��������  0@P`p��������  0@P`p�����а���������������������������������������������   ]� �_�