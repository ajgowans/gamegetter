                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��\UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�? ���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�� ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��8��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�>�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU � �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU �{UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU=� �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��? pUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��@=�|�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU= ��  �_UUUUUUUUUUUUUUUUUUUUUUUUUUUUU��� � ��?�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�  4�r��WUUUUUUUUUUUUUUUUUUUUUUUUUUU�_��  ��� ?�UUUUUUUUUUUUUUUUUUUUUUUUUUU �� @�* 0 _UUUUUUUUUUUUUUUUUUUUUUUUU�  T� @� ���UUUUUUUUUUUUUUUUUUUUUUUU�  P�  _    �_UUUUUUUUUUUUUUUUUUUUUU�  P�?  �   ��UUUUUUUUUUUUUUUUUUUUUU? �*@�?  t�* ��UUUUUUUUUUUUUUUUUUUUU�   �@�?    �* ���WUUUUUUUUUUUUUUUUUUUU
��B��    * ��V_UUUUUUUUUUUUUUUUUUUU�V���Ε�    �* �jU�UUUUUUUUUUUUUUUUUUU�@���ϊ���   �*��Z�UUUUUUUUUUUUUUUUUUU5T�����W�     �V WUUUUUUUUUUUUUUUUUUT������W�    ��U \UUUUUUUUUUUUUUUUU�@��U��_�?�����j� pUUUUUUUUUUUUUUUUU5T��_UUU=S�? ���?�Z�+ �UUUUUUUUUUUUUUUUUE��UUUU�C�? ����V�  WUUUUUUUUUUUUUUUUC��_UUUU�C�� �������+  _UUUUUUUUUUUUUUU�P��UUUUU��������@�6� �{UUUUUUUUUUUUUUU5T�_UUUUU� ��󯪪*P�*2�xUUUUUUUUUUUUUUU��UUUUUU� ����VUUE��#<�UUUUUUUUUUUUUUUC�_UUUUUU� �:��UUU��/�_�WUUUUUUUUUUUUU� �WUUUUUU5 T*�jUUU��W��C^UUUUUUUUUUUU���UUUUUUU5 T��Z��U��C\UUUUUUUUUUUU@�UUUUUUU5 P)�V���WU��pUUUUUUUUUUU� P�_UUUUUUU5 P	�U ���WUU�?
�UUUUUUUUUUU� O�WUUUUUUU5 @` �"�UUUU�j�WUUUUUUUUUU5 ��WUUUUUUU� @P �
UUUU�WUUUUUUUUUU5���WUUUUUUU-  U ��\UUUU�[^UUUUUUUUUU5���UUUUUUUU-  T ���_UUUUկ xUUUUUUUUUU5��UUUUUUUU�     *�WUUUUU�pUUUUUUUUUU���_UUUUUUUU�     *��UUUUUU�V�UUUUUUUUUU�sUUUUUUUUUU�     ��xUUUUUU��WUUUUUUUUUUUUUUUUUUUU�    ��}UUUUUU�Z WUUUUUUUUUUUUUUUUUUUUU�
�   �j|UUUUUU�n^UUUUUUUUUUUUUUUUUUUU��    �_UUUUUUUk\UUUUUUUUUUUUUUUUUUUU��+�
� �+\UUUUUUU�xUUUUUUUUUUUUUUUUUUUU����* ���\UUUUUUU�pUUUUUUUUUUUUUUUUUUUUZ+�?� ��WUUUUUUU�pUUUUUUUUUUUUUUUUUUUն�������WUUUUUUUU�UUUUUUUUUUUUUUUUUUUչ*�������WUUUUUUUU-�_UUUUUUUUUUUUUUUUUUe�
�������WUUUUUUUU� �WUUUUUUUUUUUUUUUUU}��������VUUUUUUUU� |UUUUUUUUUUUUUUUUU����������VUUUUUUUU� �UUUUUUUUUUUUUUUUUɭ��������ZUUUUUUUU�  �WUUUUUUUUUUUUUUUU����������ZUUUUUUUU�  WUUUUUUUUUUUUUUUU���<������ZUUUUUUUU�* \UUUUUUUUUUUUUUUU�?� ������jUUUUUUUU��
\UUUUUUUUUUUUUUU�����������kUUUUUUUUU��
\UUUUUUUUUUUUUUU������������UU������U��*_UUUUUUUUUUUUUUU��U��������U��UUUUU�_�_UUUUUUUUUUUUUUU��@�����������UUUUUUUU=WUUUUUUUUUUUUUUU��PUe���������WUUUUUUUU�WUUUUUUUUUUUUUUU�� U���������UUUUUUUUUUUUUUUUUUUUUUUUUU�?@Ue�����?�_UUUUUUUUUUUUUUUUUUUUUUUUUU�?PU��������W����������������jUUUUUUUUU�PU�������_�WUUUUUUUUUUUUUUUUUUUUUUUUUU�PU�������O�WUUUUUUUUUUUUUUUUUUUUUUUUUU� UU�������_�WUUUUUUUUUUUUUUUUUUUUUUUUUU� U��������_UUUUUUUUUUUUUUUUUUUUUUUUUU5 U���?3  |�UU�����WUUUUUUUUUUUUUUUUUU5@U��_������UU��WUUUUU����WUUUUUUUUUUU5@Ui�W�����UU�U��UUUUU�WUUUUUUUUUUUUUUUPU��W����? T�W�����wUU�_UUUUUUUUUUUUUT���Uգ�  ?T�_�_�U�_U�_U���_�UUUUUUUUUU U��UU�*
��T�_���_�WU�WU��U�WUUUUUUUUUBUaUU�*��W�_�U��UU�U��W��UUUUUUUUUUJU�_UU-
 ��W�_U��_U��U�_�W�_UUUUUUUUU�@IY�_UU��
�T�_U��WU�U���W�WUUUUUUUUU�PIY�WUU-� �WU�_U��WU�_U���W�UUUUUUUUUU�PR)�WUU�  �C��_U��WU�_U����UUUUUUUUUU�PP��UUU�����_U�W��_U��U�UUUUUUUUUU�WU��UUU�  ����W������_��UU�UUUUUUUUUU�T�UUU� ����U��_������W��_UUUUUUUUUU��_UU������������������������jUUUUUUU�?U�WUUU�  ��_U�UU�U��_��_�WUUUUUUUUU�?L�UUUUU  �UUUUUUUUUUUUUUUUUUUUUUUUUU��\�UUUUU  �TUUUUUUUUUUUUUUUUUUUUUUUU����U�����
��������������������jUUUUUU�����_UUUU� ������_UUUUUUUUUUUUUUUUUUUU���WUUUUU���_UUUUUUUUUUUUUUUUUUUUUUU�?���UUUUUU��U}UUUUUUUUUUUUUUUUUUUUUU� ���_UUUUUU���}UU����UUUUUUUUUUUUUUUU5 ���WUUUUU��� U�UUUUUUU��VUUUUUUUUUUUU= ���UUUUU����DUUUUUUUUUUUUUUUUUUUUUUU ��UUUUU���� U�_UUUUUUUUUUU�UUUUUUUUU����_UUUUU?��?� �_UUUUUUUUUUU�WUUUUUUUU����WUUUU�
���V�WUUUUUUUUUUU�WUUUUUUUU� ��UUUUU� �����WUUUUUUUUUUU�UUUUUUUUU5�b�WUUUU��  ���V��U��U�_UU�UUUUUUUUUUUU=�Z�UUUU���  ��U��U�����W�_�_UU��UUUUU#V}��_U��� ���U��W���������_�_��WUUUU��� �U��0��P�W��W�_�}��W���WUUU� J����W���� ���_���W_�W_������WUUU� X����_=�� � R�_��_��_��__���_}��WUUU5��}?��|?�������W��W��W���_���W�UUUU5��_?0 ?���������W}�W��W���}��_�UUUU����  ��=��������U}�W���������_�UUU����  8��꿫�����U������_���_����_�_UU��H� *����_U��U�����_���W����W�_UU��_�   ����_UU�WU�����W��}U���W�WUU��W�  �����_UUUUUUUUUUUUUU}UUUUUUU�UUU=?U50 �����UU�����jUUUUUUUUUUUUUUUU���_��������UUUUUUUUUUUUUU_UUUUUUUUUU���_U5   �����UUUUUUUUUUUUU�_UUUUUUUUUU�<�WU5�:���W	 UUUUUUUUUUUUU�WUUUUUUUUUU���_U������W��UUUUUUUUUUUUU�UUUUUUUUUUU=�U���n�UU�UUUUUUUUUUUUU�UUUUUUUUUUU��U���~�UUUUUUUUUUUU�WUUUUUUUUUUUUUU��   ��^�UUUUUUUUUUU�W�UU�_UUUUUUUUUU��?�UU� ���jUUUUUUUUU�U�_U�WUUUUUUUUUU����UU���_UUUUUUUUUUUuUU�U�UUUUUUUUUUUU���UU�����jiUUUUUUUUuUU�WUUU��UUUUUUUU��UU�������VUUUUUUUUuUUU�_UU�_�WUUUUUUUU�UUUU��g��eUUUUUUUUU�UUU�_UU�UUWUUUUUUUUUUUUUUe�����VUUUUUUU�UUU�U�_UUWUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U�W�_�UU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��WUU�_UU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU}UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���_UUUUUUUUUUUUUUUUUUUUUU��������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������                 �                �              0< �              0< �              �< �              �< �              �� �              �� �              �? �             <�? �   ;          �� �  ��          p� �  ��          p� �  ��       ����� �  ��       ����� �   #      ����� �   �     � ��� �   ��     L�� �   ��     ������ �   �?     �TU�� �   �     �_U�� �   �     0\U�� �   �     �WU=?� �   �     LUU*� �   �     ���O� �   �     ���O� �   �     ����O� �   �5     ����O�? �   �5     ����O�? �   �5     �����? �   ��     ����? �   ��  ������? �   �V�� �? ��? �   �V�   � ��? �   �Z}      �0� �   �jU5��    ��� �    �U5�<    ��� �    [U�(>     ��  �    ���:     �?  �    ���: �  ��  �     ���;  
 ��  �        0* � �   �        �   ���   �        
 <�*:   �        �  ���>   �          ���   �       � ���   �       � (���    �       0  ���;    �          ��?    �       ���/��    �      �33��    �      �?���?�     �         �     �     ��   �      �     �  �?�      �       ���     �    � P1 �0     �    �  �       �   �   ���     �  �� 
�W�0     �  ? �pP�<  � � � U
  @�  � � TU=�  @��  �� ��@U�"� �����? �\PT���@��?���3��WUU����@���������UU���/��@�>3 "����sUU��?���V �3 �����UU��T�*�V@�� (����oU��O����V@�?̠������U)?�����V@�?� �����o�ꯪ꯾�VA�?̨��������������ZQ�?��?   ����������ZQ���;    ������  �k���     �����    �����      ���      ��       �������������������������������������            ? �           �� �           ���           <3�           ���           ���         ����         �03�          �+ �          ��          ���          ��� �          � � �           � �           0 �           �? �           = �           �? �           : �    ��
    : �   પ�    : �   ����   : �   ����   : �  �����   : �  ����?  �: �  ���   �: �  ���   �: �  ���    �: �  ���    0
: �  �?��  0�: �  ��?  L�: �  ��� ���2 �  �    �@�2 �   ?  �0���> �   �   0��� �   � ����W�  �   �� ���:  �   0� � ���  �   �� ���  �  ��  ����   �  0� ����?   �  0 ����?   �   �A��   �   �_P��   � �� �T��    � � ?�T�?    � �> ��GU�?    ����  �W��    ������W��    ������Q<�    ����?�T>�    �ï����>�    �������_���     ����������     ����������     ����������     ������ ���    ������_@���    ������P���    �������>��    �����u����    ���Q��?�    ��� ��?�    ���PA����    ��� P����?    ���V ����?    ���������?    ����je�����    � ���������    � ���������   � ���������   � ���������   � ���������   �  ��������   �  ��������   �  ��������   �  ��������    �  ��������    ���������������������������������������������
  ����������ꫪ����� @����������ꫪ����*@U ���������ꫪ����
PU���������ꫪ�����GU���������ꫪ�����PU���������ꫪ�����[U���������ꫪ����0TUm���������ꫪ����0_UU����������ꫪ����0_UUÀ��������ꫪ����0�[�<���������ꫪ����0?�2���������ꫪ����0�����������ꫪ������U���������ꫪ�����V����������������;�f����*�����^C��:�O�������������Ԫ��P¾����������5����  ��먪�
j����{M���� A�)?���������{W���:@U�%�������(���_����:P�&�����������媪�:P��%�����������媪�P�������
h*
���w������������� �����w�^�����)�����`�����w�W��+��ʪ����������W�ի�����R��"�����Z����+�^�J���
�����V���0?��1��*�������귥����/��Ŭ��U�� ����W���� 
>�Ǭ��T��"����W����
~������( ���ꧾ��: �\����(�����ꫯ��:
�q���%� ����ꫫ����
8�Ǩ�*e� �������������W��j�� �������� ���q��*������꿪* TU�����j�������ꫪ
��W���W��j�j
����ꫪ����W��Ū*��
�����* @����?�Ū���*�����
����:�ű���Z*����ꫢ�����U����j�����ꫢ������_�����Z�����ꫮ��O��>|����jŪ���ꫮ�?�>�>�W̪��Z�����꫾�T�S��^ݪ���������O�?U��V{1����������*U�R���_�q����{������U�T���[�q��z�������zUU�Z�?m�Ŭ�z뮻����^Y������UŬ���媪��^V�Z����[��������WUU���[k]�����z����WUV񫵯o�U�����뮪���UeUUi����V����ﻪ���UYU�����VV���޾_檪�{UUU�����ZV�����Vڪ��{UU�ꪪ��ZU�����U����kU�������eU���z�[i���_U�鮪���iVŪ�z�n����_U������:�UŪ�j�[����_�������:�fŪ����U�ꯪ������:�VŪ����Uj�����������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?�<<����?�?��3�                  ��    ��  ������������������������ ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                            �              �              �              �              �              0              0              0              00              0              �              �              �            �             �              �              0  <            <  0              �              �          �             �    <          <    �              �        �     ?        �      �              �      �       ?      �        �?    �         �?��?           ���?            ���?           �?��?         �?    �        ?      �       �      �      �              ?        �     �        �    �              <          <              �   �          �  �              0              <            <              0              �              � �            ��              �              0              0                            0              0              0              0              �              �              �              �              ����������������������������������:������������������������������������""""""""""ʣ�����������""""""""""ʣ����������ꫪ����������#          �+          �#          �          �          �          �          �          �          �          �          �          �          �������������#""""""""""⋈����������#""""""""""⋈����������#""""""""""⋈����������������������#""""""""""⋈����������#""""""""""⋈����������#""""""""""⋈����������#""""""""""⋈����������#""""""""""⋈����������#""""""""""⋈����������#""""""""""⋈����������#""""""""""������������� �  �?  �?  �?  �  < ��� � 0�0 ��  ��  3  �3  �?  �   �   �?  ��  ��  ��  �?  <0  ��� �� ��  ��  �0  �3  �3   ?   ?  �  �?  �?  �< �33 0< <�� � �3 �� ��  �  �  0  �  �  �  �?  �?  �<  <�  <��� ������0  �?  ��  <�   3   �   �  �?  ��   �  ��  0�   0 �0 ��� ��� ��� �� <<� ����� ��?   <   �  � �� �� �� �� �?  � 0 � ���  �?    �  0  �  �  �  �  ?     � � �� 63 
� �� ?<< ��3  �  �  �  �?  ��  �� �? �? �? ��; 3 0 ?  �� ��  ��  �>  0  �  �?  �  �  �?  �?  �?  � ��� 0  0  ���� �?< �  �    �  �  �?  ��  0�  ��  0�  0� �<00 ��� ���� ���  �?  �  �  �?  �   �  �  �  �  3 ? ��  ?�� 0����  � ��  0<  �  �   �  �  ?     � <� # � � � �� �?  ��   �   �  � �  �  �  �?  �0  ��  ��  ��  ��  �� ��30���0 ��� ��� �?�<   �<  ��  ���0���������3 ?0< � 0�� 0�� ��? �� �         �? ��� ��� 3� <� ��  ?� �?������0�  �<  �  ?        �� �?������ �?<  3 ��� 0 ���0?�0��?3    <?  ��   �       <  <?  �??�3���?�?<� �00 �3 �3 �? �33  �         ?� ��? ?�? Ã?00����� �  ��  ��  ��  ��  ?  �  �  �  �       � �� <� �0 0 ��0 3<��?��� <�  �0  �3   �   �  �  �?   �   � ��� ��0 ��� ��� ������0 ?��?0 ��0 ��  �?  �?      ?   �   �    � �?������3�� ?�?��  0 ��  ��   � �  �  �   �   � �? � ����������?�� ��3? �� �  �          ����������?��? ��  �  ��  �����0��<�?��?               ��? ��? ��0 ��3 0� �� � ��< �� ����?<� �?   �?  �� �� ��< ��0 ?0 < < � �  ��  � �< ��0  �  ��          � �� 0� <�� �� �� < < �  �� ��? 0<  ��  ?                   �   � �� �� ��8 �� ��� ��� *�� ����  �� ��?  �?          ?  ��  �� 0* ,� ��: ��� .�� �ꨀ��00�� �? �   ��  �� �� �  �0  ?    3    �  �  �3  �0  �:  �?  �?  �  �?  <? �< << �0 �3 < 0 �?0  �?  �?  �?  0  �:  �?  �?  �? ��� ���  ��  �  0�  00  ��  0�  ��  ��  ��  ?  �  �  �  �  �3  �<  <0 <�< �� ���  < � �3  �?  �?  0  �  �  �           ?  ��  �� 0�> 0�� ��� �0 � �����? ?� ?�  �               �   � �� � ��  �? 0 � ��� �� ��  ?�  ��     �?  ��  ��  ��  �?  <0  �������� ��  ��  �0  �3  �3   ?   ?  �  �?  �?  �?  �  < ��� ������ ��  ��  3  �3  �?  �   �   �  �:  �:  �8 �33 �< ��� ̪���� �� ��  �  �  0  �  �  �  �?  �?  �<  <�  ������������:  �?  ��  <�   3   �   �  �?  ��   �  ��  0�   � ί: ��� �� ��� �� <<� ����� ���   <   �  � �� �� �� �� �? ��� ��� ���  �?    �  0  �  �  �  �  +     � ��� �� 6�; 
� �� ?<0 ��3  �  �  �  �?  ��  �� �* �* �
? ��; ��: �� �� ��  ��  �:  0  �  �?  �  �  �:  �:  �:  � ��� ����������� �?< �  �    �  �  �?  ��  0�  ��  0�  0� ��>0���������� ���  �?  �  �  �?  �   �  �  �  �  3 ? ��* ��� ������  � ��  0<  �  �   �  �  +     � �� ����� � �� �?  ��   �   �  � �  �  �  �:  �0  ��  ��  ��  ��  ����������: ��� ��� �?�<   �<  ��  ���0���������? �:8 �� ��� ��� ��: �� �         �? ��� ��� ?� <� ��  ������������0�  �<  �  ?        �� �?������ �*<  ? ��� �����0��0��?3    <?  ��   �       <  <?  �??�3����?��>,�� ��: �� �� ��? �3  �         ?� �: ��: ���?��ʰ������  ��  ��  ��  ��  ?  �  �  �  �       � �� ,� �0 0 ����3���?��� <�  �0  �3   �   �  �  �?   �   � ��� ��0 ��� ��� ��������?��?0 ��0 ��  �?  �?      ?   �   �    � �:��������� ����� ��: ��  ��   � �  �  �   �   � �: � ����������?�����3? �� �  �  �?  �� �� ��> 3�: ��: ��> ��  ��  � �< ��0  �  ��          � � 0� ��� ��� ��� ��> �� �� ��? 0<  ��  ?               <   �  �  � 0��   0� ��? ��? ��� �� �0< ��?@ �?      <   �  �  �� �?�  0��0 ?�0 �� �� �?�0�<? �? �  �� ��?��� ��: �� ��  � �� �� �� �� ��  ?  �  �  �  �  �?  <? �< �< �: ��; ��: ��:  �?  �?  �?  0  �:  �?  �?  � ��? �� � � �� ��  �� �� �� �� 0� 0�  �  �?  �?  �  �3  �<  <0 <�> �� ��� ��> �� �;  �?  �?  0  �  �  �           ?  ��  �� 0�> 0�� ��� �: �������? ?� ?�  �               �   � �� � �� � �� ��� ��� �� ��  ?�  ��      ��<<�      �<?3�<�<�      ����    H�Z��� �ܩ �Q��T��U� �G���E�E�;�G�: 8��E�r� Y��E���H���F�E�E�;�G�:� �Q��U 8��F�F�F�;�H�:��U��Q 8��F�D� Y�L�� Y� Y��E�;��U�G�:� �Q K��Gi�G�: 8��H�:��Q K��H8��H�: 8��H�� Y�L뛩��� ��d�(�(��z�h`�Q
��d���d�� ��`H� � 8����h`H��(�(��h`��x� �� ���4��� � H� � l�d d! :�`� ����:����;� ������`���F�;�a�Ld4�  ��� 
��4�4����T ��  � 
� 
����
�����@�ҩ
�:���� �� � �ߩ�����
���Z�;����F�;�
�: ��d4L�����4`� �����:����;� �� �ߩ������:����;� �������`���K�;�a�L �������L���L革�:���� �� � �ߩ�����
���s�;���
���K�;����_�;��: �߀���:���� �� � �ߩ�����
���_�;����
���s�;�é��K�;��`������:����;� �� �ߩ������:����;� ������ֹ���:����;� �ߩ�� 0�`�Z�

�� �ɠ�M ����� ��z�`ڥi�����:����;�  V��:�:�����`H ؅4��L��ɿ���������詃�� ��� ����Lm� 0� K�������������<��� 0� ؅4��	����L�ɿ���������⩃�� ��� ����L��h` 0����$�4������������L9���L6���������$�4������������L9���L6���������$�4������������L9���L6���������$�4������������L9���L6���������$�4������������L9���L6���������$�4������������L9���L6���������$�4������������L9���L6�������4������������L9���L6������� 0�` �ܩ�;��:�i �ߩ<�;��:�i �ߩF�;��:� �ߩP�;��:�i �ߩn�;��:�&�L �ߩ�:�  �ߩ�:�! �� ��`FZxK_s7Pi�55NNgg��    3HBP3�BLH[PL�[eHtPe�t~H�P~��H�Z�3� � �� ۡ�0 ��1 �L��� ���	���=��Z0s�qɂm�k���� �� ��1 ��X �� ۡ�1 ��K ۡ š�C��Z06�4ɂ0�.��0�� ۡ š�0 �� �� �� �� ۡ�0 �� �� ۡ ��z�h`��  ����0�`��3��5��M�	8�M� ������`��5�
��P��d����`�� ���� ���� ���� ���3�0
��P��d`��3���P�d��	��`�'i�Q�i ��"A�Q��
�������P��dL���Q��7���P��d�'��P�d��Q��
�������P��d�	�� � ��` ��.���s�����l���#D�'�'�
�������P��dL��'8�'�8���P��d�(��P�d��'�'�
�������P��d`Hڢ����P��d�:��60��P��d�'�'����P��d��'8��0
���P�d��	Ю�	�����.0���'�
����(0
���P �΢ �����.0���'8���� 0��P ���h`�P�2i�	08��P������������
������d`� �.�3�7�3�3�8��8���'8�'	��'8�'�	� ͣ���.`H�Z��Bd>d?�
�6�H�7��0��1��4�5�2�3����xd'd(d)d*d���������d d!������z�h`�����������Ώ� ��`Hd&�&�P��h`���.dN�.��� {���� 뤩 �.�N�N�
0� �!��L�� ��d>d?��@�=�(�A��:��;�R�< +�dC���D�:�E�F ܩ�B�@�<���:��0�;�' O���:��t�;� c���<��:�l�; O� ������ ��  �) ��dB��<��:�l�; O���B�)����)�������"e&mm�m�)������ �L'� 
� 
� 
ۭ�:��; c��8���;���m��: c���<��:�'�; O������<���m��:�'�; O��L��  �  �  ۭ���� i� �"i�"�  � :�`Hd>d?��=�@��A +�h`Hd>d?��=�@��A�F�< +�h` ��d>d?��@�=�(�A��:�n�;�S�< +�dC���D�}�E�F ܩ�B� �<���:��d�;�' O���:��4�;� c��*�<��:�&�; O� �� ������ �� ���#e&me(m�)����dB�0�<��:�&�; O���B���� �L�� 
� 
� 
ۭ�:��; c��i��;���m��: c��  ����O�)�� ��)��������<��:�'�; O������<���m��:�'�; O��L'�  �  �  ۭ��0�����!i�!�#i�#�  � :�`�  /01/>@?@!!                                                                                                                                                                                                         ����          ���)  jffffff   `fffff� ��������������������fffffffffffffffff�
������������������i*����������������������������������������IDDDDDDDDDDDDDDDDd�J$�aDDDDDDDDDDDDDDDDH�J$�aDDDDDDDDDDDDDDDDH�J$�aDDDDDDDDDDDDDDDDH�J$�*aDDDDDDDDDDDDDDDDH�h�����������������)(�����������������O(h                0)(                p(h                0)(                p(�                �*�                �
�                �
�                �
�                �
�                �
�                  
�                  
���������������������������������������FDDDDDDDDDDDDDDDD����FDDDDDDDDDDDDDDDD����FDDDDDDDDDDDDDDDD����������
����FDDD����
�EDDDDDD����JDDDDDD
��
�EDDDDDDDDDDDDDDDDD
��
�EDDDDDDDDDDDDDDDDD
��
�EDDDDDDDDDDDDDDDDD*h�)�EDDDDDDDDDDDDDDDDD*h�)�EDDDDDDDDDDDDDDDDD*h�)�EDDDDDDDDDDDDDDDDD*h�)�EDDDDDDDDDDDDDDDDD&()fDDDDDDDDDDDDDDDDDD��FDDDDDDDDDDDDDDDDDD�����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ���ة��  ��� � � � � �ύ& ��" � t ���d���� � �������� ��XL��H�Z�&�'��'�(��(�)��)�*��*z�h@H�Z�' )������ �� ���# �$ �% (z�hX@����2��#  �� }� g� ��d� i� ��� �� ]� a� �� h��4���� �� E� G�L�ǩN�<�  B��(�=��@� �A��B� �]�����:�>�]�;�? +ۭ    ���.��  �  � ���0"�]�;�?ʽ]�:�> +ۭ    ���ʀ� �ܩύ& `Hڪ�)�




�M��)M�& �h` ��d>d?��@�=�P�A��:�7�;�P�<� B� +۩ύ& ��:�<�;� �� �� �� :����3d d!L��L�� �ܩ�� i��:�<�;� �ߩ�:�P�;� �� ���<� �!0��̩�:���;� �߭�����:���;� �� �� �������� �ܠ	����:����;� ����0������ K���� K��� 0��� 0� ح���L�� �ܩ�� i�d>d?��@�=�C�A�
�:��;�Q�<� B� +۩ύ& ��:�x�;�  �ߩ�:���;�! �߭  ��� ��L��  ۩ �� ]� a� �꜎��
���Ņ�ƅ�&ƅ��Ņ�ƅ�&ƅ���@ƅ6�Mƅ7�Zƍ�gƍ���	���0%� ����'��d� �P��
�箍�tƅ3�R������'��d� �P���	�� ����'��d� �P�	����'��d� �P����ƅ3 l� �� Z� n� �ԩF� �˭��L�Į  ���� ����L���� P؀�����)0�݊)p�؊)`�ӊ) ��� �� ���3����)*��L:Ċ))��L:Ċ)&��L:Ċ)%��L:Ċ)(��L:Ċ)$��L:Ċ)"���
�)!�L�é�P������������E�;��� �Φ3�d
��0��;����; �Ԝ��������� �� �˩�� i�  �L�� �� �� ֤3�������L:����L:����L:���L:��	��L:��
��L:����L:ĩL:� �ܭ��� ��!i�!�#i�#ة����3������ i� �"i�"ة����3���������� i�d>d?��@�=�P�A�
�:�7�;�O�<� B� +۩ύ& ��:�#�;� �� �� �� :�  ۭ�
���Ņ�ƅ�&ƅ��Ņ�ƅ�&ƅ���@ƅ6�Mƅ7�Zƍ�gƍ� ����'��d� �P��
�� �� ]� a� ��L�ÎƎƬ������$�B�`�~ǜǺ��ǘƘƶ������.�L�jǈǦ����ǢƢ��������8�V�tǒǰ�����     



  p��p   (hHH   6::6& >��̆>7�ol   
!�@0@`dP0&
  Ȉr�����t
  ���������
8." �Ȫ������
8* (Ȉx�����p
8(($�@0TPxhF8
8$,0(� @HP 8(   (� 0(8 ( ,�`H�p�`P0
$,( Ȩ`�f�xHX
&"(�px��hh^J
"($,�hh��X^@0
L�� hץ����
���� ��L[� �� �� l� �ѭx� �ҭx� �ܜx Z݀ �� � nɦ3� �� � ����
���2���y��� �� � ��������5�P��Z� �P�E�O�;�E �� �� ,ץ3�2�5�4 �� A� Z� 7Э�� ����3��5�  ��� ����L�� �� �ץ+���� �� ֢ �E�;��
�������� �� �� ,׮  ��� �� �� �ץ+���� �ѭ��L�ĭ���	���� ��L��L�Ǧ3� �#�	�� �- Hͥ-��� �ͥ-��� �˥-��� �`� �P
��]�}��ȹ]�}'�1�'��
�ۢ �d
��0��;ȹ�E����;ȹ��E��
��`H�Z �ʭ
��3� �L�ʽ��L����h���ȹ������������ �3��� ���L��m �ȱm�ȱm �ȱm�ȱ��Ȍ�L����8�o�m�yo�ȹo�m�yo��F������0HL�ɹo�m��ȹo�m������#���� ���� �����z�h`HZ���L�ˤ3� ���P��L�����i� �'i�L������$��+�'i��8�� L�˹'i���'i������� �'i�L�������'i��i� ��'i���'i���zh`H�d>d?��=�@��A� ݭ #ݭ�< �� +��h`HZ�:�b�;�m�����x��d�
 ��zh`H��T��U�b�:�m�;��d ��h`Hڦ0�2� ���1�4���F�LEͽP�LE����8�'0^�Z�8��0O�KL2����8�'0;�7�8��0,�(L2���$�8�'�0��8��0�L2�LE���!�8�'�0���8��0���L2���$�8�'�0��	ŭ8��0���L2�LE���!�8�'�0���8��0���L2���!�8�'�0��ŭ8��0���L2ͭ8�'0����8��0�������3 �Ω�����-�h`Hڦ0�2� ���1���L�ͭ�H�L�ͭ8�0)�%���!����P���8�'�0��L�ͽP����'8�0������3 �Ω��-�h`Hڦ0�2� ���1���L�έ�H�L�έ����(�P�U�8��0J�F�'8��;��07L������/�P����!�8���0��'8����0L��L������,�P�����8��0��ۭ8�'����0�L������%�P�0�8��0��8�'��0�0L�Ω���3 �Ω��-�h`�Z� ��	���


}P�����d���


}P����Νdz�`HZ�2� �"��H�����A�4�y��F��� ��L�Ϡ �8���0&�"�8�'0����3  �  �L�� ��L����
-L4Ϥ0�2��1�8���0��8�'0��0���zh`��F�L���G��C� �2�8�8���0-�)�8�'��0��3�2� �����������
п`�3� �8���0$� �'8�'�0����'НP�/Нd���0�`�3� ��L�� �ϥ3�2����ﭑ����㜑��3��3�	�Թ'8�'P��	0�3��8�'0�� ������J��J��J�S������������<�����0%�$0����������������P �Μ�`���>�3� ��6�1��0��0�8��8���'8�'	��'8�'��3`�	�8���0��8�'0
����3`��2����0 5Ѧ3�	�"�	 � ��.ɨ0*�(�3��0 �  � ���	������
�
�����`���3� �C�	�?������H�1��0*�#&�0�0�0�8��0��0	�����`HZ�x���/�8�<���F�а[�8�70��L�ҭ8�60��b�L�ҭ�p���E��A��p���4��0�3��	�&�������3�0�
���������3��L�ҥ88�0���L�ҩL�ҥ98�0�'�8�60���L�ҥ88�0���L�ҩL�ҭ8�60���L�ҥ88�0����xzh`Hڦ3� �L�ӽ��L�Ӯx���7�L���7�7L�����7��6�L���6L�ӥ6���6�7�7L�����6��L����&�6��9���L���7�7L�ӥ9���L6��6�7�7L����	�9����L����&�9����8�<�L���6L�ӥ8�<�Ld��6�7�7L����	�8�<��L�ӥ6�	�8�<�L�ӥ8�<�L ��7�7�6L�� �Ӏ�x�h`Hڦ3�����(�M��N��O��P���M��N��O�
�P�x���78�M��7L��d7L�����78�N��7�68�O�	�6L��d7��d6L�����68�P���6L�����7eNɐ��7�ʩ��7�����7eMɐ��7L�ԩ��7L����!�7eNɐ��7�6eO���6L�ԩ���������6eP����78�N��d7���h`Zک�WdV� ������
����  ����
0�z`Hd>d?��=�@��A��Ci�D�'�Ei�F�C�6��8��8�D�8�C��@�L�եD�6��8�6��@�6�C�8�@�>�E�7��9�ۥ9�F�8�E�3
�A��F�7��8�7�#
�A�7�E�8�A�?�C ݥE #ݹ;�< �� +�h`H�Z� �� �:�X �;�c �A�n �@�y �V��W� �եViP�V�Wi �Wz�h`�X �D�c �EdOdC� ڦE�V�����Z�D��C��Cz�O�O�y ��D��dO�X �D�E��n ��`H�Z�	�� ���,�V8�P�V�W� �W�X �:�c �;�y �T�n �U�V��W� �ֈ����z�h`�
�D�(�E��� �dOdC� �E�V�����D��C��C�C�(��i(��i �dC�O�O���D��dO�
�D�E��м`��� ��
�:�(�;��T��U ��`H�Z�;�N�:�DdOdC� �;�V�����C�%�D��C�C�(��i(��i �dC�O�O�T��D��dO�:�D�;��Uк�N�;z�h`H�'���'� �+�(���(� �,h`d$�7�)�����%�����%���%`�*���*�%��$����� ��)�!�7�)��$�8��$��%��%�Y�$������`�
�:�(�;� �ߥ% �ߩc�L �ߥ$ �ߩ
�:�2�;� �ߥ  �ߩc�L �ߥ! ��`Hڢ��'��+�(��,�h`H�Z�5�)�� P�LL؊) � ��LL؊)� �LLحO�E�)� ��LL؊)� ��LL؊)� �LL؊)� #�z�h`H�Z V� �ש�)��&  �� 
ۭ  )��� �� 
۩ύ&  ��z�h`�  ���� ��  � 
�`�3� �L��0�������
�������)*��L�؊))��L�؊)&��L�؊)%��L�؊)(��L�؊)$��L�؊)"����)!�
��P�� ��`�3� ��0�5L������������I����)��Lxي)��Lxي)��Lxي)��Lxي)��Lxي)��Lxي)����)�
��P�� ��`�I�����P��)	�	��P��
�)
���P� ��'ɠ	�� �P�
�� �΀�d`�I���	��P���)�	��P���)���P�� ��'ɠ	�� �P�
�� �΀�d`��P��d� ��� ��`��P��d� ��� ��`�8��8��T ,ݥE�M�F�N�'8��8�'���T ,ݥEeM�M�NeF�N��MdN`HZ� �/��U� �2��/� �ڥ/�0�
�U��/��2��/� �ڥ/�1zh` 7ڥM�O�N�P��2�# 7ڥN8�P��M8�O��/�N�P�M�O���0���U��`H�  ����h`Hd&�  ����&�0�h`H�Z�/���� ���� ��z�h`Hd&�&�
0�h`H�Z�<
����轁��?� ��e=��i ����e>��i �� ��@��;� ��i0��i ����e:��i �� � ڱ�B� ���1�
���Q���@�����A��i0��i ��e=��i ���z�h`H�M�C�D�N�E�P�F ܥM�C�O�D�N�E�F ܥO�C�D�N�E�P�F ܥM�C�O�D�P�E�F �h`H�Z�C�D��E�F��F�K�E�JL�ܥE�K�F�JL�ܥC�D��C�J�D�KL\ܥD�J�C�K�K�J�K�L��)� ���IL������IL�����0�IL�ܢ��I�E�V�����JJJ��EI��JL^��K�J�K�L�ܥC)� ���IL������IL�����0�IL�ܢ��I�J�V�����CJJ��EI��JL��z�h`H�Zd�@�� � � ��������z�h`H8�6�:h`H8�7
�;h`HڥT
�EdF�TJ���T�� � �eEH�Fi �Fh�� ���E�h`H l� }� �� �� \�h`H�6i(�8�7iP�9h`�Z� ����7�
�����L���9��E�
����Cȹ��D�6�C��C�8�D��D�C ݥ:

�C�E #ݥ;�E�F�D ݥ:

�D �L��z�`�Z� ����6�
�����LY��8��C�
��7�X����Eȹ��F����Eȹ��F�7�E��F�ŅE�9�F��E���F�C ݥ:

�C�D�E #ݥ;�E�F #ݥ;�F �L��z�`�Z� �����������L�ީ�<���E���F�7�E02�0�FͰ�8�E
�?�F8�7
�A�7�E� ݥE #ݩ�=�@ +�d?Lbޥ9�E0��F0
�� �Ad?��8�E
�A��Lb�z�`�7�=�;�&�$��E��A��<��=�@� ݥE #� +�d?LU߅E8��?�8�7
�A���|0��9��0�����0���Ad?�̅E��<L��8��
�A��`H�Z�'�-��U���Q�;�V�����:�Q��i��i �ȲQ��i��i ���Q��z�h`H�Z
������ ��$��b��a��'�8�7�L �� 
�Ȁ�z�h`H�Z�)�JJJJ�L �ߊ)�L ��z�h`H�Z�L�a��$��b��%��'��'��c��&��-��U���M�;�V�����:�%��Ȳ%����M���:�:z�h` 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P�� P�� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____________MODEbbSELECT$babEXERCISE$bbbCHAMPION$bPUSHbSTART$TIMEbSELECT$bbabTHREE$bbbbFIVE$bbbbEIGHT$bbTEAMbSELECT$SPAINbbbRUSSIAN$ITALYbbbHOLLAND$FRANCEbbENGLAND$SWEDENbbGERMANY$bbSPAIN$RUSSIAN$bbITALY$HOLLAND$bFRANCE$ENGLAND$bSWEDEN$GERMANY$VS$EXERCISE$CHAMPION$TIMEbb$SCOREb$YOUbLOST$TRYbAGAIN$YOUbWIN$TRYbNEXTbTEAM$HAbbIbKICKbIN$TIMEbOUT$WEbARE$THEbCHAMPION$�������������
��"�2�B�R�b�j�r�z������������������������          @ ` ���� � ` @     @```@@� 8p���8(080(8(08�8  8�Ш����Ш����8H`pp����������/�I�c�}�� � �F � �G � �H � �G � �F�����F����G����H����G����F�����F����G����H����G��� F���F�	�G��H��G��F�  F  G  H   G $ (F�F	G
HGF���F��G
��H��G� F���F��G�
�H��G��F�	
  	
  !!"###$%%%JJKK  &'()*+,-..//00112233445566778899::;;<D==>>??@@AABCCCDEEELLMM   ���� �  �   ���� �  ���x�w�w�w�����������7�w�7�w�����7�w�����7�w�����7�w�����7�w�����7�w�����7�w�7�w�7�w���������7�w�����7�w�����7�w�����7�w�7�w�����7�w�����7�w�7�G�@�W��������� � �@�@����  0@P`p��������  0@P`p��������  0@P`p����������������������������������������� ������ ]� a� � � � � � � � �* d�dܜ ����d�`�������� ]ꥱ� ���  ��渥�ų� �祑������ a꥾� ���  
��ť���� 襏���J�������� ]꥕� ���  饑������ aꥣ� ���  d�朥�ŗ� [�檥�ť� |����� o� ��`������ȱ���ȱ���ȱ���ȱ���)
������􅛥�)0��ȥ���������Ȅ�d�d���� �L褞 ��� �
��� �d���Ȅ�d���������ȱ���ȱ���ȱ���ȱ���)
������􅷥�)0��ȱ������Ȅ�d�d���� �� ��� ��)��	����d� �`������ȱ���ȱ���ȱ���ȱ���)
��������ĥ�)0��ȱ������Ȅ�d�dƥ�� к� ��� ��)��@Ы����d� �瀠������ȱ���ȱ���ȱ���ȱ���)
������􅩥�)0��ȥ���������Ȅ�d�d���� е�� ��� �
��� �d���Ȅ�d�����
������ٱ؅�ȱ؅�`��
�����轉�ٱ؅�ȱ؅�`H�Z��)?	@�Ȥ�;��%ȅȤ������)@��J��ȅȥ��8������)0��Ȅ������Ɲ��d��ȍ z�h`H�Z��)?	@�Ȥ�;��%ȅȤ������)@��J��ȅȥ��8������)0��Ȅ������ƫ��d��ȍ z�h`H�Z��)?	@�Ȥ�;��%ȅȤ������)@��J��ȅȥ��8������)0��Ȅ������ƹ��d��ȍ z�h`H�Z��)?	@�Ȥ�;��%ȅȤƱê��)@��J��ȅȥ��8��ǀ��)0��ȄƱ�����ƥ�dƥȍ z�h`� `� `�թ��� o�`H�Z������֩��Յܥ�)?
�����轐��d� ��z�h`dܜ* d�`�ݱޅ�ȱޅ�ȱޅ�ȱޅ�)
��������Υ�)0��Ȅ�d�dϥ�� ��d�`H�Z�����Le�ʅӥ�;��)��Ӥϱͪ��)@��J��Ӆӥ��8��Ҁ��)0��Ȅϱ�����ϥ�dϥ�)�ȥ�)����
�@����ȅȥӍ( ������* ���̥���� ��z�h`H�Z�  ��  ��d�d������ [� |� � d� o����z�h`H�Z��� ���� �dۥ�)?�ېD�� �>��
���􅯽����􅰽��d�d�� ������)������ ������ �� o�z�h` �2�� �2�� �2�� �2��.2�� �2�� �2��.2��.2��}2��.2��}d��}2�� �2��.2��.2��}2�� �2��.2��.2�� �2�� �2�� �2�� �d��     ��2�}2�}2��2�\2��2��2�\2�\2��2�\2��d��2�}2�\2�\2��2��2�\2�\2��2��2�}2��d�     � �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D �2�D 2�D �2�D 2�D 2�D     � d2�D w2�D d2�D w2�D K2�D w2�D K2�D w2�D _2�D q2�D _2�D q2�D q2�D �2�D q2�D �2�D T2�D q2�D T2�D q2�D C2�D T2�D C2�D 2�D     �O2���2��h2���2�\2���2��h2���2�O2���2��T2���2��2���2��T2���2��2���2��}2���2��2���2���2���2�     ��2���2���2���2�\2���2���2���2�O2���2��}2���2�\2���2��}2���2�O2���2��2���2��2���2��2���2�     �O2��2�h2��2�\2��2�h2��2�O2��2�T2��2��2��2�T2��2��2��2�}2��2��2��2��2��2�     ��2��2��2��2�\2��2��2��2�O2��2�}2��2�\2��2�}2��2�O2��2�2��2��2��2�2��2�     � 2�� 2�� 2�� 2�� q2�� q2�� q2�� q2�� d2�� d2�� d2�� d2�� T2�� T2�� T2�� d2�� ?d��     �\2���2��\2���2��:2���2��:2���2���2���2���2���2���2���2���2���2���d��     � ��� ��� ��� ��� �2�� �2�� �2�� �2�� �2�� �2�� d2�� 2�� �2�� d2�� 2�� �2�� ?2�� T2�� d2�� ?2�� T2�� d2�� ?ȧ�     ��d��d�Td� �d�T2��2��2��2��d�}d�     � ��� ��� ��� ��� ��� ��� ��� �� q�� d�� _�� T�� K2�� T2�� ?d�� 2�� 2�� ?2�� 2�� 2�� 2�� ?2�� 2�� �� q�� d2�� _�� T�� K2�� 2�� ?2�� q2�� d2�� _d��     ��2��2�}d�     � �
�� /d��     � ��     � ��     � _ȧ �     � ȧ �     � ���� _���     �����������  �O
   �O
   �o
   �
      d
   �
      �J   �J      �   �     ( �
     ( �
    	

			�

		�
	�
�
	

�
	
	 ������������������������  ����  |��|�|�$��  |��|�|�P���  ��  �  ��  �  R�  $�  <�N�r�~�<�Z�f�~���?�J�Y�h�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           F� �g�