                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�   % UU%        VUeUUVUe          Ve        UVUeVUeU           	 % � VY	e%�UVVYYee��VVYYee   V Ye�VVYYee��VVYYee��VV � X�UXU        U�UY�UYU         @ T@�TY        �UYUU�UY           � ` X V��`eXYUV��eeYYVV��eeYY @ P T �@ePYTV��eeYYVV��eeYYVV��   0      0      �0      33    �����     �;   �������?< �:<    <    (��(??���?������������������������������UUUT���?�?�?�?�?�?�?�?�?�5�5�5TTPP� ������wwwUUT T <������UUUU???7��?_���_��?����=�=���__�� ��� <�<??      T��T       @   P  P  �  � T�U�~T� �  �  P  P  @           @U   @Y   ��  �� P��_T��_���T��_P��_ ��  ��  @U   @Y                T    U   e  @�  ��  �� P���T���U����YT���UP��� ��  ��  @�   U   e   T                 ��?              �� � �*� � �        �� ��?� � �?    �         �         �         �         �         �         �        �        �
       ���?       �>    ���������� ����0     ��        <<                                        .        .       ��      ����     ��   ��������? �3���    ��                                   ��?     .   ������� ���33    �                    �,?   �  ����� 3��         ����?      �         �         �         �         �         �         �        0      �?��     ��   ��������� �γ��0    ��       �        �                                                        3      �?�     ��   ��������? �3���    ��       ?                                     3    ����    ��   ������? ����    ?     0    0    0    0   �3?   �  ����� 3�3  �   �             �      0                �  0 �0   � 0�        ��     ̯    ��    0�     ��    ���    0�?    �     �      0      �           �     0                      �    0          � �0  00�  ��  ��  ��  ��   ��   �   0        3   �    0                  �    0    �    �  �<   0?   �0   �   �          �   0    �                    0      �            � �   0 0   �0     �     <�     ��     ;�     0     �<    �    ��0     <�            0      �            �      0      �               0    �    0� �  0  3  ��  �  �3   �   �3   ��        0    �        �    0    �        0    �     �  ��   �<   �3   0�   �<   ?    �        �    0    �             � � 3  ��  ,  �  � ��  0  �   0                    0      �             �   3 0   �0    0�     ��     �     ��     �?     ��    �:    ��0     �            3      �      0            0      �               0    �    0� 0    3  ��   ��   ��   ;   �0            3    �    0        0      0  �0 03  �  �  �  �3   �   0   �                  �      0               �   0 �0  � 0    3    ��     �?     ��     ��    ��    ��    0�        �      0           3     �      0                      0           �  �0 0  03  ��   ��   ��   ;   �   0        3   �    0            @ � YT� �
�*�J�����f��"�IZP��U �@�� @�j  ��j	 QTR	 QUV� UV�UV�"UE�T!��%U�VQT(Y��H Z�j ��U D      ��V ����P��V�iVA�e�
X��YE�*��
��Ui��RU ( V@ ��R (e ��� ���Q@����U�je�j*d	�Z��JDVR �VYV�� PU   T     dU    PU�	   P    T�*U �U��VU d����U �Z��VV��iVU��e�
��Y��YU��*���$��Ui���RU ��%V@ �Q�R (e�� ��D�� ��T�U@��T��U�jUe�jjhe��ZV P���JT�fVR Z  �VYV  ���  ��V�  XfUU    AU    TU     �     ��    P��	  @P�   @ �  �VU� �F��
 ��
��* h���  X����� X��T( Z��A` (PB�eV% ��	� @�j
�Z@U"�T @TU
�U  DU)�U D�&�U�HU�UfUHf*hf	DU)P�UUZ	�FV�iZ
 ���Z�
@�f��@J�J @Y�PU*  �V��
   � * ����;  ���? ������ �   �� � ��� ������
��� �   ��  ���� �� ����������*��������  �    ���   ������ ���   ���*  �����? ������ ������������誫����믿�� �
 ��
��ww����* �� w������_���_www_���_���*  ���*  ���  333��*�����33333�����33333����������  �����  ����z  ����_���<��\���������<��<�s�������<��<�s������� ������   �����z   �����^   �����_       \��������ܪ��    ���z��������_       \��������\       \��������_       \��������\       � ��������?  �  ���������� � ��� �>���������  �   ��  ���� �����������������������   �    <�    ��  �����? ����������������������������������                               @                   �   �                      � �                            ���  ���                     �         �@             @   �            �                            �      �      �     �     �     �   � �@   � �   �     �    ��     ��                 �*  ��
                           � �         �    �   �@� �    �@  �     �    �      �     �      �      �           ������������������������������������������������������������������������������������ ��0���������������������������������������?��                        �������������?��                        �������� ��0��                        �������������?��                        �������������?��                        �����������0 ���������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU    @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU UUUUUUUUUU��������������������UUUUUUUUUUUUUUU������������������������������UUUUU����������������������������������������������������������������������������������������������ZUUUUUUUUUU��������������������������������������������������������������������������������Z�����������������������������������������������������������������������������������������������UUUUUUU�UUUU����������뿺~UUUU����������������j������������������~��������_���������������������������~��������_����������UUUU�����?  ���~UUUU����_�������������������   ����������������������������������     ��������������������������������~UUUVUU���������������������������    �      ������������    ����?� 0    �     @���3����0    ��??�����??    ��      @����<�<���?    ��?������??    ��     @��3�<�����?    ��?�� � ??    ��      @��3������0    ��?�����??    �;@UUVU@��3���?���?    ��?������??    �;@    @����<�<���?    ��?���<� ??    �;@   @���3���0    �����������    �@    @�����������    ����������������@ TV @�������������������������������@ @ @�������������������������������@ C @�����������������U��U���UU����ȏ��������������������U��U���UU���@ C @�����������������U��U���UU���@ @ @�������������������������������@ TV @�������������������������������;@    @�������������������������������;@   @�������������������������������;@    @������������������������    ����@UUVU@�����         �������?    ����      @����?         ���������?    ����     @����?         ���������?    ���      @����?    <    ��������?    ���     �����?         ���������?    ���>      ����?         ���������?    ����WUUVUU�����?    <    ��������?    ��﫪�    ������?         ����������    ��뫪�? 𯪪����         ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������*�

(�*�*�*�*
(�*�*
(
(
(
 
 
(
(
(
 
 �*�*
(�*�*�*�*
(�*�*
 
(
( (
 
 
(
( (
 
 
(�*�*�*
 
(�*�*�*                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<3<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  ��<� ��<�<��   �� ��� �� �       ���        ������                ������       ������     ������            �?�?      PRESSaSTART$TOaPLAY$LEVELaSELECT$PRIMARY$MIDDLE$ADVANCED$MISSION$C$O$M$P$L$E$T$I$N$A$G$V$R$bbbbbbbbbb$baREWARDab$MISSIONaaCOMPLETE$BONUS$TOTAL$BANK$BEFOREHEADaCOMPLETE$eeeeeeeeeeheeeeeeeee$MUNITIONSafEQUIPMENT$eeeeeeeeeegeeeeeeeee$GUN$MISSILE$FUEL$FUELTANK$ARMOUR$SELF$GENETAL$ADVANCER$SPECIAL$SMALL$MEDIUM$BIG$LIGHT$HEAVY$eeeeeeeeeeieeeeeeeee$eeeeeeeeeeeeeeeeeeee$WIN$RESULT$dddddddd$COMPLETE$HITaFIGHTER$HITaTANK$HITaWARSHIP$APPRAISE$SCORE$ENTERaSIGNATURE$CONTINUE$END$COST$�����	���!�#�%�'�)�+�-�/�#�1�+�#�%�7�3�+�5�9�;�F�;�Q�c�t�c�i�o�������ǃ��˃��Ӄ��؃���#��8�����������M�Q�X�a�j�v��������bhn������
Tf	Qamy(
2222222222222222
22

&
.>JXdt� 
  " *2 :B JR Zb j r zFIRST$SECOND$THIRD$FOURTH$FIFTH$SIXTH$SEVENTH$EIGHTH$NINTH$������ÅʅЅօޅ�(0 P0daENEMYaaFIGHTERa$aaENEMYaaaTANKaa$aENEMYaaWARSHIPa$ORDNANCEaFACTORY$
��,�
��,�
�,�=�P�)�)�)P     000Hڭ���� ����� �
��녍� �녍�  g� �̩ 6��  ��[ �̩�� �2�� �d�� �  ���  ��= ������`��� �a��� ʽN��� �N���  g� �̭��� �	��� ���� ���h`Hڢ� 6� ������ �ũ�H *� �� ���h`H� �Ω� �ϩ�8� �� � �� �ԭ  ���� �� ��� �� �� ���h`Hڢ� 6� �� ������ �� �� �� ���h`H�Z��� ��� �: ����� ��� �; ����� �3�� �< ����� � ���$�� �8�X��  ����� �E�� �= ����� � ���� �� �ʀ��� �W�� �> ��� ��"�� �� ���� �i�� �? ��� ��"�� �� ���� �{�� �@ ����� �	8�mX�	��#�<�mm�����"�����P������m�����i
��  �� 툩�� ���� �A ����� � ���} �� �ʀ�  ��� �� �� `� ��z�h`H��������&8��������8����~i�~�i ��Э��8����~i �~�i ��⭄�8����~i0�~�i �����h`H�Z� ��  � #��|0N��~�{0D��}�z0:��y0P��~�x0F��}�w0<��v0J��~�u0@��}�t06��L � 6� V��^� �b��������- |��^� �n�������� � i��^� �h������� ��z�h`�w�z�x�{�y�|� �h�n����`�t�w�u�x�v�y� �b�h����`�}�t�~�u��v`�}�w�~�x��y`�}�z�~�{��|`H�Z��� �L���(�� ��� �B �� �� Ћ������ � �'��  �̭� H�a�� �����  ��h�� ���  ���' 9�������  �����  ���
 9��������� �'� y�LI��
�� LI������ �'� ��LI��#�� LI��� �� %��U %������  �� 9�L����� P������  ��� ��� P� ��L�����L�� P������  ������� P� ��L��z�h`��� �K�� �C ����� �d�� �D ����� �}�� �E ��`��� �K�� �v ���u ���t ����� �d�� �y ���x ���w ����� �}�� �| ���{ ���z ��`Z�
������ ȹ���� ���� �'�i7��^��z �� 9�`Z����
������ ȹ���� �����^�8�7��'�� z`H�Z8�7�� �� ͘ �� ��'�� h`H�A8�7�� �� ͘ �Ξ ��'�� h`H�Z��  �ϩ2�J  �� ͩР��������J �<��J ��J �m �m )�խ ��
 �ө�m �ĩ�� �N�� �9 ���  )��� �� �� ��z�h`H� �� �
�� �S�� ��� �/��  U�h`H�� � �  ҍ� �  �έ �\� ҍ� �  �έ  ��)LF����� �  ҍ�  �έ  ��� ɐ0�����  �Ω�� � � ҍ�  6�� 6� �h`H !�� 6�� 6�� 6�� 6�h`H� �ϭJ 8� �J ��� � �� �  I� ��� �h`Hڽ �	0� <��h`ڢ�m )�ɀ0 rӭ� � ��m )��m �
�� ��#���� �`Hک� � � X��	�� J�� I��h`H�Z� ��� ��� �a�� �� �� ���� ���  U� �̩ �� �� �� ���  UΠ��   ����V���!� � �� �� 8��� ���� �y�� ������� �� �� i�� ��� � ����8�� ���� УLp�� ���� � ����	������W���	����z�h`H�Z�
��N��� �N��� �
������ 轼���  g�z�h`� � � � � � � � � � � �( �) �* `Hڜt�u�v�w�x�y�z�{�|� �^�b�h�n����$�b�h�n�h`� � ��Y`�m�� � ��V� �	�
���0������8��;�7�0�<��B�?�C��U� �F�,���������}�~���� � �' �J �m ��#�� �� ����� �
�� ��X�W���`� �����!� �)�-�.�3�9�A�J�� �T�%���S�7��7���?���K��L�M�P�N�
�4��
�5��@���,�=�*�����/����+�����b��� �k��=�t��>�
������ ����� 轭��� ����� �!����
��=


m�6� �Z��[`H�Z�� 6� �� ������ �� �� �� �� ���"�� ��� � �� �̭  ��� ��z�h`H� �� �� �(�� ���� � ��  U�h`H���%��� �J�� �b��  ���i�� �	�
�p� �=��� �d�� �b��  ��� �	��>�
�=�G��
i`�
�i ���=���!�"��� �t�� �b��  ����mi�؀	�"� V�� ���h`H�Z��� ���� �b��  ���a�� � �������� � ��� Z�� �ʀ�z�h`Hک ���	 Z�� �ʀ��h`H�Z��
���N8�����
�8��
��� �t�� �a�� � ��������  ���i��i � V���������z�h`H�Z��)�JJJJ�� ����a�� ���� ���)�� ������a�� ���� ��z�h`H�Z��)�JJJJ�� ������� ���)�� ��������� ��z�h`H�Z�)�JJJJ��  ���)��  ��z�h`xH�Z�� �a��$�>�b��%�6�c��&�.�d��-�&�e��(��f��)��g��*��h��+��i��,��6��� �d��� ��� �� ����� ����� �� ��-� ��� Ȳ�-� ��� �Ζ ��� � z�hX`H�Z��1 �� �ԩ�' �"�J �c� ���"��/� 6��"��.��J� ���1��"��  ����� �"�� ����1�
���2��3 ���2��  ����� �2�� �< ��B��  ����� �B�� �7�;����  ���  ���A�;����
�������m7���� � �� ���i���؍ ��R��  ����� �R�� �;���4�
���5��6 ���b��  ����� �b�� �8���7�
���8��3 �� Ӗ��� ���� �H ����� ���� ���� ��� ���  U� ���  � 9��  ���� �̘) ��J �r�� ԞL���)�'��\�\��]��^�;i�_�8�`�`�N�)���\�0�]�2�^��_��`�. ��)��J i�t��"�J �)��J 8��"��r�J L���J �"� W�L���2� ��L���B� m�L���R� U�L���b� ��L��L�� � �� �� ��z�h`��� ���� � �� ��� �	��  U�`��� �a�� � �����`H�Z����� �ԭ, �� �� �� � �Ȁ��, �����z�h`H�Z��2 �Ϡ � 9� 9� � 9����
 J��
 ���
 �ީ���� �ԭ, �&� �� ��, �����z�h`H�Z���L���\����"��  �� ���\��/��� �"�� �2 ����� ����  .����  ���  �� ��Lݗ�а��� �"�� �3 ����� ����  .����  ���  �� ���  ���� �̘) �W�)��\��	��\L���\Ld��)��\Ld� ��)��J i�t��"�J L���)Ь�J 8��"��r�J L���\��"����8��� V� Ԟ����UL���������8��� V� Ԟ����Uz�h`H�Z�<ə�Li��2��  �� ���]��/��� �2�� � ����� ����  .����  ���  �� ��LC��]� �/��� �2�� �  ����� ����  .����  ���  �� ��LC���� �2�� �0 ����� ����  .����  ���  �� ���  ���� �̘) �u�)��]�0���]L����]i�]�L���)��]���0�]L����]8��]�L�� ��)��J i�t��"�J Li��)Ў�J 8��"��r�J Li��]��3�<ə�)���"�8��� V� Ԟ�<ɐ��i�L�����<Li�� �1�<ə������8��� V� Ԟ�<ɀ��i ؀���<���0�/�<ə�����8��� V� Ԟ�<�p��i0؀���<z�h`H�Z�7�;�LQ��B��  �� ���^��,��� �B�� ���  ����� ����  .��P ���  ��L���/��� �B�� � ����� ����  .����  ���  �� ��L���� �B�� �2 ����� ����  .����  ���  �� ���  ���� �̘) �|�)��^�2���^L{���^m^�^�L{��)�#�^���2�^L{�����^L{���^L{� ��)��J i�t��"�J LQ��)Ї�J 8��"��r�J LQ��^��A�7�;�6��P���*��8�P��� �� V� Ԟ�7i�;��;�7LQ���0�7�;������8��� V� Ԟ�7i�;��;�7���2�.�7�;�����8��� V� Ԟ�7i�;��;�7z�h`H�Z�;��L���_�;���R��  �� ���_��/��� �R�� �5 ����� ����  .����  ���  �� ��Lל��� �R�� �6 ����� ����  .����  ���  �� ���  ���� �̘) �c�)��_��	�;�_L���_i�_Lb��)��_8��_Lb� ��)��J i�t��"�J L���)Р�J 8��"��r�J L���_������8��� V� Ԟ��;L���������8��� V� Ԟ��;z�h`H�Z�8��L���`�8���b��  �� ���`��/��� �b�� �8 ����� ����  .����  ���  �� ��L���� �b�� �3 ����� ����  .����  ���  �� ���  ���� �̘) �W�)��`��	�8�`L���`L���)��`L�� ��)��J i�t��"�J L���)Ь�J 8��"��r�J L���`������8��� V� Ԟ��8L���������8��� V� Ԟ��8z�h`H�
������ 轼���  g��h`HZ �� � �� � �̈��zh`Hڭ�� �' �� �J ��  ���h`H�a�� �' �� �J ��  ��h`H��� �f��  ��h`H�b��  ��h`�Z�P��������z�`HڽJ m �J �h`HڽJ 8� �J �h`H�Z� ���$�0�a�#�b��c��d��e��f��g��h��i�8�7��  ��Ȁ�z�h`� �� �� �� ��  � #� � � � � � � � �� �� ��I�ߍ& `H�	��� �
��� ��� �
�� ��� ����  7�h`��? �����       0� ������       ��<� �?� �0�  <�  ��� � �  <�  ��� � ��<�  ��� �0��<�  ��� ��<�  �� 0� ��<��  0� �? �� < � ?� � `% Z	�V*�Z� P �
P�@�ZH�Z� ������������������� ����  ҡ���r� W���8����ܩh��������8����� ���� � �������� ҡ��8����� ���� ��������� ҡ���D� W�L� W� W����� ������� � ����� G���i����  ҡ���� ������ G���8�����  ҡ���\� W�L}�z�h`xH�Z��
������ 轚��� ���� ���� �� ����� ����� �� JJ���-� ���� i�� �� i �� Η �� � �Ȁ�Ζ �� � �
���� �L��z�hX`H� ��  ҡ���� h`H�Z�/���� ���� ��z�h`����? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                          m���            �                         �                        �?                       ���                       �[�                       �[�                       �k�                       �k�                       �f�                 ���  �f� ���             ��� �f� ���            �UU �f� |U�            o P= �e� _@>           �[ @� �e��[ @�           ����e���
�          �AU��!��dU�          o PP�ZP�od@>         � @@�_T�K d  �         � @F
 Q�U hd  �        � @e@Q�UQ@D  �        o  e ]�U@$  T>       �[  d \�U@  P�       �V �d ]�U@� P�      �U  hD ]�U@P
 @�      oU  Z` ]�E@P) @U>     �[ �V  ]�E @�  U�     �V �  ]�E  � T�    �U h   ]�E  T
 T�    oU ZX  ]�E @	P) PU>   �[U�V V  Q�E @%@� PU�   �VU��  U�U  � �PU�  �UU xp T�T TT@U�  oUU@^\ T�T  4PPm@UU> �[UT�W W� P�T  �E5@�aEU� �V����t  �� @� Ն�U��U%%yp}  �� @PTV�lUII^]w  �� @7PTmXXUkUR�WW�q  �� @�@5P�aaU:���佪�p  �� @C�����Ū:���~��U�UU��sU�U��K���:���PU  ��������  @U���?           ��                      ��                      ��                      ��                      ��                      ���                      �?�                      �?�                 �             �            �?           ���           �[�           �[�           �k�           �k�           �f�       �  �f�  ?    � �f� ��   �� �f� ��  �> �e� ��  �1� �e��_L>  o���e��3�  �P�%�|E�� ���A�jT�_@0��1�T� 4L�� TU�TU s��   �T   @C�  0�U  @p�  0�  t�  p�U  D� p�U  @� t�U 4@�A t�U 4A�  4�Q 4 @�A t�U 4A� t�Q 44@�A< T�T <4A�, T�T 84@�A T�T �4@�A� @�T  �7A�q�  �  @?M�q� �� @?M�q� �� @3M�q� �� @3M�q� �� @�M��� �� @�_���WU��sU�_�5 ������� \�=   ��   |�=   ��   |�?   ��   ��   ���   ��   ���   ��    ���    0    �?�         �?�                 �?                        ���?                     � ��                     �� �                     ���                     � �                      � �                  ��  �� ���             ��� �� ���            �VU �� |U�            �  = ��   >            /  � ���  �           �  ����  �          �  @lT|   �          �|   =lT   @>          o�  �_T�    �         �[�  PUU    �        �V|           �        �|             P>        o|    ��     P�       �[|    ��w     @�      �V|   |����   @�      �U |   �����    U>      oU �  ����    U�     �[ � �����    T�    �V |  ����� w  P�    �U | ���������� PU>    oU | �����������@U�   �[U | ���w�����@U�  �VU | ��������@U�  �UU | ���������! UU>  oUU@| ��������UU� �[UT�| ��������цU��V�������������AVV��U%%y����}�����mXXU>lUII^ |  ����� ���aaU9kUR�W    ��  �  @Ն�U����ZU�|UU���UU=_U�~�꫺�~���?�����������/�������       ��       ����           ��                      ��                      ��                      ��                      ��                      ��                      ��                <          <          <          <          <         ��        ��        ��?      ������?    ������?  ���������������������    ��        ��         �         <        <        <        <        �       ��      ��     �����   ������? ���������   ��       �       <      <      <      <      �     ��    ��   ����? �������   �     <    <    <    <    �   ��? �����  <        �� ��?� � �?�       �   �  �   �?  �������   ������  ���������������  �����+            �   0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���ة��  ��� � � � � �ߍ& �� ��"  `�� t ����� ��� �� � ������ ��� ��XL �H�Z� �Z��Z�%��%�,����*�*��=�*  � <ۭ@��@�I��I� ���I�G��� ��(z�h@H�Z�' )�2�,���% �� ��� � �� �ڜ �.�/� ��.��# �$ �% z�hX@                                                                                                                                                                                                                                                                                �ߍ& ����  �� �� �� ͠ �� �� �� �̩ߍ&  ����E�� �ũ�H *� Ǐ @��p�� �̈�!�  ���� ��������� �E �� [� �� �� ӏ �ũ<� �ũ�H *� �έE� 1����  �Ω�  �ϭ� ɠ� 7�L�� F� }� �� �� ��X��#  v���a���& �� ɠ� ϭa��a� �Ω�%�%���S��S @� %� ӭ� ɠ� Z� �� �� �� 
� 5� >π
��%�%������" �� %� ӭ� ɠ� �� �� �� 
� 5�L�ĭ���LA� �ϭ5��5�4��4�E�'�F�F)��-��  ��
�>�0�L� ��x ��L"  �  ���	������LaĊ��L"��8 w�x���& � � �*  �� �̭  ��� ��X���& � ��  wΩ��� L�­� ɠ���� �̩����ɿ� �� �̊)� �Ɗ)� 'Ǌ)� �Ǌ)� �ǭ4��)� �ȩ
�4�5��) � 9ȩ8�
���5 �٭�2�� ɠ�
�a���a +� �� �حS���SL�©ߍ& � �,x o� �� �ŭY��L"©�� �<�� �F ����� �X�� �G ����' �<�J �c��  힬  ���� �� ��)��,�)��J �<��X��<�J �)�ϭJ �<��X��<�J �� �� Ԟ �έJ �<�	�Y ��LoY ��L"©ߍ& � �,x �� ��Y V����	 O��Lu�� �� ��L"����  ��� ���`H�� �ߍ& �
�� ��� ��  �� t�h`H���G � #�h`H� �Gh`H�Z�� ɠ����� �%�� � �� 7� �� �� %� ���#�� � �� �H�m )�� ���' �0� �d�J �0���' �(� �d�J ɰ�
��' �� ɐ������� ����#Ю�W�m�� � �%  Fʢ� �>�m )�� ���' �F�J �,� �0���' �Z�J �#� ɰ���' �<�J �� ��#иz�h`H�Z�2�%��%8�2}J �J ��28�%�� 8�J � �J z�h`H�Z�� ɠ��a�I�"�' �@�' �H �8 ������S�� � ���2� �	�2��4�  ���#��' ����' z�h`H�Z�� ɠ0�a�I�"�' ��@�' �H �8 ������S�� � ���� �	����  ���#��' �0���' z�h`H�Z�� ɠ��a�H�"�J ɇ�?i�J �k i�k �.�S�� � ������5�J  ���#��J �Ai�J z�h`H�Z�� ɠ��a�H�"�J �2�?8��J �k 8��k �.�S�� � ���9���U�J  ���#��J �!08��J z�h`Hڭ��; �����4�  d����� ɠ��@� �ɀ��� ɠ��( �π ����h`H���'�<�"� d�� ɠ� ɀ [����<8��<�h`H� �������� �� �� �� �� �h`H� ����$��� �ʽ����� �� �� �� ��' �h`H�Z C��#�� �2� ���!� ���!� ���!����� ���8 ��z�h`H�� �	�m )��0���#��h`Hڢ"�' ��� �(���#���� ����� �����  ʜ� ����h`�� � �m )�ɀ0�' ��m8�0�0	��#�֩ ���`H�/��� �h`H���� �h`H�'�� � �h`H�&��� �h`H�Z ������� �Ϡ"�' m�' �J �J z�h`��! �ϩ�" ��`��! �ϩ�" �ϩ ��`Hک��� �7�� ����  �ʭ7i�� ��� �?�� � �� ���h`�k i�� ���  U�`H�Z���� �8�;��� �m;��  ��z�h`H�#�� �l i�� �< <�h`H�
�� �l i�� � <�h`H��� �l i&�� � <�h`H��� �l i&�� �= <̩"�� �l i&�� �> <�h`Hڭ� ɠ�I�� �=�i�9�J �n�2 �˽' ��%��!�J ɉ�Ɍ��A�	8�

�A� ��A ����!й�h`�' ��)��%�J Ʉ�ɒ��Z��[�
��[�8�Z ���[`H�Z�' 8�����D�� �7��� �J �� �B��� ��� ����� ����� �� �� �� ��
.Η �������ȭ���� �� ���C��D�� � ��z�h`Hڪ��� �)�JJJJ W̊) W��h`xH�Z��6��� �d��� �� �� �� ����� ����� �� ����� Ȳ���� �Ι ��� � z�hX`H�Z����� ���  �� ���� ��z�h`H�  )@��h`H�  ���� ��h`H�  ����h`H�� �  ����� �0�h`H�Z������� ���� ��z�h`xH�Z �ͽ/��� ����� �ɀ� �̀ �� β�-� �� !���� Η ��z�hX`xH�Z�� �ͽ��͖ �� 8� �� �/�͗ �� ��� ���� ?�L�ͭɀ� �̀ �� β���� !����� m� �� �� i �� � Η ��z�hX`�)�����	�)���`�' �� �J �� � �ʊ`8�
������ 轿� �͍� `
������ 轿� �͍� `�� �� �� ����� ����� �� `�� i�� �� i �� �Θ `H�Z β�-� �� !���� Η ��z�h`H�Z έ� -� ���Θ 0
��� Η ��z�h`H�Z����� ��� �͍� �
�� �
�� ��� �4��  7�z�h`Hک � � ��#���h`Hک � �� �����h`H�Z�� �@�� � � � ������ ���z�h`H�Z������ ����� � � ����(����m��z�h`H� ��  � U�h`H�Z� ����� ����� � � ����(����P��z�h`HڭV���	� X������ �V�h`H�Z������ ����� � ��	�����(����m��z�h`Hڽ' �� �J �� � �ʽ���� �(8� ͖ �� �/��� �K8� ͗ ��� �h`H�Z� ������ ��z�h`H�Z� ��z�h`�_�� ����' ���J ���m `H�Z� �� ɠ�q�E��F)��-�� ��  �)� �ЭS� vЊ)� �ЭS� �Њ)� �ЭS�� ���J�J �)� ѭS�� ���J�J �S��%�z�h`HZ� �4��5��2�
�2��3��� zh`HZ� ������
������ zh`�� ����#��`� ���#��' �0���' � �`� ���#��' ����' � �` ���#��J �608��J � ` ���#��J �2�i�J � `Hڢ � �� �р ;��h`H�Z��U�� � �� �(�� ����� ��� ���m�� ��  U�����)�� ����� ���'�ˢ:��z�h`H� �����
���������� ����������������  +ҀD�2�������3��������4������
�������  n�h`H�Z�J ����m�,�� � �� ��
�� Ẅ��� W���m� ���z�h`HڽJ ��(���m�0�� �8���� � W̭� �(�� Ẁ�m� ����h`H������h`Hڢ � ��J�� �� �h`���������� `Z ����)�� � ���� �Ѐ vЩ��� z`H�x�� �C�!0���� � Z� �ʀ,�� ɠ��J �n��m )�ɐ��������n�K �ԩ��K��#гX�h`Hڽ � Ͻm )� ��� ���h`H�Z��� ���������_��ʽ����� ����	���� �<�(8�' �01��08�J��' 8��' ��8�J}' �(��'�' ���� ��m z�h`H�Z�� ժ�� �� ���K8�J �� � �ʽ/�͗ ��� z�h`Hڽ �ʽ��8� ��ɀ�8�
����m�� 轿�i  �͍� �
����m�� 轿�i  �͍� �h`H ���� Ԁ � I�h`H�Z���' �. ����'�m ɀ� )����
�� �Ԁ� �ʽ����� ��z�h`Hڽ � ����� � �� ��������� ��� �h`ڽ � �� �	���������`H�Z�m )�� �_�� ���C���m �m � �(� ���!� �Հ'�m ��' � ���!��m ��' 8�J ��J � ��z�h`�� ���' ����!��`�� ���' ����!��`�D ��8�' ��
0 fր�'  5�`�% �8�' ��
0 fր�'  5�`8� ��U���
����m )m� �й' `8� 

����m )m��' `�J �� ���i��J 8���� t�8�J ��J ` t��' m�' `ڭ�� �*��������`�, ��i�8�' ���
0 �ր�'  5�`�= ֍8�' ���
0 �ր�'  5�` t�8�' ��' `�Z��J �J ���ʽ/�����}J ��L��ʽ/�yJ ��J �7�' �' ���ʽ���}' ����ʽ��y' ��' ����� z�`H�Z� ��� ���m )�ɀ� ������ �� �׀��!��z�h` wٹ' m�'  AڹJ m�J `ڹ ��� ɠ��?��J �F��?��7�� �ʽ��m � d� ���`� � �m )�ɠ����
���ɐ�$�-���i����i ��؀���i��؀���i��عm )���� )����� 



����i�ح�����`H�Z� ��� �*��m )�ɠ�ɰ������� ������ �� �׀��!��z�h`Hڢ�� ɠ�T� �H�m )�� �(�0�; b׽ �3�m )�
� � ��"�m �J �J � kؽ ��m )�� � ���!Ю�/� �%�m )�� ��0� b׽ � #Հ kؽ � ?���!���h`H�Z�m )�� �_�� ����U	 �m � �2� �Հ ���m z�h`H�Z��������ݟ�08���J�z�h`Hڢ� ��� � ��!���h`ڢ � ���!������`H�Z�� ɠ�W�� �K�m )�ɀ�B (����; �����9��� �Ϲ � w��' m�(��'  A��J m�J �� � ��!Ыz�h`�' �0�%�J �0�i���`H�Z����/����/�08�/�J�z�h`Hڜ�� �%�m )�ɀ0��)����



�����!���h`H�Z� ��� cڭ��W �����P��!��"�(��� JJJ���"�#����� JJJi�#�h �ϭ"�J �#�' �!�!����!� ��z�h`H��.�����������	�� �ۀ �ۀ ���h`H��-�-�+�;�)�� �����0���)�)�����+� �-�� )i�L�� )?i�N�h`H�G�"���# ��h`H�S�"���# ��h`H�0���M�"�Ѝ# �ۀJ� �ۀ ��h`H�Z�+�-��O�)�J�#� cڭ��: �����3��" �ϭ2�1i)�J �� JJJ���"�' )����m�/� �.z�h`H�Z�P�T�3���'�(�� �L�� �Խm )��`� ��L��ɀ0| �ɰ��T Y�<��� ��3ɠ� � 9ހ'��� � $���3���R����ɐ���� 4ݽ ��+�� �&�m )� �ӽ �� ������ �� � � �m ��!�LAܭ� ���� �� �3��	�2�1�3z�h`H�P�P

mL�'��&�Qh`H�Z ������' �� �� z�h`H�Z �ݭ)�� � � �>�RJ� �ݭ� ɠ�+�2�1�#�8�1}J �J ��18�2��J 8��J �J z�h`�� J��  �)��' ��)��' `Hڽm )��m � J�� �
� �� � �h`H�Z�� ɠ��J �m��0��J ɝ�	�0 ��� � z�h`H�Z�J �� ��� � z�h`�' �'�� � ������� ��	� �� � ���`H�Z �ݽ ��y�y�Ɂ�ɉ� �ހh�z�ɂ�Ɋ� �ހT�{� �߀KɃ� ��Bɋ� ��9�|� �߀0Ʉ� 7��'Ɍ� ���}� �߀Ʌ� ^��ɍ� �� b� ��z�h`HڽJ ���J ��J �h`H��J �h`H�Z�� )i��� )i���m )�d�� �L�߬  �)��)��' ���' �%��' �
�' ���' �)��J ɖ��)��J ɀ��J ���J ɛ�@�J �;�J �6�J��
�J��m �%�J�' ��� ��%�' �`�J � ����m  ��z�h`H ��h`H ��h`Hڭ  )��J �J ��J�� ���h`H�Z�  �)� 	��J �� J��Q�' ��' ��' ��' � �� ��z�h`�S�	� 8�� `�S�	� i� `H�� ɠ� 	�2�& ����2�& ��h`H�� ɠ� 	�N�& ��� �����A�& ��h`Hڭ� ɠ� 	�P�& ��� �����P�& ���h`H�Z�J �&��J ��  )�� Ƀ�Ʉ����J z�h`H�Z�J�B�"�J �J ��J �J ��J ��)�' �' �!��' � �Ȁ�' ��' � �� �Ȁ�' �J �&��J z�h`H�Z�  �)�
�(�" �߀�)�
�'�% 	�� �J�-�' �Q�%0�' � �� �Ȁ�' ��' � �Ȁ�'��' z�h`Hڭ� ɠ� ��J �N��  )��J ��J ��J �h`H�Z�  �)��)��' �Q��' � �� �Ȁ�' ��' � �Ȁ�' z�h`H ��h`H ��h`Hڭ  )��J �J ��J�� ���h`H�Z�  �)� ���J �� J��Q�' ��' ��' ��' � ��z�h`H�Z �ݽ �L��f�� �(��n�	�v�� �' ����'�(L��e�� �(��m�	�u�� �' ����'�(L��d� ��w�l� ��n�t� ��e�c� ��\�k� ��S�s� ��J�b� ��A�j� b�8�r� �/�a�� �(��i�	�q�� �'�� ɠ��i�  ���(�' ��z�h`H�Z�� ɠ�G�J �n� �ހC�' � �Խ' ��� � �Ȁ�' ��!��' � 	�J �N��J ��J ��Z�& 7�z�h`H�Z�� ɠ� 	�K�&  � �����K�& 7�z�h`H�Z�� ɠ� 	�N�&  � �����<�& 7�z�h`H�Z�� ɠ� 	�-�&  ��-�& 7�z�h`H�Z�� ɠ� 	��&  ���& 7�z�h`H�Z�� ɠ� 	��&  ���& 7�z�h`H�Z�J �&��J ��J z�h`H�Z�J�B�"�J �J ��J �J ��J ��)�' �' �!��' � �Ȁ�' ��' � �� �Ȁ�' �J �&��J z�h`H�-�&�� ɠ� P� 7�h`H�<�&�� ɠ� P� 7�h`H�N�&�� ɠ� P� 7�h`H�-�&�� ɠ� �� 7�h`H�N�&�� ɠ� �� 7�h`H�K�&�� ɠ� �� 7�h`�Z� ��& ��" ��� ��?� �I �' �l �J � d���z�`H�Z�  �)��'� 	��J �� J��Q�' ��' ��' ��' � �� ��z�h`H�Z�  �)��(� ���J �� J��Q�' ��' ��' ��' � ��z�h`H�Z�6�LR�


��� )m������>)m�6��� cڭ��M �����F�� �w��� ɠ�:���� �' i�(��'�' �J i�J � ʭ� ɠ���i����m �6z�h`H�Z�T

mL�$��!�M�T


mN�i��P�O �ݽ �LY���J�m )�	�H�' m�
�'�' 8����J m���J 8��d� ��LY�m )�� ]�LY�� ɠ�I� �� �ݬ  �)��)��J��' �M��' ��' � ��
�)��)�4�J �O�,�J �1�m )�%� ��& ��" ��� � ���J �J �J �� � z�h`Hڽ' ���' ��' �J �<��J ��J �h`H�Z �ݽ ��+�m )��& ��" ��� � ���J �J �J �� � z�h`Hک �  ���h`H� ����?��_� �I �' �l �J �a�m �h`Hڭ� ɠ����V� d�78�8�7� �7�?����h`H��>��=�8��=�`�>8��>�h`H�@��?JJ�?��7��7���?��@h`Hڪ�� ���� ����� �� ���� �h`H�Z�� ���C�� 
����� 轇�� �� 

����$�* ȱ�



�� �� ȱӍ) ȱ�� �( �� � ��z�h`�� �* `�� ���Q�� ���.�� � 쭥 �� � �  뭹 � #쭲 �� � �  k�� �� ͧ � j�� �� ʹ � Iꭡ ���.�� � � #쭿 �� � � � �  ���� �� �� � ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��K �K Ȍ� �� �� �� � �LHꮮ �H�� ���� �� ��� ��� � ��� ��莮 �� ���� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��K�� �K�� Ȍ� �� �� �� � �#� ��  � #쭥 �� � � �� �� � � `�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��K �K Ȍ� �� �� �� � н�� �H�� ���� �� �� ��� � ��� ��莻 �� ���[ �[ `�5 �5 `�q �q `�c �c `�= �= `�} �} `H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����έ �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����κ �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� �Ī�� )@��J��� �� Ȍ� ������� �� �� �� � �� � �� z�h`� �� `� �� `H�Z�H�� ���� h� �윢 �� ��� ��  j� I� � k���� z�h`�5 �= �6 �> `�[ �c �\ �d `�q �} �r �~ `H�Z�C �D �� ���  �� ����� z�h`H�Z�E �F �� ���  �� ����� z�h`H�Z�G �H �� ���  �� ����� z�h`.� �� �� �� ���.��@���� �� �� �� ���� �� ��� ��   @�.� �� �� �� ���.� �� �� ��   � ��� �� �� ��� ��@�.� �   \���\���\���\�������\��������\���   \������\���\��������\���\�\�    �    �� �� �� �� �    �� /2�   �
	�
�
�
	�	�

		�%����   �X�  �����  ����������������)�  �����"�f���  ��-�b����  $����O�  ����  

  �� �� �� �� �$� �� �� �� �� �H� ��    �� �� � $� �� � �� � qH� d� q� �    q� q$� �� � q� �� �H� �� �� � q0� d� q� � �� �� �� �� �H�   ��������h�h�����   ����������.�.���.�.���������T�T�T�T�T�����   ��T�T�T�������T���T���T�T�   ������ ��T�T���h�����h���������h�T�T���   h���h�����������T0�    ?� ?� ?
� ?
� ?
� G
� O� G
� T
� O
�    ?
� (� G� G� G
� G
� G
� O
� T� O
�    T
� _
� �
� (� 
� _
� T
� O
�    ?
� G
� ;
� ?
� /
� /� /� /
� 5
� ;
� ?
� � G
� ;
� ?
� /
� ;
� /� 5� ?
�    
� G
� ;
� ?
� O
� ?
� T
� ?
� _P�    
� �
� 
� �
� 
�
� 
�@
� 
�
� �
�@
� 
� �
� 
� �
� 
�
� 
�
� 
�@
� 
�T
�    
� �
�}
�T
� 
� �
� 
� �
�}
� 
� �
� 
�}
�    
� �
� 
�}
� 
�@
� 
�@
� 
�@
� 
�T
� 
� �
� 
�
� 
�}
� 
�T
� 
�    �
� 
� �
� 
� �
� 
�T
� �
� �
� �
� �
� �� ��   +.148<AGMSZahpx�����+036:>DJPW^elt|����-037;?EKQX_fnv~����/259=BHNU\cjrz�����    ���������������������������������������������������������������������������������������������������������������������������������������-�C�[�s�������� �8�O�g�����
 �� 
 ���  ��� 
 ��� 

 ��� 
	 ���� 	

 ��� 	
 �� 	
 �� 
2->:64(<20(6<&.40*3:"6.,(&0,*$.,!($/"'"$ ($"
	
           	
   !"#$% '()*+,   012345 789:;<= ?@ABCD   HIJKL NOPQR TUVW YZ[\  _`abcdef  ijklmn  qrstuv  yz{|}~  ������  ������      
          "!          





  





  





  





  





  





  ����  cB� g
 mIIUF2
2P �<diZF2 ddl_K7- dcqvvU cciZF2 cci_K7- 2<FPZ 2<FPZ 2<FP 2<FP    ��nZF2  ��nZF2  ��nZF2  2FZn�  2FZn�  2FZn�    ������� �RR���� �B/44444 ??!!!!!! /���� ee44444 ee!!!!!! ����� ����� ���� ����  dd������  ������  ������  ������  ������  ������    	 (($$   	    
    	
  
	  
  
  	
  
  113/  
 		3GGG	 	  
G 	  	 	
 	   !  
      
    ������F��������A����c��������A�B9S�U�������C�C�B�B�B@C���A�C�A�AB=BYBdB���A�AmB�B�B�B�B�B���A������������9MN�AB=BYBdB��SL�LmB�B�B�B�B�B���N�N�NO>O���O�O�O�O<P���P�P�P)Q��������������hQRR�CEK�K�I�C�C�����C~D�D0E�C�C�����C�I�JK�C�C�����CXE
H�G�FmE�����CXE�FxFFmE�����CXErII_HmE���� �] 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p�����Ѐ���������������������������������������������Kd}bhn                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          O� ���