xآ���ɍ& ���  ��� ����� � � � �H�H�H� H� �� ������������� ��h� h�h�h� E� w�����!���� �" ��{� ���� � � ����� i� �i ���� ��� )��;�<���[ �)��=��=�;)�S�<��L����:���9��� s��<���:� �9���i s��<L�@@@@@@8  0@P`8@@@@@@p�����Т �{�	�}8��}�����p��{�	�}i�}���������#�;i�;�;ɀ�L��d�ɴ�
�	���	��L��

�����{���Á���ā���:�z�~i�����9�}��i����� �|������`	
+,)*78'(56%&34#$12!"/0 -.���!��"��4�7�+��'�$���,�-������q�� Ǘ Tũ�� W��-�	��)� �ϭ	���� ��L热-�,��+�1�-�>�@����$�'����0 �� E� �� �i��j���� C��� )��� )�L�Thin Chen Enterprise
      presents



   @1989 & @1992

      PYRAMID



Design by:
     L.C. Tchacvosky
Artist by:
     Shyh-Dwo Maa
Music by:
     L.C. Tchacvosky  E����	� �� �ϭ���� ��	���� ��-I�-L`�`8`�x�j�
�i�-
�������LC���˃  PYRAMID  
  T-BLOCK     RYRAMID  
  T-BLOCK   ����� � � �� ��� ����� ������
��&���'��l 6�6�9�I�w�S�9���L���3���� �3L���3�����3��1�4�r��� �4�� �L��

�3���4:�r�:Le��5�0��1 �L��� �� ��3����J�K�]��j�i�
H��q��r� K���i�b���  �Lʄz�g���h�� �������`l �4
�����LK����  EASY  NORMAL    HARD  �5	0 썩 L썭6	0 썩 L썭7
��G��H�LK�M�R�W�off    1    2  `@HPX`$$ (��,�9�\�{��������� difficult  start level  start line  music  play � ��$�%�& E� )��+�7�6�2���� )��)�� ������ ������� )���ҩ�������� Ǘ�a������  �� �� �� � �� �� a��� �� ����� a������� �� � �������@�Z�+� ��� ��������8���


�� 4�z�����Μ�L/������	����� �� � � 㻭���) ���$� ������ ��
������ޭ�п���L6����
��2�	
��$���%�� �L�l 

D���Ň	���'�b��c�x���b�b�b�b��� ҿ�5��)���Hi��� ҿh�����Hi��� �h��`���
�`����  ҿ���)���Hi���  ҿh���ѭ�H8����  �h���`��)�� ҿ�2��Hi��� ҿh�����Hm.m.)��� 4�h��`���`�+�
���2��1�	 ƽ�1L��`�����H�)����)������H}������)�� ҿ�%��Hi��� ҿh��� 4��h�� Ќ�`�h�����`                        ��������������H�)���ʊ)������H}������)�� ҿ�%��Hi��� ҿh��� 4��h�� Ќ�`�h�����`  �R�������� �	���	���	��� � ������� �L"� @ H P X`�2������h��i��`�2��㭕�0��8���`�2��� ;���`�+�`�)��A�?�A�@07�	�@ ��L쉮>�	����$���	�@�>L�JJJJ�?�	�)�@�> ��8`hh�<L)��?
��$���%��l�@�P ����Q� �Q�Q��A�Q�Q �0���� E������ک��� ���  � � ы�� ��L4� �ĩO�� W��j�(�i�1�� C���j�(�i�8�� C��@��(�� ǘ�i(��i ��O ǘ�i��i ��i0��i ����������i0��i ��8�0��� �� )���	� ?�L���)����$�!�-�� ��ߢ� W��)��)��A��A)� �L� ��L�L�GAME OVER ��H�H�O8� ǘ�i��i ��i0��i ��Oe ǘ�i��i ��i0��i �������� ������%��i0���i ���8�0���� �L��h�h��`ZڠP� �������z`�0����.����/`   � � �@�� �� � �������`� ��z�[���`e���`�  �  ���  �����  ���  ����`@Hm��Hm��Hm�m � ���
��
���  I���
>���	��+����xL� �� ��h�h�h@�B�� �C� �����CmG�C�H��B`
�
e�� �ꌙC������B`�,
��� 8� � 
�@@ 
��<� �<�@S0����+�LE��7
��*��+�LW��\�Z�TRADE MARK "SACHEN"�J��K���i�N�j�O� ���
���*�	�-��, � ɍL[�`�N�i�jiɪ�骍jLt�� �i��Lt� ɍ�H)�KhJJJJ�JLt�HJJJJ ��h)	0�:�iL����`�ڍS�T�U َ��V	0 ���`�L�MH


iǅ��i �hJJJJJe��j ǘ�mi��i ���P� ��JH�K��JJj.Q.R
.Q.Rh���Q�ȭR� 䛥i0��i ��Pн ���L�M`�h� �U,�-�^��SI��S���Si�S� mT�T� mU�U� َ���V�����V	0�^��h��� �^��h��� �^`�SH�TH�UH�� �V�����S8�G��S�T��G��T�U��G���U�V��L򎈈�SyG��SȭTyG��T���о�S�Vh�Uh�Th�S`���@B��' � d  
  � �U�T�]�S��UH�TH�SHS.T.US.T.UhmS�ShmT�ThmU�US.T.U�VmS�S� mT�T� mU�U��`                                                                                                                                 08<80                                                                                                                                  <<  cc"     66666 ?T>~ac3c 6;nf; 00`     000   66   ~    0    ~           0` >cgksc> ? >c0c >cc> 6f `~c> 0`~cc> c >cc>cc> >cc?<       0 0`0   ~  ~  00 >cc  |�����| 6ccc ~33>33~ 3```3 |63336| 14<41 14<40x 3`oc3 cccccc << f< s36<63s x00001 cwkccc cs{ogc 6ccc6 ~33>00x >ccko> ~33>63s >c`c> ~Z< cccccc> ����f< �����ff �f<<f� �f<< C1 <00000< `p8 << 6c                  <>f; p0<633n   >c`c> 6ff;   >c`> 20|00x   ;ff><p06;33s    f<p036<6s    v{kkk   n3333   >ccc>   n33>0x  ;ff>  n300x   0> ~   ffff;   cc6   ckwc   c66c   33<  ~0~ p   pp ;n       6cc  ?_/W(T �����
(T(W/_?

����� �����     �����(T(T(T(T



88((88� ���     ?��     ���     ��� 4  b  � �� � ?�  � ���������!�����	���������q�pa� � � �  �@@@` ��,.((�h  `�  �        ������������������������  U�U�  ((((��������癙~~�����������$B��$$<<$$�B$(O��O(��                                                        ��ժ������U�U�����W�]����������������������������������ժ����U�U�����]�W�            �   �       �    �   �                                                                                                                                                        �        			`�������
�l`   �ff<8    �����`�` `����  >>6~`&<��~nz�>6   X� ������p	~d|a ؠ�`���?�?                                                                                                                                          ���{����� �������i��i ��i��i ���ة{����j�i� � G�����jɨ��`�Z��iJ�&�jJJ��a�e&�'�b�i �(�H� �'hz��t�u�



e��i ��JJJJe��j ǘ�mi��� ��ȱ��i�� e��i0��i ���� ���u�t`�j�i���0�� iɪ�骍j�i`H)��★hJJJJ�
ei@}�` 0`��� P���@p��      �)��}�`�}�#��d#�[���� �0n�iȱ�j
��a�mi��b�i �ijjj� � G��i��i �L�{�����#;Sk������+C�@ �[����;� �;��� �|){�Z ��z������ ���`�z�vJJJ�j�{�w�|�x�}�yJJJ�iJJJ�k�x)�i�p�JJJ	�s�x)J�i�q�J	�r�j
mjmk��i)��s�l�Z�iH�r�m�;=���%�;���;Z� �i�ȭj��i��i �z�m��i���Ƣ ���h�iz��j����lФ�0�$d%�v�xmp:H���%E$�$h ǘ�yJJe��i ��w�



He!��"i ��xJ�jJJJHe�he �he��i ��y)�t�q���k,xp���k��0�� �ڪ�����k��t�#8.k.l.m.n.o8.k.l.m.n.o��ݬq�k1����q� �k,xp���k��0�� �ڪ�����k��t�!k.l.m.n.ok.l.m.n.o��߬q�kQ����e$��e%��mq��i ��mq��i ��p�L��`���`���`��}�`�}� � �Z�[�z��\�{��]�|��^�}�L�])\��[�v�\�w�]�x�^�yZ ��z�z�[�{�\�|�]�}�^�|){� y�z������Љ`�z�v�{�w�|�x�}�y�x)i�p�x)Ji�q�0�$d%�v�xmp:H���%E$�$h ǘ�w�



e�� i ��xJ�jJJJe��y)�tNyNy�q� �k,xp���k��0�� �ڪ�����k��t�!k.l.m.n.ok.l.m.n.o��߬y� �(��@�	� �kQ����q��e$��e%��mq��i ��p�L��` @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��Hژ��7
�h�+h�*`�F�G� �FH
������������ �����`l���Ϟݞ� �F� �����`� �F� �����`� �F�( ��������F`� �)��� �)��)�� �~��� �~��"�� � � �( ����`d) ��!���~���(���)��` W��)��`�(t)���!�~��L��~�2�3� � �2�*��������7� �4�����:�;�<�)`�)�`�:��L�����;��;�`� �:�<m~�;�7�
�4�	�4�� L�������*�0�+�1�:� �00LB����LE����L^����� �7����� ��0�<m~�; �LΟ��� ��0���08��0�1� �1LΟ���Le�������}�����0���1 �LΟ���- ��0H ��0H�}���0���1����h�1h�0LΟ���' ��:���� �0��������0i�0� e1�1�:LΟ��� ��0Hȱ0�1h�0LΟ���2�����)���:��� ��� ��0�����:�4Lw� � �LΟ����:���)���)����� ��:LΟɀ�(逼��

��Ţ���Ƣ���Ǣ���Ȣ�� ��:LΟ�:��������<�� �p�� ��� ���  �� �0�����:�4 ��:
��0�*�1�+�:����ޚ��`�9��6��6�L��� �.���� �9L����� ��.���.8��.�/� �/L��

� ��.�����6 �����( ����) ���)�* 	�* L��   �0��1`�.��/`H����
��hJH��m���hn�n��뮟��`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P             	        
                                                                                       !"        #$%&                                                        '        ()*+,                
����h� >P����������*� �Uݪ�]�]��A��]�������_u�uO3_3�u������ww�3�3 wU����� �
�_) ����UU������

��

��UU������""""����������>�����������������""""����""""����

��

��

��

������֧v���~�����v�v�֧����TUTU ?��UUUU  �?� �� �?UUUU  ���� ��UU5 8�88888TUTU ���UUUU  C�0�0�0CUUUU  �����3��UU5 8?8�8?8�8?8         8 8 8 8 8 8 8 8      ����            ���� 8 8 8 8 8 8�:�?     ����TU          ����UU 8 8 8 8 8�:�?UTUTU �����UUUU   � � � �?�UUUU  ���<���<��UU5 88 88 88UUTU �UUUU  �3<0��<���UUUU  �?��?��?UU5 88888�8������>����������������Ƿ��T>P X��~���U�U� �?�����wUwU3 3�w������ )O)���/�                 @ � � �@�P�Կ�� 	 ) � ��
�+����P�@� � � � @  �:��� =     ��Y�i����֥��k����~������}�]���UUVU
P
P
P
P�j�����
�
#ȏ���5�����     PTUUUUUUUUTP�
�*���������*�
��?���������?������0?�  ??0��  ?�� �  �����������                         	
            !"#$%&'()*+,     -./0123456789:       ;<=>?@ABCDEF        GHIJKLMNOPQR         STUVWXYZ[\          ]^_`abcdef          ghijklmnop         qrstuvwxssyz        {|}~�������            ����                ����                 ��                                                                                                                                       ������           ��          ���?          �?�?�_          ������          ���               @          	 	 (                �          ?�?���           �?           �?�?��          ������          ��?�������������������_�����_�WU�?���������T�Q��_�W�W�U�UOUOUU��������������������_�_�U UT @PTTUUEQ( � ���
�
�*�� � �   0 0 < � ����������������??� � � ����?�?�?�?�?�?�?�?��������������������������������        �O�O�O�O�OUE@PUUUUTUPU@U U Q�E���� T  @TP@@@@ @U@����������UQTEPPU� ��OUEUQUQQ�T�T�U�U����������������� �������*U�T�T�?�?�?����EUQTE����?�?TUUA�?�?�?�?�?TUU����������PUTUE��������WTUU            @U U T P        E      UU              UUUATEPU@U      UU@U U T P      UTTU�U�@P�T����T6jZ����jK��wF�	�f��*���Qk
���J�J�*�**���F*UQUTUEU     ��UPTEUAU      ��U@QUU      ��UQUTUE      ��U              PP@U U U T        ������U�        ��������   @ @ P�T�**Ņ\!������
{zԿ��$�U�`d�������������o�熹���j_��8 2 � � ��)�%�+�        ��������        ������� � � *�*�
���  T P @ @        U�U�U�U�U�UUTUPU�����������*�J�JJ�R�R�TaT�U�UU�q��zZp
�@Y�kO��BE@A��TT@϶�� td h i@jQj�ժ��������媔����•����P���������������������������������*� * 
 
       PU@U@U U T T P P�R�R�TUUEUQUQU���jEU��``��j@e����U��� ���_UPUUPVTZ�����Q��������ڪ����j����jU ������P��*�/�*P*�*����������������*�
�
�� � * *  @     @ @ P T TTTU�U�U�U�U�����?�?j�������� ��� ���@���@�g�꧵��������Z�Z���������UU @�� P�� ��� ��*�ʿ�*����������ꧪ����������    
 
 * �  U U@UPUPUTUU��������������������������X���X��@���@���@���@꧸W�����[�������������n��k��@��/P*����ʥ�������������������������������� ���
�
�*����   @ @ P T T U@UU�U�U����������������������������h�c������������A���A���E���F�������� �?�?�?��[ ��[@��[@��jP�ƥ����i�o�����������������  
 
 * * � �@UPP�T�����    ��  ��������    ��  ��������    �  �j�j����    V*�J���������PU�?U�*�*����������i���ii�R�����FU�����������*��UU��������    �UU��������    ��
�
j)���Z    PU@U U U T T P @����������U�U�U����������������*�
�
�� � * 
  @              U�U�U�T�PUPU@U@U��������*�*�
�

              U T T P P @    �� � ) ) 	                      P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������2��͍�`����������ΑL��/����)�� ҿ���.Hi��� ҿh�����Hm.�� 4�h�����L���������� ЌΏ���� &��������L�`��)��m�)�����)��m�)�����������ʸ����)��J��JJJJ���
�����H����I�J� �H�����̒��eH�H�Ii �I�Ji�Γ��`�"���(�j��������ʸ����
�����H����I� � �����i� �J� �����H����  �ȦJ�������   ��ji�j������`��������ʸ��� ��
�����H����I� �H0�����{ Z������� ��i����i0����� �|���}i�����z������i��Γ��`         Z�]�`�c�f�k�p�u�z�}���������������������������������ȹϹֹݹ����� �����#�*�1�8�?�F�K�P�U����� � � � ��������� � � � �����  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ������H��I`�+����p��`   Z�-�ĺ�4}ƺ����mmm )m���ɺ� �	͜��L����

z`   0            			

		

	
��� �����`����JJJ}���	�8�`��)���J��JJJ}ʸeJ��὚����ʸ���J


m�)��J��JJJJ���
�����H����I�J� �H���H]�� �5���0�H�,������ ��̒�ԘeH�H�Ii �I�Ji�Γй`8� `����`
�����H����IlH  �L� ����ʸ����)��� �J����������Δ��J��ȥJi�Γ�׌�� �������`�)�͟����� Ќ���Ξ� �� f��̖��`� ��ک�J����� ����J��h8���Ly��̖�٘m � �i � ��Ώ�-������1 �ĭ��-�
 � � �ĭ0�	�#8�5
�������� ���	�0 �� ��` ( < P d x � � � ���
��\�m$�$�]�m%�%� m&�&��$�!������`�$�!�%�"�&�#�`  P � @�ZH)�i ǘh)
i�e��i �� �I�������0���z�`� � �������`�Z�H)�i�jh)
i�i�����  �z�`�2���z��{��|�H�}���� W�`�2
�����H����IlH �� �+�`�)�͠���� ;��2������������`�`�)�͠�ˍ�� Ќ����&�����}ƾ�z����{� �|��}���}�`�� �z��4��� �2��)�J��Jy��0����y��ɐ�
�� ��� ����L��  $(,0

 ���
��8�)�ɀ��J��8�0JJJeJi����`
�� ����)����Hi�� �h��`����JJJ}���	�8�`��������ʸ����)��J��JJJJ���
�����H����I�J� �H��H�H]�� �b���]�H�Y����.��*��I�������o��;�p��6������H���)�#��̒���eH�H�Ii �I�Ji�Γ�LX�`8� `
����JJJ���`��������ʸ����)��J��JJJeJ���
�����H����I�J� �H�������� ]����������H�o��+�p��&����̒�ǘeH�H�Ii �I�Ji�Γ�L�`8� `� ��@���������`�����[������d���ͦ���� �� �������魪����i<���`

�� ���� � �����`� �/ ����Χ`������@�]�<��8� ǘ�i0��i �������������i0���i ���㭩���  P­��a�1�]�-�D ǘ����ȑ�� ��� ��i0��i ���ߩ��� ���_��a�Ș �����a�����`�`���Ψ`���M�]�I��8� ǘ�i��i ��i0��i �������������i0���i ���㭪��� P­��a�1�]�-�D ǘ��ȱ����'��� ��i0��i ���ߩ�����a�����`�`



}����i ��J��� ǘ���e��i ������`�� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �+�� �i�h�j����LC�Demo �#�i�h�j�J��K�0	0L썩�i�h�j�J��K� �S��T َ�L7ũ�i�0�j�J��K�1LЍ��i�j�!�S�"�T�#�U َ�L7Ŝi�j�$�S�%�T�&�UL�ʠ �V�� �� ��0��I0 ���`�x�j�i�c��LC�
      PYRAMID       

    @1989 & @1992
Thin Chen Enterprise �i�(�j����LC������� OPTION ������









�������������������� ��i�@�j��� C���i�P�jL�HI-SCORE ����%��G���  

	�  	�  

	�  	�  
	�  �  
�  �  

�  �  
	#�  $�  


	$�  �  
0���  $            
  
  
  
      
  
  
  

  
  
  

  
  
  
                              
  
  
  

  
  
  
                                    
  
  
  

  
  
  
                        �    ��b���&���  "0((((('�  &(����������������	#   	 	# 	 #	#    #	"	��  2((((('((((('((((('(                                                        ��                     �	`���Q���  $
		
		0	""		0��  #	                        �UΛ�����  /���  3										����7φ���  /	���  4(		���Ϩϲ�� �  &      ��  20 �����  ͬ�I�  �������=���9��2���	�- E� ����i�8�j� ��Ii�z��<��z� C�L�Ϝ�`IIIIIIA*@XPP[cc=! 'I*!,'I,'=,;9; :,ccIIIIII9;,:,'=:i���������  /���  3										����7φ���  /	  O  ���  4(		���Ϩϲ�� �  &      ��  20 �����  ͬ�I�  �������=���9��2���	�- E� ����i�8�j� ��Ii�z��<��z� C�L�B  P  Ϝ�`IIIII                        ������           ��          ���?          �?�?�_          ������          ���               @          	 	 (                �          ?�?���           �?           �?�?��          ������          ��?�������������������_�����_�WU�?���������T�Q��_�W�W�U�UOUOUU��������������������_�_�U UT @PTTUUEQ( � ���
�
�*�� � �   0 0 < � ����������������??� � � ����?�?�?�?�?�?�?�?��������������������������������        �O�O�O�O�OUE@PUUUUTUPU@U U Q�E���� T  @TP@@@@ @U@����������UQTEPPU� ��OUEUQUQQ�T�T�U�U����������������� �������*U�T�T�?�?�?����EUQTE����?�?TUUA�?�?�?�?�?TUU����������PUTUE��������WTUU            @U U T P        E      UU              UUUATEPU@U      UU@U U T P      UTTU�U�@P�T����T6jZ����jK��wF�	�f��*���Qk
���J�J�*�**���F*UQUTUEU     ��UPTEUAU      ��U@QUU      ��UQUTUE      ��U              PP@U U U T        ������U�        ��������   @ @ P�T�**Ņ\!������
{zԿ��$�U�`d�������������o�熹���j_��8 2 � � ��)�%�+�        ��������        ������� � � *�*�
���  T P @ @        U�U�U�U�U�UUTUPU�����������*�J�JJ�R�R�TaT�U�UU�q��zZp
�@Y�kO��BE@A��TT@϶�� td h i@jQj�ժ��������媔����•����P���������������������������������*� * 
 
       PU@U@U U T T P P�R�R�TUUEUQUQU���jEU��``��j@e����U��� ���_UPUUPVTZ�����Q��������ڪ����j����jU ������P��*�/�*P*�*����������������*�
�
�� � * *  @     @ @ P T TTTU�U�U�U�U�����?�?j�������� ��� ���@���@�g�꧵��������Z�Z���������UU @�� P�� ��� ��*�ʿ�*����������ꧪ����������    
 
 * �  U U@UPUPUTUU��������������������������X���X��@���@���@���@꧸W�����[�������������n��k��@��/P*����ʥ�������������������������������� ���
�
�*����   @ @ P T T U@UU�U�U����������������������������h�c������������A���A���E���F�������� �?�?�?��[ ��[@��[@��jP�ƥ����i�o�����������������  
 
 * * � �@UPP�T�����    ��  ��������    ��  ��������    �  �j�j����    V*�J���������PU�?U�*�*����������i���ii�R�����FU�����������*��UU��������    �UU��������    ��
�
j)���Z    PU@U U U T T P @����������U�U�U����������������*�
�
�� � * 
  @              U�U�U�T�PUPU@U@U��������*�*�
�

              U T T P P @    �� � ) ) 	                      P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������2��͍�`����������ΑL��/����)�� Ͽ���.Hi��� Ͽh�����Hm.�� 1�h�����L���������� ͌Ώ���� #��������L�`��)��m�)�����)��m�)�����������Ǹ����)��J��JJJJ���
�����H����I�J� �H�����̒��eH�H�Ii �I�Ji�Γ��`�"���(�j��������Ǹ����
�����H����I� � �����i� �J� �����H���� �ȦJ�������  ��ji�j������`��������Ǹ��� ��
�����H����I� �H0�����{ W������� ��i����i0����� �|���}i�����z������i��Γ��`         W�Z�]�`�c�h�m�r�w�z�}�������������������������������Ź̹ӹڹ����������� �'�.�5�<�C�H�M�R����� � � � ��������� � � � �����  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  ������H��I`�+����m��`   Z�-����4}ú����mmm )m���ƺ� �	͜��L����

z`   0            			

		

	
��� �����`����JJJ}���	�8�`��)���J��JJJ}ǸeJ��ὗ����Ǹ���J


m�)��J��JJJJ���
�����H����I�J� �H���H]�� �5���0�H�,������ ��̒�ԘeH�H�Ii �I�Ji�Γй`8� `����`
�����H����IlH ��I������Ǹ����)��� �J����������Δ��J��ȥJi�Γ�׌�� �������`�)�͟����� ͌���Ξ� �� c��̖��`� ��ک�J����� ����J��h8���Lv��̖�٘m � �i � ��Ώ�-�������1 �ĭ��-�
 � � �ĭ0�	�#8�5
�������� � ��	�0 �� ݋` ( < P d x � � � ���
��Y�m$�$�Z�m%�%� m&�&��$�!������`�$�!�%�"�&�#�`  P � @�ZH)�i Ęh)
i�e��i �� �I�������0���z�`� � �������`�Z�H)�i�jh)
i�i����� �z�`�2���z��{��|�H�}���� T�`�2
�����H����IlH ����(�`�)�͠���� ʾ��2������������`�`�)�͠�ˍ�� ͌����&�����}þ�z����{� �|��}���}�`�� �z��4��� 2��)�J��Jy��0����y��ɐ�
�� ��� ����L��  $(,0

 ���
��8�)�ɀ��J��8�0JJJeJi����`
�� ����)����Hi�� �h��`����JJJ}���	�8�`��������Ǹ����)��J��JJJJ���
�����H����I�J� �H��H�H]�� �b���]�H�Y����.��*��I�������l��;�m��6������H���)�#��̒���eH�H�Ii �I�Ji�Γ�LU�`8� `
����JJJ���`��������Ǹ����)��J��JJJeJ���
�����H����I�J� �H�������� ]����������H�l��+�m��&����̒�ǘeH�H�Ii �I�Ji�Γ�L�`8� `� ��@���������`�����[������d���ͦ���� �� �������魪����i<���`

�� ���� � �����`� �/ ����Χ`������@�]�<��8� Ę�i0��i �������������i0���i ���㭩���  M­��a�1�]�-�D Ę����ȑ�� ��� ��i0��i ���ߩ��� ���_��a�Ș �����a�����`�`���Ψ`���M�]�I��8� Ę�i��i ��i0��i �������������i0���i ���㭪��� M­��a�1�]�-�D Ę��ȱ����'��� ��i0��i ���ߩ�����a�����`�`



}~��i ��J��� Ę���e��i ������`�� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �+�� �i�h�j����L@�Demo �#�i�h�j�J��K�0	0L鍩�i�h�j�J��K� �S��T ֎�L4ũ�i�0�j�J��K�1L͍��i�j�!�S�"�T�#�U ֎�L4Ŝi�j�$�S�%�T�&�UL�ʠ �V�� �� ��0��I0 ���`�x�j�i�`��L@�
      PYRAMID       

    @1989 & @1992
Thin Chen Enterprise �i�(�j����L@������� OPTION ������









�������������������� ��i�@�j�
�� @���i�P�jL��HI-SCORE ����"��D���  

	�  	�  

	�  	�  
	�  �  
�  �  

�  �  
	#�  $�  


	$�  �  
0���  $            
  
  
  
      
  
  
  

  
  
  

  
  
  
                              
  
  
  

  
  
  
                                    
  
  
  

  
  
  
                        �    ��_���#���  "0((((('�  &(����������������	#   	 	# 	 #	#    #	"	��  2((((('((((('((((('(                                                        ��                     �	]���N���  $
		
		0	""		0��  #	                        �RΘ�����  /���  3										����4σ���  /	���  4(		���ϥϯ�� �  &      ��  20 �����  ͬ�I�  �������=���6��2���	�- B� ����i�8�j� ��Ii�z��<��z� @�L�Ϝ�`IIIIIIA*@XPP[cc=! 'I*!,'I,'=,;9; :,ccIIIIII9;,:,'=:i���������  /���  3										����4σ���  /	  O  ���  4(		���ϥϯ�� �  &      ��  20 �����  ͬ�I�  �������=���6��2���	�- B� ����i�8�j� ��Ii�z��<��z� @�L�Ϝ�?  P  `IIIIIIA*01:get_scr_adr
9909/001909/01:draw_sprite_all
99C8/0019C8/01:draw_sprite
9BEB/001BEB/01:inc_sou_adr
9BF2/001BF2/01:inc_sou2_adr
9BF9/001BF9/01:xor_sprite_all
9C80/001C80/01:xor_sprite
9D90/001D90/01:hori_inverse
9E90/001E90/01:minsert_channel
9E9F/001E9F/01:meffect
9EF6/001EF6/01:pausemusic
9F29/001F29/01:replaymusic
9F44/001F44/01:mwaitsong
9F4C/001F4C/01:mdismusic
9F5E/001F5E/01:mplaymusic
9F8F/001F8F/01:music
A308/002308/01:p_game
A498/002498/01:d_game
A768/002768/01:spr_pic
A878/002878/01:p_title
AA08/002A08/01:d_title
B308/003308/01:p_sachen
B698/003698/01:action_block
B72D/00372D/01:set_block
B7AA/0037AA/01:print_next_block
B81A/00381A/01:draw_block
B8A1/0038A1/01:blk_xsize
BA68/003A68/01:get_block_type
BB30/003B30/01:clear_block_buffer
BB3B/003B3B/01:check_drop
BBEA/003BEA/01:check_line_finish
BD1E/003D1E/01:add_bonus
BDA0/003DA0/01:print_block_all
BDAC/003DAC/01:print_single_block
BDCD/003DCD/01:set_bomb
BDEE/003DEE/01:action_bomb
BED4/003ED4/01:check_bomb
BEF7/003        �UΛ�����  /���  3										����7φ���  /	���  4(		���Ϩϲ�� �  &      ��  20 �����  ͬ�I�  �������=���9��2���	�- E� ����i�8�j� ��Ii�xة�& L �N�����