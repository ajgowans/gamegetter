 8� Q����{���| t�d������o��p��u���v w���� �׭  )����  )����ע� �ש2H H�h:��`��i� Z��o�	�p�)
����u���v��H �� ���iz���`�i�:�����`       ��
                                     ( �   �
  �   �
 �� �
�
 �
                        ��             �             ��              `UUU%  V%  V   V%  VV`% V           XUUU� �U�  V  �U�  VV`��U           XU�U� �U�  V  �U�  X�� ����            VUVU�U�  V  �U�  X�� �Ub�            V� XU�U�  V  �U�  `e%  Vj%            V% `U`�U V  `�U `U%  VU%            �* ���*� �  �*� ��
  ��
            �* ���*� �  �*� ��
  ��            �* ���*� �  �*� ��
  ��             �* ���
�
 �  �
�
 ��
  ��             �*    ���
 �  ���
 ��*  ��             �*    ���
 �  ���
 ��*  ��             �*    ���
 �  ���
 ���  ��             �*    ���* �  ���/ ���  ��             �/    ���/ ��� ���/ �� ��             �/    ��/ ��� ��/ �� ��             �/   ��� �����࿀� � ��             �/   �� �� ����� ���� � ��             �/   �� �� ����� ���� �
 ��             �/                                      �/                                      �/          �*                          �/    ����* �� � �������
��            �/    ����/���� ���������            �/�������/���� ���������/            �/�������/�/�� �������
��            �/���� �/��� ���/  ���            �*���� �*�
�
� ���/  � �            �*���� �*�
  � ��
�*  � �            �*���� �*�
  ����
��� ���            �* ����
�*�
  ����
��� ���            �* ����
�*�
  ����
��� ��*            �* ����
�*�
�
����
��� ��
            �� ����
�*�
�
� ��
�%  VZ            VUVUX �%`	X	� X`	�%  �X	            XU�U� X �%`	`	� X`	�%  �`	            XUUU� X �%`	`	� X`	�%  �`%            `UUU% X �%`%X	� X`	���
��%            �     � ���  �  ���                 � �  �  �  � �             ( �  � �* � � ��
���
� �             ��
        �*                                                                                                                       @                                     @  @                                                                                                                @                               @@    @                                  @      @                                 A                               @ @ �   A                               T                                 @D   T A                             @ A  T   @                             @ T                                   X                                   U	                                @)                                    P��   @ @                             P�                                    P�                              D  ( P� �                               PU� �                              � PQ� p                               Q PQ� `
                               } TQ��                        @@   � U��
�                             ��`U��*�                             ��rU��:�/                               l�n�W���/ @@                        X�n����?                            @  W�{���꫿  @                       @   V�j����j�   @@                         U�n����j�                             V�~����k�  @                      @ D PV�k����j�
                             �U�ju��j�+                          �U�~U���k��                          @�V�nUU��j��                       @  ��V�kUU����
                          d�U�zUT����[)                        ��U�nUT����k�                          i�V��UT�꪿[�                           ��V��T��k���                           ��U�^T��j��*                       ��U�[yTn����
                           ��V�V�U[���                          �V�V��V���*                             �^�U��V���                          �zeU��V���                               �uU��V��; @@                          �U��V��                             �nQ����                              �jP����                         �zP���/                             �zP�����                            @�jХ����                             ��j��֯��                         @��j5��լ��/                            ��j	�����?                           ��j	�����/ @@                          ��j��@��                        @ @ ��  �  �                             �   U  ��                               �   (                              � �?   @                            � �?                                  � �  @                          @  �
* ��                              �
* ��                              �� j�
                                 �Zj ��@                            ��j ��                                P�Z �� @                            P�Z ��                              P�V �j                               P�U UZ                                 @U TU                                 U PU                                   U PU  @                                T @ @                                 P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ����      @            @            @            @            @            @            UU           U            U            U            U           U        P U U      P U A      P U A      PTUTA      TU  A      TU  A     @TUU  UA    @  T   @    @  T   @    @ T   @    @ T        @ T        @ T        U TU    P   A TU        A TU      PUA TU    TUTA TU     @TA TU     @TA  U     @TA  U     @PUA T@    TU  A T@       A T@       UPUU   P   @PUU        @PUU        @PUU@ @      TU@ @       TU@ @       TU@ @     @ TU@ @    @ TU@      @ TU@      UPU    P   APU        APUU T     APU      APU      UUUUPTUP   @  @  @    @  @  @    @  @  @       U             A   A        TA TA                                                         TA TA       TA TA       TA TA       TU TU       TU TU       TU TU        U   U         U   U         U   U          @            @            @            @            @            @            U�
           U�
           U�
           U�
           U�
           U�
        P U�
 �      P U�
 �      P U�
 �      TU��A      TU��A      TU��A     @��VU��VA    @��V*�@    @��V*�@    @��V*�@    @��V*�     @��V*�     @��V*�     j��VU���j   j��VU���*   j��VU���* �Vj��VU���*�V�Vj��VU���*�B�Vj��VU���*�B�Vj��U�
 �*�B�Vj��U�
 �*�B�Vj��VU�
 �*�V  j�
T@��*   j�
T@��*   j�ZUU����j   @�ZUU����*    @�ZUU����*    @�ZUU@���*     �
TU@��B      �
TU@��B      �
TU@��B     @�
TU@���*    @�
TU@���*    @�
TU@���*    j�Z�U�
��j   j�Z�U�
��*   j�Z�U�Z��*   j�ZU�
��*   j�ZU�
��*   j�ZU�
��j   @  @  �*    @  @  �*    @  @  �*       U             A   A        ��* ��*       ��* ��*       ��* ��*       ��* ��*       ��* ��*       ��* ��*       T� T�       T� T�       T� T�       TU TU       TU TU       TU TU        U   U         U   U         U   U          @            @            @            @            @            @            U�
           U�
           U�
           U�
           U�
           U�
        P U�
 �      P U�
 �      P U�
 �      �TU���      �TU���      �TU���     ���VU����    ���V����    ���V����    @��V����?    @��V����?    @��V����?    @��V����?    j��VU�����   j��VU�����   j��VU����� �Vj��VU�������Vj��VU�������Vj��VU�������Vj���U�������Vj���U�������Vj���U������  j��Wկ���   j��Wկ���   j��Wկ���   @�ZUտ���*    @�ZUտ���*    @�ZU����*     �
T����      �
T����      �
T����     @�
T����*    @�
T����*    @�
T����*    j�Z�տ����   j�Z�տ����   j�Z�տ����   j�Zտ
���   j�Zտ
���   j�Zտ
���   @  �?  �*    @  �?  �*    @  �?  �*       �             �   �        ��* ��*       ��* ��*       ��* ��*       ��* ��*       ��* ��*       ��* ��*       T� T�       T� T�       T� T�       TU TU       TU TU       TU TU        U   U         U   U         U   U    (c)1992Thin Chen Enter. � ��@���������`�����[������ds���s������ k� %������������si<�s��`

�� �c�� � �����`� �/ ������`������@�]�<��8�� k��i0��i �������������i0���i ��������  դ���a�1�]�-�D k�����ȑ�� ��� ��i0��i ���ߩ��� ���_��a�Ș N����a�����`��`�����`���M�]�I��8�� k��i��i ��i0��i �������������i0���i �������� դ���a�1�]�-�D k���ȱ����'��� ��i0��i ���ߩ�����a�����`��`



}����i ��J��� k��
�e��i ������`�� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 ���  ��� � � � � � �� � �( ���򩧅��� b��@�d�� �������`��������� 7��s)��������)�S����L������������� !��������� ������i !���LƧ@@@@@@8  0@P`8@@@@@@p�����Т ���	��8��������p����	��i��������������i����ɀ�L]�ds�sɴ��  ����  ����`

��o����p����q����r���������i����������i����� ��������`	
+,)*78'(56%&34#$12!"/0 -.                   P @  T   @  @@@@ UPUTUTTUPU@U UUUUUUU          @ T U@UPUPTTUUUQPPP T@UPUTUTUUU U UUTPP  UUUUUUUUUUPPPPPPUU UPUTUTUUUUUUUUUUUUUU    UUUUUUUUUUUUUUU@U@U@UAUEUEUUUUUT @   P@@@@  @  T P @    UUUUUUU UUUTUUU TUTUUUUUUUUUUUPPPPPUUUTTUPU@U T  PPTUUU  UUUUUUUUUUPPPPPPPUUUUUUUUUUUUUUUUUU    UUUUUUUUUQUAUUUUUUUUUUUUUUTUPU@U   � 
�    �((  * �   * ���� ������*������ �������     
 *    � � ������*�*�*�*�*�*�*�*�*�* ��������
���
 � ��
�
�*�*  �����������*�*�*�*�*�*�*�* ����������������*�*�*�*�*    �*��*�����������������������������(( (  �  
 �*�� ��    �*  � � �    ������� ��
�*�*�*�
� �������
�
�
�
�
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*�����������������*�*    �*�*�*�*�����������������������������s)����`����������0'� �����������������Z ��z�����۠ �������������������Z ��z�����ة ��`��������������������� k���JJe��i ����



e��i ��JJJJe���)�������������
.�.�
.�.����Q�ȭ�Q�ȭ�Q��i0��i ��i��i ����L �`es�s��`� �����`H)�����hJJJJ�
ei@}���` 0`��� P���@p��      
�*�*�*�*�*�*�*�*����
������ �  �*�*�
�
�� 
 ����������*�*�*�*�*�*�*�*���������+6]
		XCHG	AX,SI
		MOV	AX,DATA_129[SI]
		CMP	AX,[BP+0AH]
		JNE	SHORT LOC_2178
		LES	BX,DWORD PTR [BP-10H]
		MOV	AX,ES:[BX+6]
		MOV	DATA_129[SI],AX
LOC_2178:
		PUSH	WORD PTR [BP+0AH]
		PUSH	WORD PTR [BP+8]
;*		CALL	FAR PTR SUB_7		;*
		DB	 9AH, 7DH, 00H, 00H, 00H
		MOV	DATA_246,0
		MOV	AX,[BP-0CH]
		MOV	DX,[BP-0AH]
		MOV	[BP-4],AX
		MOV	[BP-2],DX
		MOV	AX,[BP-4]
		MOV	DX,[BP-2]
		MOV	SP,BP
		POP	BP
		RETF	6
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		SUB	SP,4
		nop	                        ;*ASM fixup - sign extn byte
		MOV	SP,BP
		POP	BP
		RETF
			                        ;* No entry point to code
		ADD	[DI-75H],DL
		IN	AL,DX			; port 0, DMA-1 bas&add ch 0
		MOV	AH,0FH
		INT	10H			; Video display   ah=functn 0Fh
						;  get state, al=mode, bh=page
						;   ah=columns on screen
		XOR	AH,AH
		POP	BP
		RETF
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		XOR	AX,AX
		MOV	ES,AX
		MOV	AH,ES:equip_bits_
		MOV	AL,[BP+6]
		CMP	AL,7
		JNE	SHORT LOC_2179
		OR	AH,30H			; '0'
		JMP	SHORT LOC_2180
LOC_2179:
		AND	AH,0CFH
		OR	AH,20H			; ' '
LOC_2180:
		MOV	ES:equip_bits_,AH
		XOR	AH,AH
		INT	10H			; Video display   ah=functn 00h
						;  set display mode in al
		MOV	AH,5
		XOR	AL,AL
		INT	10H			; Video display   ah=functn 05h
						;  set display page al
		POP	BP
		RETF	2
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	AX,1111H
		MOV	BX,[BP+6]
		CMP	BL,6
		JNE	SHORT LOC_2181
		MOV	AL,12H
LOC_2181:
		MOV	BL,0
		INT	10H			; Video display   ah=functn 11h
						;  load 8x8 font, bl=block
		POP	BP
		RETF	2
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	AH,0BH
		MOV	BH,0
		MOV	BL,[BP+6]
		INT	10H			; Video display   ah=functn 0Bh
						;  set color from bx (CGA modes)
		POP	BP
		RETF	2
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	DH,[BP+8]
		DEC	DH
		MOV	DL,[BP+6]
		DEC	DL
		XOR	BX,BX
		MOV	AH,2
		INT	10H			; Video display   ah=functn 02h
						;  set cursor location in dx
		POP	BP
		RETF	4
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		XOR	AX,AX
		MOV	ES,AX
		MOV	DL,ES:video_options_
		MOV	DH,DL
		OR	DH,1
		MOV	ES:video_options_,DH
		MOV	CH,[BP+8]
		MOV	CL,[BP+6]
		MOV	AH,1
		INT	10H			; Video display   ah=functn 01h
						;  set cursor mode in cx
		MOV	ES:video_options_,DL
		POP	BP
		RETF	4
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	DH,[BP+8]
		DEC	DH
		MOV	DL,[BP+6]
		DEC	DL
		XOR	BX,BX
		MOV	AH,2
		INT	10H			; Video display   ah=functn 02h
						;  set cursor location in dx
		XOR	BX,BX
		MOV	AH,8
		INT	10H			; Video display   ah=functn 08h
						;  get char al & attrib ah @curs
		POP	BP
		RETF	4
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	DH,[BP+0AH]
		DEC	DH
		MOV	DL,[BP+8]
		DEC	DL
		XOR	BX,BX
		MOV	AH,2
		INT	10H			; Video display   ah=functn 02h
						;  set cursor location in dx
		MOV	AX,[BP+6]
		MOV	BL,AH
		XOR	BH,BH
		MOV	CX,1
		MOV	AH,9
		INT	10H			; Video display   ah=functn 09h
						;  set char al & attrib bl @curs
						;   cx=# of chars to replicate
		POP	BP
		RETF	6
			                        ;* No entry point to code
		MOV	DI,CX
		MOV	CX,1
		MOV	BH,0
LOC_2182:
		AND	DI,DI
		JLE	SHORT LOC_2183
		MOV	AH,2
		INT	10H			; Video display   ah=functn 02h
						;  set cursor location in dx
		LODSB
		MOV	AH,9
		INT	10H			; Video display   ah=functn 09h
						;  set char al & attrib bl @curs
						;   cx=# of chars to replicate
		INC	DL
		DEC	DI
		JMP	SHORT LOC_2182
LOC_2183:
		RETF
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	CX,[BP+6]
		AND	CX,CX
		JLE	SHORT LOC_2189
		TEST	BYTE PTR DATA_254,0FFH
		JNZ	SHORT LOC_2188
		MOV	AX,[BP+0EH]
		DEC	AX
		IMUL	DATA_264
		ADD	AX,[BP+0CH]
		DEC	AX
		MOV	DI,AX
		SHL	DI,1
		CLD
		MOV	SI,[BP+8]
		MOV	ES,DATA_263
		MOV	AH,[BP+0AH]
		MOV	DX,DATA_262
		AND	DX,DX
		JZ	SHORT LOCLOOP_2187

LOCLOOP_2184:
		LODSB
		MOV	BX,AX
LOC_2185:
		IN	AL,DX			; port 5500H ??I/O NON-STANDARD
		TEST	AL,1
		JNZ	LOC_2185
		CLI
LOC_2186:
		IN	AL,DX			; port 5500H ??I/O NON-STANDARD
		TEST	AL,1
		JZ	LOC_2186
		MOV	AX,BX
		STOSW
		STI
		LOOP	LOCLOOP_2184

		JMP	SHORT LOC_2189

LOCLOOP_2187:
		LODSB
		STOSW
		LOOP	LOCLOOP_2187

		JMP	SHORT LOC_2189
LOC_2188:
		MOV	BL,[BP+0AH]
		MOV	DH,[BP+0EH]
		DEC	DH
		MOV	DL,[BP+0CH]
		DEC	DL
		MOV	SI,[BP+8]
;*		CALL	FAR PTR SUB_623		;*
		DB	 9AH,0ECH, 00H, 05H, 01H
LOC_2189:
		POP	BP
		RETF	0AH
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	AX,0B000H
		MOV	ES,AX
		XOR	SI,SI
		MOV	AL,ES:[SI]
		MOV	AH,AL
		ADD	AH,5AH			; 'Z'
		MOV	ES:[SI],AH
		MOV	BH,ES:[SI]
		MOV	CL,0
		CMP	AH,BH
		JNE	SHORT LOC_2190
		MOV	CL,0FFH
LOC_2190:
		MOV	DI,[BP+0AH]
		MOV	[DI],CL
		MOV	ES:[SI],AL
		MOV	AX,0B800H
		MOV	ES,AX
		MOV	AL,ES:[SI]
		MOV	AH,AL
		ADD	AH,5AH			; 'Z'
		MOV	ES:[SI],AH
		MOV	BH,ES:[SI]
		MOV	CL,0
		CMP	AH,BH
		JNE	SHORT LOC_2191
		MOV	CL,0FFH
LOC_2191:
		MOV	DI,[BP+8]
		MOV	[DI],CL
		MOV	ES:[SI],AL
		MOV	AH,12H
		MOV	BL,10H
		INT	10H			; Video display   ah=functn 12h
						;  EGA/VGA special, bl=function
		MOV	AL,CL
LOC_2192:
		MOV	CL,0
		MOV	CH,0FFH
		MOV	DI,[BP+6]
		MOV	[DI],CL
		MOV	DI,[BP+0CH]
		MOV	[DI],CL
		MOV	SI,[BP+0EH]
		MOV	[SI],CL
		CMP	BL,10H
		JE	SHORT LOC_2195
		MOV	[DI],CH
		CMP	BH,0
		JNE	SHORT LOC_2193
		MOV	DI,[BP+8]
		MOV	[DI],CH
		MOV	DI,[BP+6]
		MOV	[DI],CH
		JMP	SHORT LOC_2194
LOC_2193:
		CMP	BH,1
		JNE	SHORT LOC_2194
		MOV	DI,[BP+0AH]
		MOV	[DI],CH
LOC_2194:
		AND	AL,0FH
		MOV	BX,204H
DATA_192	DW	0D72EH
DATA_193	DW	488H			; Data table (indexed access)
LOC_2195:
		POP	BP
		RETF	0AH
			                        ;* No entry point to code
		ADD	[BX+SI],AL
		ADD	BH,BH
		DB	0FFH,0FFH
DATA_194	DW	0			; Data table (indexed access)
		DB	 00H,0FFH,0FFH,0FFH
DATA_195	DW	0			; Data table (indexed access)
		DB	 00H, 00H, 55H, 8BH
DATA_196	DW	0B4ECH			; Data table (indexed access)
		DB	 0FH,0CDH, 10H, 8AH
DATA_197	DW	0B4C4H			; Data table (indexed access)
		DB	 00H,0A3H, 4EH,0EBH,0B4H, 12H
		DB	0B3H, 10H,0CDH, 10H
DATA_198	DW	0FB80H			; Data table (indexed access)
		DB	 10H, 74H, 10H,0B8H, 30H, 11H
		DB	0CDH, 10H,0B6H, 00H
DATA_199	DW	8942H			; Data table (indexed access)
		DB	 16H, 50H,0EBH, 88H, 0EH, 5AH
		DB	0EBH, 5DH,0CBH, 00H

;��������������������������������������������������������������������������
;                              SUBROUTINE
;��������������������������������������������������������������������������

SUB_930		PROC	NEAR
DATA_200	DW	0C923H			; Data table (indexed access)
		DB	 7EH, 1DH,0F6H,0C6H, 80H, 75H
		DB	 1EH, 23H,0D2H
		DB	74H
DATA_201	DW	0AC15H			; Data table (indexed access)
		DB	 8BH,0D8H
LOC_2196:
		IN	AL,DX			; port 0, DMA-1 bas&add ch 0
		TEST	AL,1
		JNZ	LOC_2196
		CLI
LOC_2197:
		IN	AL,DX			; port 0, DMA-1 bas&add ch 0
		TEST	AL,1
		JZ	LOC_2197
		MOV	AX,BX
		STOSW
DATA_203	DW	0E2FBH, 0C3ECH
LOC_2199:
DATA_205	DW	0ABACH
DATA_206	DW	0FCE2H
DATA_207	DW	8AC3H
DATA_208	DD	9AD78BDCH
DATA_210	DW	0ECH, 0
DATA_212	DW	0FA8BH
DATA_213	DW	80B6H, 8BC3H
DATA_215	DW	0C4EH, 0C13BH
DATA_217	DW	1A7DH, 0C82BH
DATA_219	DW	0CB3BH
DATA_220	DW	27EH
DATA_221	DW	0CB8BH
DATA_222	DW	5350H
DATA_223	DW	8A51H
DATA_224	DW	866H
DATA_225	DW	0B3E8H
DATA_226	DW	59FFH
DATA_227	DW	585BH
DATA_229	DB	3
DATA_230	DB	0C1H
DATA_231	DW	0D92BH
DATA_233	DW	347EH
		DB	 8BH, 4EH, 0AH, 3BH,0C1H
LOC_2201:
		JG	SHORT LOC_2203
		CMP	AX,[BP+0CH]
		JL	SHORT LOC_2203
		SUB	CX,AX
		INC	CX
		CMP	CX,BX
		JLE	SHORT LOC_2202
		MOV	CX,BX
LOC_2202:
		PUSH	AX
		PUSH	BX
		PUSH	CX
		MOV	AH,[BP+6]
		CALL	SUB_930
		POP	CX
		POP	BX
		POP	AX
		ADD	AX,CX
		SUB	BX,CX
		JLE	SHORT LOC_2204
LOC_2203:
		CMP	AX,[BP+0AH]
		JLE	SHORT LOC_2204
		MOV	CX,BX
		MOV	AH,[BP+8]
		CALL	SUB_930
LOC_2204:
DATA_235	DW	55C3H			; Data table (indexed access)
		DB	 8BH,0ECH, 1EH, 8BH, 46H, 0EH
		DB	 48H, 36H,0F7H, 2EH, 4EH,0EBH
		DB	 03H, 46H, 10H, 48H, 8BH,0F8H
		DB	0D1H,0E7H,0FCH, 36H, 8EH, 06H
		DB	 4CH,0EBH, 36H, 8BH, 16H, 4AH
		DB	0EBH, 36H,0F6H, 06H, 22H,0EBH
		DB	0FFH, 74H, 0EH, 8AH, 76H, 0EH
		DB	0FEH,0CEH, 8AH, 56H, 10H,0FEH
		DB	0CAH, 8BH,0FAH,0B6H, 80H
LOC_2205:
		MOV	BX,[BP+16H]
		CMP	BX,1
		JLE	SHORT LOC_2206
		MOV	AX,1
		DEC	BX
		LDS	SI,DWORD PTR [BP+18H]
;*		CALL	SUB_931			;*
		DB	0E8H, 62H,0FFH
LOC_2206:
		MOV	BX,[BP+14H]
		AND	BX,BX
		JLE	SHORT LOC_2207
		MOV	AX,[BP+16H]
		LDS	SI,DWORD PTR [BP+1CH]
DATA_237	DB	0E8H
		DB	52H
DATA_238	DW	8BFFH
		DB	 46H, 16H, 03H, 46H, 14H, 8BH
		DB	 5EH, 12H, 3BH,0C3H, 7FH, 09H
		DB	 2BH,0D8H, 43H,0C5H, 76H, 18H
		DB	0E8H, 3CH,0FFH
LOC_2208:
		POP	DS
		POP	BP
		RETF	1AH
SUB_930		ENDP

			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		PUSH	DS
		MOV	CX,7FFFH
		MOV	SI,[BP+6]
		MOV	SI,[SI]
		AND	SI,SI
		JZ	SHORT LOC_2211
		MOV	DI,[BP+8]
		MOV	DX,[DI]
		MOV	CX,[BP+0EH]
		SUB	CX,DX
		JL	SHORT LOC_2209
		MOV	BL,4
		JMP	SHORT LOC_2210
LOC_2209:
		NEG	CX
		MOV	BL,8
LOC_2210:
		MOV	DS,SI
		CMP	CX,4
		JL	SHORT LOC_2213
LOC_2211:
		MOV	AX,[BP+0EH]
		CMP	AX,CX
		JGE	SHORT LOC_2212
		MOV	CX,AX
		XOR	DX,DX
		MOV	BL,4
		MOV	DS,[BP+0AH]
LOC_2212:
		MOV	DI,[BP+0CH]
		ADD	DI,2
		MOV	AX,DI
		SUB	AX,[BP+0EH]
		CMP	AX,CX
		JGE	SHORT LOC_2213
		MOV	DX,DI
		MOV	BL,8
		MOV	DS,[BP+0AH]
LOC_2213:
		MOV	DI,[BP+0EH]
		CMP	BL,4
		JNE	SHORT LOC_2216
		XOR	BX,BX
LOC_2214:
		CMP	DX,DI
		JGE	SHORT LOC_2219
		MOV	AL,[BX+2]
		CMP	AL,3
		JNE	SHORT LOC_2215
		MOV	AL,[BX+3]
		XOR	AH,AH
		ADD	AX,DX
		CMP	AX,DI
		JG	SHORT LOC_2219
		MOV	DX,AX
		MOV	DS,[BX+6]
DATA_241	DW	0E3EBH
LOC_2215:
DATA_242	DW	8E42H			; Data table (indexed access)
DATA_243	DW	65FH			; Data table (indexed access)
		DB	0EBH,0DDH
LOC_2216:
		XOR	BX,BX
LOC_2217:
		CMP	DX,DI
		JLE	SHORT LOC_2219
		MOV	DS,[BX+0AH]
		MOV	AL,[BX+2]
		CMP	AL,3
		JNE	SHORT LOC_2218
		MOV	AL,[BX+3]
		XOR	AH,AH
		SUB	DX,AX
		JMP	SHORT LOC_2217
LOC_2218:
		DEC	DX
DATA_248	DW	0E6EBH
LOC_2219:
DATA_249	DW	7E8BH
DATA_250	DW	3608H
DATA_251	DW	1589H
DATA_252	DB	8CH
		DB	0DAH
DATA_253	DB	33H
		DB	0C0H
DATA_254	DB	1FH
		DB	8BH
DATA_255	DW	676H
DATA_256	DW	1489H
DATA_257	DW	0CA5DH
DATA_258	DW	0AH
DATA_259	DW	8B55H
		DB	0ECH, 8BH, 4EH, 06H, 23H,0C9H
		DB	 7EH, 11H
DATA_260	DW	8E1EH
DATA_261	DW	0A46H
		DB	 8BH, 7EH, 08H, 8BH, 76H, 0CH
		DB	 8EH, 5EH, 0EH,0FCH,0F3H,0A4H
		DB	 1FH
LOC_2220:
		POP	BP
		RETF	0AH
			                        ;* No entry point to code
		PUSH	BP
DATA_263	DW	0EC8BH
DATA_264	DW	4E8BH
DATA_265	DW	2306H
DATA_266	DW	7EC9H
DATA_268	DW	1E0BH
		DB	 07H, 8BH, 46H, 08H
DATA_270	DW	7E8BH
DATA_271	DW	0FC0AH
DATA_273	DW	0AAF3H
DATA_275	DW	0CA5DH
DATA_277	DW	6
DATA_279	DW	8B55H
DATA_281	DW	8BECH			; Data table (indexed access)
DATA_283	DW	84EH			; Data table (indexed access)
DATA_284	DW	0C923H			; Data table (indexed access)
DATA_285	DW	2C7EH			; Data table (indexed access)
DATA_286	DW	71EH			; Data table (indexed access)
DATA_287	DW	768BH			; Data table (indexed access)
DATA_288	DW	8B0AH
DATA_289	DW	0FCFEH			; Data table (indexed access)
DATA_290	DW	61BBH			; Data table (indexed access)
DATA_291	DW	0BA7AH			; Data table (indexed access)
DATA_292	DW	5A41H			; Data table (indexed access)
DATA_293	DB	8AH
		DB	66H
DATA_294	DW	2206H
DATA_295	DW	75E4H
		DB	 02H, 87H,0DAH

LOCLOOP_2221:
		LODSB
		CMP	AL,BL
DATA_296	DW	0D7CH
DATA_297	DW	0C73AH
		DB	 7FH, 09H, 2AH,0C3H, 02H,0C2H
DATA_298	DB	0AAH
		DB	0E2H
DATA_299	DW	0EBF0H
DATA_300	DW	4703H
		DB	0E2H,0EBH
LOC_2223:
		POP	BP
		RETF	6
DATA_301	DW	8B55H
DATA_302	DW	33ECH
		DB	0DBH, 8BH, 4EH, 08H, 23H,0C9H
DATA_303	DB	7EH
		DB	42H
DATA_304	DW	0F983H
DATA_305	DW	7502H
		DB	 28H, 8BH, 76H, 0AH
DATA_306	DW	8AACH
DATA_307	DW	0ACE0H
DATA_308	DW	0FC80H
		DB	 41H, 7CH, 08H, 80H,0FCH, 5AH
DATA_309	DB	7FH
		DB	3
DATA_310	DW	0C480H
DATA_311	DW	3C20H
		DB	 41H, 7CH
DATA_312	DW	3C06H
		DB	 5AH, 7FH
DATA_313	DW	402H
DATA_314	DW	0F620H
		DB	0E4H, 25H, 7FH, 00H, 8BH, 7EH
DATA_315	DB	6
		DB	89H
DATA_316	DW	8B05H
DATA_317	DW	0A76H

LOCLOOP_2226:
		LODSB
		CMP	AL,41H			; 'A'
		JL	SHORT LOC_2227
		CMP	AL,5AH			; 'Z'
		JG	SHORT LOC_2227
		ADD	AL,20H			; ' '
LOC_2227:
		ADD	BL,AL
		LOOP	LOCLOOP_2226

		AND	BL,7FH
DATA_322	DW	0C38BH
DATA_323	DW	0CA5DH
		DB	6, 0
DATA_324	DW	8B55H
DATA_325	DW	8BECH
DATA_326	DW	64EH
DATA_327	DW	0C923H
		DB	 7EH, 1BH, 8BH, 76H, 0AH, 8BH
DATA_328	DB	7EH
		DB	8

LOCLOOP_2228:
DATA_329	DW	8AACH
DATA_330	DW	471DH
		DB	 3AH,0C3H
DATA_331	DW	774H
		DB	 80H,0EBH
DATA_332	DW	3A20H
DATA_333	DW	75C3H
		DB	 06H,0E2H,0EFH,0B0H, 01H,0EBH
DATA_334	DB	2
LOC_2229:
		XOR	AX,AX
LOC_2230:
		POP	BP
DATA_336	DW	6CAH
		DB	 00H, 55H, 8BH,0ECH, 8BH, 5EH
DATA_337	DW	8B06H
DATA_338	DW	0AC36H
		DB	0EEH, 03H, 76H, 0AH, 8AH, 66H
DATA_339	DB	8
		DB	0AH
DATA_340	DW	74E4H
DATA_341	DW	0FE14H
		DB	0CCH,0ACH
DATA_342	DW	413CH
		DB	 7CH, 06H
DATA_343	DW	5A3CH
DATA_344	DW	277H
		DB	 04H, 20H
LOC_2231:
		CMP	AL,[BX]
		JNE	SHORT LOC_2234
DATA_345	DW	0EB43H
DATA_346	DW	0ACE8H
		DB	 3CH, 20H, 74H, 04H, 3CH, 5DH
		DB	 75H, 05H
LOC_2233:
		MOV	AX,1
		JMP	SHORT LOC_2235
LOC_2234:
		XOR	AX,AX
LOC_2235:
		POP	BP
		RETF	6
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		PUSH	DS
		POP	ES
		MOV	AX,[BP+0EH]
		MOV	BX,[BP+8]
		MOV	DX,[BP+0CH]
		CLD
LOC_2236:
		MOV	SI,AX
		MOV	DI,BX
		MOV	CX,[BP+6]
		REPE	CMPSB
		JZ	SHORT LOC_2237
		CMP	AX,DX
		JE	SHORT LOC_2238
		ADD	AX,[BP+0AH]
		JMP	SHORT LOC_2236
LOC_2237:
		SUB	AX,[BP+0EH]
		JMP	SHORT LOC_2239
LOC_2238:
		MOV	AX,3E7H
LOC_2239:
		POP	BP
		RETF	0AH
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		XOR	AH,AH
		INT	16H			; Keyboard i/o  ah=function 00h
						;  get keybd char in al, ah=scan
		POP	BP
		RETF
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	AH,1
		INT	16H			; Keyboard i/o  ah=function 01h
						;  get status, if zf=0  al=char
DATA_348	DW	275H
		DB	 33H,0C0H, 5DH,0CBH, 55H, 8BH
		DB	0ECH, 33H,0D2H,0B4H, 02H,0CDH
		DB	 17H, 80H,0E4H, 09H, 75H, 0CH
		DB	 8AH, 46H, 06H, 32H,0E4H,0CDH
		DB	 17H, 80H,0E4H, 09H, 74H, 05H
LOC_2240:
		MOV	AX,1
		JMP	SHORT LOC_2242
LOC_2241:
		XOR	AX,AX
LOC_2242:
		POP	BP
		RETF	2
			                        ;* No entry point to code
		MOV	BX,BP
		MOV	BP,SP
		MOV	AX,[BP+4]
		AND	AX,AX
		JNZ	SHORT LOC_2243
		MOV	AX,[BP+2]
		MOV	DATA_384,AX
		MOV	AX,[BP]
		MOV	DATA_385,AX
		MOV	DATA_386,BX
		MOV	DATA_387,SP
		MOV	BP,BX
		RETF	2
LOC_2243:
		MOV	SP,DATA_387
		MOV	BP,SP
		MOV	AX,DATA_385
		MOV	[BP],AX
		MOV	AX,DATA_384
		MOV	[BP+2],AX
		MOV	BP,DATA_386
		RETF	2
			                        ;* No entry point to code
		MOV	AL,0B6H
		OUT	43H,AL			; port 43H, 8253 wrt timr mode
		MOV	AX,533H
		OUT	42H,AL			; port 42H, 8253 timer 2 spkr
		MOV	AL,AH
		OUT	42H,AL			; port 42H, 8253 timer 2 spkr
		MOV	AL,4FH			; 'O'
		OUT	61H,AL			; port 61H, 8255 B - spkr, etc
						;  al = 4FH, speaker on
		MOV	CX,32C8H

LOCLOOP_2244:
		LOOP	LOCLOOP_2244

		MOV	AL,4DH			; 'M'
		OUT	61H,AL			; port 61H, 8255 B - spkr, etc
						;  al = 4DH, enable keyboard
		RETF
LOC_2245:
		MOV	AH,1
		INT	16H			; Keyboard i/o  ah=function 01h
						;  get status, if zf=0  al=char
		JZ	SHORT LOC_2246
		XOR	AH,AH
		INT	16H			; Keyboard i/o  ah=function 00h
						;  get keybd char in al, ah=scan
		JMP	SHORT LOC_2245
LOC_2246:
		RETF
		DB	1, 0, 2, 0
DATA_349	DW	3
		DB	 04H, 00H, 55H, 8BH,0ECH
DATA_350	DB	0B4H
DATA_351	DW	2E35H
DATA_352	DW	20A0H
DATA_353	DW	0CD06H
		DB	 21H, 33H,0C0H, 26H, 81H, 7FH
		DB	 02H, 50H, 45H, 75H, 11H, 26H
		DB	 81H, 7FH, 04H, 32H, 69H, 75H
		DB	 09H, 26H, 81H, 7FH, 06H, 6EH
		DB	 74H, 75H, 01H
		DB	48H
LOC_2247:
		POP	BP
		RETF
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		PUSH	DS
		LEA	DX,[BP+6]
		INT	67H			; ??INT NON-STANDARD INTERRUPT
		POP	DS
		POP	BP
		RETF	14H
			                        ;* No entry point to code
		ADD	AX,600H
		ADD	[BX],AL
		ADD	[BX+SI],CL
		ADD	[BP],AH
		ADD	[DI-75H],DL
		IN	AL,DX			; port 0, DMA-1 bas&add ch 0
		MOV	AH,35H			; '5'
		MOV	AL,CS:DATA_60
		INT	21H			; DOS Services  ah=function 35h
						;  get intrpt vector al in es:bx
		MOV	SI,[BP+8]
		MOV	[SI],ES
		MOV	SI,[BP+6]
		MOV	[SI],BX
		MOV	CS:DATA_61,DS
		PUSH	DS
		PUSH	CS
		POP	DS
DATA_356	DW	85BAH
		DB	 06H,0B4H, 25H, 2EH
DATA_357	DB	0A0H
		DB	 2EH, 06H,0CDH
DATA_358	DW	1F21H
DATA_359	DW	0CA5DH
DATA_360	DW	4
		DB	 09H, 00H, 0AH, 00H, 0BH, 00H
		DB	 0CH, 00H, 55H, 8BH,0ECH, 1EH
		DB	 8BH, 56H, 06H, 8EH, 5EH, 08H
		DB	0B4H, 25H, 2EH,0A0H, 2EH, 06H
		DB	0CDH, 21H, 1FH, 5DH,0CAH, 04H
		DB	 00H, 0DH, 00H, 0EH, 00H, 0FH
		DB	 00H, 10H, 00H, 1EH, 2EH, 8EH
		DB	 1EH, 2FH, 06H, 50H, 9AH, 63H
		DB	 08H, 00H, 00H, 1FH,0CFH, 11H
		DB	 00H, 12H, 00H, 13H, 00H, 14H
		DB	 00H, 15H, 00H, 16H, 00H, 17H
		DB	 00H, 18H, 00H, 00H, 55H, 8BH
		DB	0ECH, 33H,0C0H, 8BH
		DB	76H
DATA_361	DB	6
DATA_362	DB	0B9H
		DB	 40H, 00H

LOCLOOP_2248:
		ADD	AX,[SI]
		ADD	AX,[SI+2]
		ADD	AX,[SI+4]
		ADD	AX,[SI+6]
		ADD	SI,8
		LOOP	LOCLOOP_2248

		POP	BP
		RETF	2
			                        ;* No entry point to code
		PUSH	BP
DATA_366	DW	0EC8BH
		DB	 8DH, 3EH, 50H,0EFH, 1EH, 07H
		DB	0B9H, 81H, 00H,0FCH, 33H,0C0H
		DB	0F3H,0AEH, 23H,0C9H, 74H, 22H
		DB	 4FH, 8BH,0C7H, 8DH, 0EH, 50H
		DB	0EFH, 2BH,0C1H,0B1H, 03H,0D3H
		DB	0E0H, 8AH, 15H,0BBH, 00H, 01H
LOC_2249:
		MOV	DH,DL
		AND	DH,BH
		JNZ	SHORT LOC_2250
		SHL	BH,1
		INC	BL
		JMP	SHORT LOC_2249
LOC_2250:
		XOR	BH,BH
		ADD	AX,BX
LOC_2251:
		POP	BP
		RETF
			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	AX,[BP+6]
		MOV	BX,8
		XOR	DX,DX
		DIV	BX
		LEA	DI,CS:[0EF50H]
DATA_368	DB	3
DATA_369	DB	0F8H
		DB	0B3H, 01H, 8AH
DATA_370	DB	0CAH
		DB	0D2H
DATA_371	DW	8AE3H
DATA_372	DW	3205H
		DB	0C3H, 88H, 05H, 5DH,0CAH, 02H
		DB	 00H, 00H

;��������������������������������������������������������������������������
;                              SUBROUTINE
;��������������������������������������������������������������������������

SUB_932		PROC	NEAR
		CMP	SI,BX
		JB	SHORT LOC_2253
		PUSH	AX
		PUSH	DX
		PUSH	DI
		PUSH	ES
		PUSH	BP
;*		CALL	FAR PTR SUB_1		;*
		DB	 9AH, 01H, 00H, 00H, 00H
		MOV	CX,AX
		POP	ES
		POP	DI
		POP	DX
		POP	AX
		MOV	SI,[BP+0AH]
		MOV	BX,SI
		ADD	BX,[BP+0CH]
		AND	CX,CX
		JZ	SHORT LOC_2252
		MOV	AH,CL
LOC_2252:
		CMP	SI,BX
		JB	SHORT LOC_2253
		MOV	AL,1AH
		MOV	BYTE PTR [BP+5],0FFH
		RETN
LOC_2253:
		TEST	BYTE PTR [BP+5],0FFH
		JZ	SHORT LOC_2254
		MOV	AL,1AH
		RETN
LOC_2254:
		LODSB
		CMP	AL,1AH
		JNE	SHORT LOC_2255
		MOV	BYTE PTR [BP+5],0FFH
LOC_2255:
		RETN
SUB_932		ENDP

			                        ;* No entry point to code
		PUSH	BP
		MOV	BP,SP
		MOV	BP,[BP+6]
		MOV	SI,[BP+0AH]
		MOV	BX,SI
		ADD	SI,[BP+6]
DATA_374	DW	34EH			; Data table (indexed access)
		DB	 5EH, 0CH,0E8H,0ABH,0FFH, 3CH
		DB	 0AH, 75H, 03H,0E8H,0A4H,0FFH
LOC_2256:
		CMP	AL,1AH
		JNE	SHORT LOC_2257
		MOV	AH,1
		JMP	SHORT LOC_2263
LOC_2257:
		PUSH	DS
		POP	ES
		MOV	DI,WORD PTR DS:[0EEACH]
		INC	DI
		XOR	DX,DX
		MOV	AH,0
LOC_2258:
		CMP	AL,0DH
		JE	SHORT LOC_2262
		CMP	AL,1AH
		JE	SHORT LOC_2262
		CMP	AL,9
		JNE	SHORT LOC_2259
		TEST	BYTE PTR [BP+4],0FFH
		JZ	SHORT LOC_2259
		MOV	CX,DX
		AND	CX,0FFF8H
		nop	                        ;*ASM fixup - sign extn byte
		ADD	CX,8
		MOV	AL,20H			; ' '
		CMP	DX,CX
		JGE	SHORT LOC_2261
		CMP	DX,0FFH
		JGE	SHORT LOC_2261
		STOSB
		INC	DX
DATA_376	DW	0F2EBH
LOC_2259:
		CMP	DX,0FFH
		JGE	SHORT LOC_2260
		INC	DX
		STOSB
		JMP	SHORT LOC_2261
LOC_2260:
		MOV	AH,3
LOC_2261:
		CALL	SUB_932
		JMP	SHORT LOC_2258
LOC_2262:
		MOV	WORD PTR DS:[0DF80H],DX
		MOV	DATA_170,0FFH
DATA_380	DW	762BH
DATA_381	DW	460AH
DATA_382	DB	89H
		DB	 76H, 06H
LOC_2263:
		MOV	AL,AH
		MOV	AH,0
		POP	BP
		RETF	2
		DB	 00H, 55H, 8BH,0ECH, 8BH, 7EH
		DB	 06H
DATA_383	DW	58BH
		DB	 8AH, 66H, 08H, 8BH, 5DH, 02H
		DB	 8BH, 4DH, 04H, 8BH, 55H, 06H
		DB	 8BH, 75H, 08H,0CDH, 21H, 89H
		DB	 05H, 89H
DATA_384	DW	25DH
DATA_385	DW	4D89H
DATA_386	DW	8904H
DATA_387	DW	655H
		DB	 89H, 75H, 08H, 72H, 02H, 33H
		DB	0C0H
LOC_2265:
		TEST	BYTE PTR DATA_241,0FFH
		JZ	SHORT LOC_2266
		PUSH	AX
		MOV	AH,30H
		INT	21H			; DOS Services  ah=function 30h
						;  get DOS version number ax
		POP	AX
LOC_2266:
		POP	BP
		�`	md	fE8�^	�jEEA�f	�<�b	md	8�f	�E�E�+�a	me	fE8�_	�jEE�g	��c	me	8�g	�E�E�8``xآ��� IՅ �I� �)d ��� �� ������ ��Ս ��� �� ��L�� �� ����dddddL��
������ iܘ
�������� �� �� 8� ��dddd���������Y��Ą������Ƅ �� ă o� � �� � ݈ F� � � �� � ɂ �� ����  <� O� u�� ��2�L����L�� H�LV���������o�	�p�n�u���v w�P H���LV�            Game Over             dddd|�F�	�x�
��������m�s��s����������������������'�������N���O�1�������d�`�1���q���g���h�rI��i� 1g�g�i�01g�g�i�`1g�g�F}x�x� ��0}eg�g���@eh�h���`���Lr��r� g�g�r�0g�g�r�`g�g���1�����` R�)i���@�� R�)�����r R�)���������@ R�F`0 ` � � 0� @�� )�`���y�\�z�L�Z �8�y�~�y�z��zz���`� ����yȭ���y�0ey�y��z� ����yȭ���y�0ey�y��z� ����yȭ���y�0ey�y��z� ����yȭ���y�0ey�y��z� ����yȭ���y�0ey�y��z� ����yȭ���y�0ey�y��z� ����yȭ���y�0ey�y��z� ��yȭÃ�y�0ey�y��z`� �t�7tp�
�	�o�
�p�0 � J)��>��u�?��v�J��<�H�:�z� L������ �ץJH)��M��u�N��vhJ��G�eo�oɠ�do�J�ep�p�����o��A��D�� L��B�΄         @   @	  @@	 @S� ��� @�� `Z�; fZ�fz��`��; @V�  R� @R� `f�; `F�; @   00   DD   FE  VV  ��  ��  ��  ��        00           @   @	  @@	 @S� ��� @�� `Z�; fZ�fz��`��; @V�  R� @R� `f�; `F�; @  ��   ��   ��   ��   00  ��� S�݅7�  �?   ��� 0�������� ��V�� �jUU��ZUU��VT��V @�>�U @�>�  �>�  �>�  �>�U @�>�V @�>�VT��ZUU��jUU���V�� ����� 0��� ���   �?    ��   �  �V�� �kUU��[P��Z@��V  �>�V  ���V  �>�V@��[P��kUU� �V��  �   ��     ��     �j��   ����� �U    U� �����   �k��     ��   �	
	���`�  )�`��̆�g� ��0 φ��g���`�
�������O�
��^�e	��e
�"�1�@��Z ��z�` ��9����Ǣ�� ����`��o�"�p���u���v�OjjjjHj)�}1�1h)��	�(}�ɠ�3�^jjjjHj)�}@�@h)��	�(}"�"ɠ��i���L���i�L��� ���� ��0`���΁`�  )�`���`���������e	�����
������`����È�g�Ј�h��dg��h��eg��8���g��8���h���  ����0`ڽ��oɘ�-���pɠ�$� )��g��u�h��v�i��J����H���z ���`���i� ���`k���� ph
llllllll�lP	$$$d��@@� ph
llllllll�l  �@         ��0`���Ί`�  )�`���ɀ����Ɂ������`��������e	���e
���������)

	���
��`���� V����`���%�}�����}����oɠ�C�5�}����-�}����pɠ�+ު���� �����M�H�
��=��u�>��v�i��zL�螌�i�L��ڢ ��)?������(���`}��gɠ��ڊ}�hɠ������h*���g*)�8�������)���}�)��`  ���   � ���  � �   �U�c�q�}���������� pppp��
 ;�&�9n�� �    �V5� � � �n�9�& ;�
�pppp� � ��
l.�� ;     �/W%�/  ; � �l.�
�� �����������(�������������(�0����~	�	�m0`�ɀ��Ɂ���mn�n�mɃ�� %�� ���mnH ~�ɀjɀje	i�o�oh ��ɀjɀje
i�q�pɠ�!�oɠ�� )�����u����v�i���L��i�L�� ������� ����lQl]������ ����kf:��9��9kf:�����s��s`�mɃ�`�  )�`�mɃ��p�g�r�h o�g�q�h��t��`�gɐ��x�h�|���t��s`��t� "����`�R�u���v�x�o�|�p8�|��|���o�t�i���L����zk���dd\7L7"    ��`�����o���p�����)��
L�� R�)L�� ��`�����o���p��.�V�Ȍ�~�茝�`}ujZG1 �Ϲ������������ 1GZju} 1GZju}}ujZG1 �Ϲ������������ ��`�����o���~�p��.�V�����` ��`�����o���p�`dg T�� eg�g��` ��0�����o�.���p�V��g��` ��`�����o���p��.�V�����` ��`�����o���p��.�V�����` ��`�����o���p��.�V�����` ��`�����o�~�p������` ��`�����o���p������` ��`��������.�V�����~�����������������������,��L�� ��`�����o���p��.�V�����~���  �������i����
�윪�����T��L�ע'����`�'���� ӎ��`)?
��䎅u�厅vlu ���㐚�������������������q�j�s�a�O�����+�ܨ�`������yh��o�yl��p�������o�
��X��u�Y��v�e��d�H�`�zL��p�����   �? �����Z�>�UU:�P�kA�k@�kD�kA@�P��UU:�Z�>���� �?  � ��? �� �V��U�o�o�o�o��U��V��� ��?  �  � ����>�U:oU�kA�kA�oU��U:��>�� � ��:k���k�:�����)�����u����v� �~�
}.�.�}����oɛ�� ���
}V�V�}��pɛ������o�o�^	�p�_	��b	�c	�	�`	�
�a	��d	��e	��f	�g	  �j��e���L�軐Őϐِ� ���� 0 � �� 0 � �g�� � ���� ��
����u���v�M}V�V� }�ɔ������p�}��� ��ɀjɀj}~��ɔ����oڊi��� ����o�^	�p�_	��b	�c	�	�`	�
�a	��d	��e	��f	�g	  ��`ک ��ܠ <��������	���
����"��F`���`�`mNm�N�����`mNm�N����	���ɂ�`������`�N��N��m�	��mɃ�`�m��m�m`
�.�R�v� � ����:( )+)�+)�+)�+ �(�*,�:�� �  � ���A:�A*�A�A�A�A꨾*�A:�� �  � ���:�e9K��������!��:� �  � ����:�U+{A�{ �{ �{A��U+��:�� � ���o��p�� v��
���  <�Lx���)
����}V�V���}�ɐ����o������J)�� ��u�"��v�i�����L��  d � j��� ���j� d $`��            B�  �  uu@YY @Hm @t	@Y� my � �        �  P 0� @^u�e �����PP@�]� d]0��  @ 0     ���o��p����� )}V�Vɐ�	����	��`�� ��ɀjɀj}.��ɐ�F�� ~�ɀjɀj}V�ɐ�/� J)��+��u�,��v�� v��
���  <�Lx��i���L�����	`/�g� *� �)hp)hLii1 Ye  �� ���b���b Z�  Ye Lii1p)h�)h *�  �
  �:  �� �� `	  �)  � � h+  `	 �� ��  �:  �
 ���o��p�P}V�V� }�ɖ�	����	��`��=�����������������#ڥoHi�o R�)i �� R�)i ��h�o����L:��d}.�.� }����	����8}.�.��}����� v�}���$��
�����u����v�����H���H�i�zhL�螶����	�Ƞ  <�Lx�
��ݕ�ݕU�ݕ�
� �E�Z*��e��i��k�[nh��P�W  �� @� ��$  V	  X  �  �� L	��f�	��	��	�~
T_H��G `� `� �$   �  L	  �� f����	��	T/�	H�~
�_`�`G ��  �   $      �   ��L	�	��	f�	�~
�_��T�G H?� � `$ ` �     ���o��p�� v������	���,� <�Lx�����JJJ)�����ɐ�	����	��`���H���H�
����u���v�i�zhL���9�     @  �� �������+��������  �  h
  P  @   @   � �(�
����+�������  �  h
  P  �  �  ���o��p�� v�}���2����	���^� <� x��o�o�o�o�p�p�p�p�)H ��hi� ��`��	����	��`����JJ)��u�v�i���L���.� U P� $�j �������������V��������v������� �� @U  U P� $�j 	U�	U�YU�	U�	u�Y��iͥ�u������� �� @U ���o��p�� v�}�������	����� <�Lx���ɠ�	����	��`�}��� ��ɀjɀj}~���oɐ����o����JJ)��u��v�i���L���3� ��  �1  �1  �1 ���?ж��m�@۶@�m m�  �v  �-  d  �  �  @  ��  �!  �!  �! ���?P۶жm@m�@۶ �m  mk  �  �  P  �  @ ���o��p�� v�}�������	���  <�Lx��7}V�V� }�ɠ�	����	��`���  R��}�/��)?��&J)�Z�����	������Z}V�V� }�z���u���v�J���H�i��zL���@� * �� `�`�X�������������  ?     ���
��*��*��;�������� � ���o��p�� v�}���2����	���^� <� x��o�o�o�o�p�p�p�p�)H ��hi� ��`��)�#ڥoHi�o�pHi�p�}���) ��h�ph�o��� �ߠ Hh�}.�.�}����U}V�V� }�ɠ�	����	��`����JJ)��2��u�3��v�i���L��:�v���� � ��  �
�*�����1C�T0p0C�T0��1����%0�
��  �
  �
 ��  �
�+��A�"!�"!�%�
!�n����
 ���  �
  �
 �� 0)���Y2�Ƥ2�r�2�Ƥ2c�2��) ��  �  � �� 0�����n�#Ja!�$aR(2�A�2���+0�
��  �  ��`�����o���p��.�V�����`���o��pڽ���̜

�Ϝ� v�}���	����	��`��



}V�V��JJJJ(}�ɠ�	����	��`ڽ�
��Ҝ�u�Ӝ�v����̜�Ϝ�H�i�hL��؜�$��	�#N7�6���p/� �  �=  ��؍=<�u}]�$1Ƈ|��]��?t�=F� }� r� �?  �  �s ���B �Aw�? �)��( x	�6�>G�W�+�T})N/���A}<�?A����/�  W��I�
�lI�A�;Q;;W{�6<.�W��|.�3��� �K��	 ����  ��\  ��+   �   ��`���� R�)�g R�)eg����.�V R�)������ R�)��)?��)i�����`���o��p�� v�}�������	���^� <�Lx���
 �߅gdh
��h�	ɠ���eg�g��eh�h���	�
��eg�g��h�g}.�.�h}��������L�����	�*ک<���oHi�o�pHi�p� ��� ���	 ��h�ph�o��M}V�V� }�ɠ�	����	��`�oɠ�`����)H����u���vhJ�����g���h�i��g�hL���X���̟̟��X�� �
 ��� �W���x
h�j)-�
-d-�-Z�-x
h�	��W����  �
  T @�Z ����g���y�By(�y�h�"Jy�@���W����@�Z  T      T @�Z P�k������)�����!��'����P�k@�Z  T           P � �@.n@�l@.n � � P ��`�����o���p��.�V R�����``�ȅ���d�S����Ȱ! R�)?}��o R�)?8�}�p�x�  <�Lr���������F ��G ��� iܘ
��������L����h���m���� m��������d����m�����m�����m���� m����� ��ɀjɀji(���� ~�ɀjɀji(����o��p�P�( v�� eo�o� ep�p�� v�����}������o��p� J)�����u����v��(�G ��F �譪�"Ϊ� eo�o�ep�p��u���v���F �� )��`��2��� }��o� }�p� ����� ��`�����o���p����`��ˤ         $                 �  0          
 �� �   @ j�  �% �� X  ��h�  �� �� V  �R)��
 �% ��? X ���
��% �% ���> X X�
�j�� �5 �]u: \ FF���F�� ��: V������j � �
; �  $�� ��e$ V�Ɠ>�� Y��  ���% X�Ɠ?�% X��?  ��Ɩ �9��l ���  ��  ���o  �� @j՗� @�����o ��W� �Z�� @��瀾 o�*  ������
����ZR�  �F
�F_�������  ��h��zl9���b)��   �Z�h�N����n)J��    ��V�Kp����P�?    ���vr�󍝎&��     �j`����O�n	��      �k���}}��^$�      P�Z�KqC�M�^��     ��o���O�n�_j    ��ڿ�:�s�c�����    	������а�_��`    d��j��ʣ�����    �����~���:����>    ����o��+����    h�_��#��V/ȫ��)    ��忺 l��9 ��[�z    ��?����k��
�>��    ����/\��W�5�N�_     Z��+������Ϫ�      ����޾����ë�      �� \�[�N5� �:      � �
��
  �            `	                 ��        `      ��      	�
 �   ��    �@�
 �  �@>  � �d�j� �	  �@�  ` ��j�
�%  �@�  X�
� ��%�%  k���  XXZ�  ����5  �T�  \F��  �F�  ;$�  �����  �j� o�
� �& $�>  ��e$`
 o�C� �	Y�  ���%����C�0nX��  īƖ &9��K>l� ���  X�� 89�&�>l, ��%  �՗� |9�ڧl= ��W
  ���� @��ڧ�� or�
  ������
����Z��  ��F
�F[少����  ��h��zl9���b)��  ��j�h�N����n)J��   ��V�Kp�������    ����vr�󍝎&��?    ��j`����O�n	��     �k��nsι�^$�      P�Z���@�^��     ��o��nC¹�n�_j    ��ڿ���pO�����     ����������_��     	��j��ʣ�����?`    �����~���:����    �����o��+�����?    �_��#��V/ȫ���    ����� l��9 �~Z_     Z�����k��
����      ��/\��W�5�Ϋ�      ���+�������:      ���޾�����         \�[�N5�            �
��
                `	         qC�O¹�sO�N�F�S�\V�5�*���(UU(�Ԣ��C�*��I��aT���P P ��
��Ȩ}.�.�ɨ}����oɐ�4�Ҩ}V�V�Ө}��pɐ��� v����u���v�i���L�螶�i�L�� �? �W�p�j���6��6�@��  ��  ��  ��  ��@ۜ�6���6p�j�W� �? ,���  s � � ,� �ȅ���<�  � H�`����Ȱ  R�)?�}��o R�)?}�p�� <�Lr���������'��ɀ����� ��� iܘ
��������L������� ��}!� �߼� �ۘ����}!�
 �߼� �ۘɀjɀj}�����
�Ȣ ک�u���v��i}��o���p����� �����	�֥ JJJ�ˠ���[���u�v��}�i�o���p�g�E8�g��
�( ��(�( v�� )?��`)�` ��`�����eo���ep�`"*17<@CE 	$-6?HQ   �    �     ���  ʛ    ����ڛ    �۩�j��   ��۩�j��  �曧:�ڛ�  �&�z��  �曧��ڛ�  �v��Z��  ��E\��u��   �Z���V��   ����Z����   �ڪ�VU���   �ۺ�UA���    o�U��z>    ���V���:   ��������   𪫫���z�  ��j���l��  \�J�[�X�  ��R�o�\��; ��T�[���� ���ÿ�����j��[��Z�������o��������>���:��  ��꿪����  ﾖ������> ���Z�i�o��� ��o���o>�� �����Z�����  ���V����>  ����V����  hj�j�U�^j*  ZY�V%V�~Y9  ��oU	XU��) ���^���F�� ���^X	P��� ���n�X�_��� ��ﺿ����� �j뺭�j��z� �k�������{�  j�������{*  k����i��{:  ���������  ���jUU���  ���VUU���   @��UUU��{    ��UUU��;    �UUA��    ��U ��    ��V  ��     �V @�+      �ZP�       �U�*        ���                             $        F�       ��      �Z��     ��k�    �����    ����    ����*    �+�z�n    �)n�hj   �����rn? �k��_R��0�v~��n��߻�z�!JC���my����̊>l9��3��7 � ����Y `	 e���V� X% ���̪� h) j�3��� �� ����:[���N��>l9�������.������Z����k��V���k��Z���k��j����  ����>  �:� k�  ��  �0  P:  ��  ��:  ����Z�  �^�
��   LUTU1     @T               $        �       ��      �Z��     ��k�    �����    ���j    ����*    �+�z�n    �)n�hj   �����rn? �k��_R��0�v~��n��߻�z�!JC���my����̊>l9��3��7 � ����Y `	 e���V� X% ���̪� h) ��3����&������[%�N���>l9��B:k������k�V����>�k�U�  kU>�k��:  ��>鬽�  ��~:���  ��O:���    �C:�    0��      ��*      � k      �  �=    |�  |�    �=  \�    j5  �  �Z  @U
  �U   T  P   �* �V�`�	��'ب*'6���6���6���6���6���6���ب*'��'`�	�V� �*  ����V���� hj�j�U�^j ZY�V%V�~Y ��oU	XU�����_���F�����_X	P�����o�X�_�������������j��������k������ j������� k����i�� ��������� ��������� ��������� @�������  �������?  �������  ���ZU��  ���UU��   ��U��?    �V��     ���?      ���   ���o��p�}�ɠ��� v��V�u���v�i���L�螶����	`<;;�999999999999<� �b	�c	�o�^	�p�_	� �� ����g`�	�`	�
�a	��d	��e	��f	��g	  �j�`��f	�g	dg α �� 2�Lh���d	�e	����`	�"�a	  ��
�g���o	���`��d	��e	��f	�g	�mɃ�� �� �o�`	�q�a	  ���g`��d	��e	��f	��g	�  M����0`���`	���a	  ��`�g`��d	�e	��f	�g	������`	���a	  ��
�g����	����`�`�  )��
�
�
����
�  )��
�
�
Ɉ����
�  )�
�	�	���	�  )��	�	�	ɐ����	`� )�`��o� �p�5�u���v w��=��>��?� �@ m�H ��G ��F ��EL��SCORE: e��e�����`�  )�� H�  )��� H�  )��� H�  )���`�s�8�����`���`��������`� �������������`e���ȱ
�ȱ�oȱ�p�e����߳�u�೅vlu /�E�t���!�����h�*������`��dX,WORD PTR DS:[2]
		ADD	AX,WORD PTR DS:[4]
		ADD	AX,WORD PTR DS:[6]
		ADD	AX,WORD PTR DS:[8]
		ADD	AX,WORD PTR DS:[0AH]
		ADD	AX,WORD PTR DS:[0CH]
		ADD	AX,WORD PTR DS:[0EH]
		INC	BX
		LOOP	LOCLOOP_2310

		MOV	CX,ES:DATA_5E
		SUB	CX,ES:DATA_4E
		MOV	BX,ES:DATA_4E

LOCLOOP_2311:
		MOV	DS,BX
		ADD	AX,WORD PTR DS:[0]
		ADD	AX,WORD PTR DS:[2]
		ADD	AX,WORD PTR DS:[4]
		ADD	AX,WORD PTR DS:[6]
		ADD	AX,WORD PTR DS:[8]
		ADD	AX,WORD PTR DS:[0AH]
		ADD	AX,WORD PTR DS:[0CH]
		ADD	AX,WORD PTR DS:[0EH]
		INC	BX
		LOOP	LOCLOOP_2311

		SUB	AX,CS:DATA_55
		SUB	AX,WORD PTR CS:[3B2H]
		MOV	BX,ES
		MOV	DS,BX
		MOV	CX,0FFF8H
		SUB	CX,SP
		SHR	CX,1
		MOV	SI,SP
		ADD	SI,6

LOCLOOP_2312:
		ADD	AX,[SI]
		ADD	SI,2
		LOOP	LOCLOOP_2312

		SUB	AX,DS:DATA_7E
		MOV	CX,DS:DATA_3E
		SUB	CX,DS:DATA_2E
		SHR	CX,1
		MOV	SI,DS:DATA_2E

LOCLOOP_2313:
		ADD	AX,[SI]
		ADD	SI,2
		LOOP	LOCLOOP_2313

		RETN
SUB_938		ENDP

		DB	7 DUP (0)
		DB	 01H, 02H, 03H, 04H, 05H, 06H
		DB	 07H, 08H, 01H, 02H, 03H, 04H
		DB	 05H, 06H, 07H, 08H, 01H, 02H
		DB	 03H, 04H, 05H, 06H, 07H, 08H
		DB	 01H, 02H, 03H, 04H, 05H, 06H
		DB	 07H, 08H, 01H, 02H, 03H, 04H
		DB	 05H, 06H, 07H, 08H, 01H, 02H
		DB	 03H, 04H, 05H, 06H, 07H, 08H
		DB	 01H, 02H, 03H, 04H, 05H, 06H
		DB	 07H, 08H, 01H, 02H, 03H, 04H
		DB	 05H, 06H, 07H, 08H, 00H, 00H
		DB	 05H, 00H, 29H, 45H, 3CH, 2DH
		DB	 2DH, 00H, 00H, 00H, 07H, 00H
		DB	29H
		DB	'E     Personally Developed Softw'
		DB	'are  '
		DB	 19H, 00H
		DB	')EFor IBM Personal Computers  '
		DB	 17H, 00H
		DB	 29H, 45H, 2AH, 2AH, 2AH, 2AH
LOC_2314:
		ADC	AL,[BX+SI]
		SUB	[DI+2AH],AX
		SUB	AH,[BX+SI]
		AND	[BP+SI],DL
		ADD	[BX+DI],CH
		INC	BP
		AND	[BP+SI],CH
DATA_395	DW	202AH			; Data table (indexed access)
		DB	20H
DATA_396	DW	420H			; Data table (indexed access)
DATA_398	DW	2900H			; Data table (indexed access)
		DB	'EPersonal Editor II  '
		DB	 05H, 00H, 29H, 45H, 2AH, 2AH
		DB	 20H, 20H, 12H, 00H
		DB	')E *****'
		DB	 12H, 00H, 29H, 45H, 2AH, 20H
		DB	 20H, 20H, 14H, 00H
		DB	')E (C) Copyright IB'
LOC_2315:
		DEC	BP
		AND	[BP+DI+6FH],AL
		JC	SHORT LOC_2322
		AND	CS:[BX+DI],DH
		CMP	[BX+SI],DI
		XOR	CH,[SI]
		XOR	[BX+DI],DI
		CMP	[DI],DH
		AND	[BX+SI],AH
		SBB	[BX+SI],AX
		SUB	[DI+20H],AX
		PUSH	DI
		JC	SHORT LOC_2323
		JZ	SHORT LOC_2324
		OUTS	DX,BYTE PTR GS:[SI]
		AND	[BP+SI+79H],AH
		AND	[BP+SI+69H],CL
		INSW
		AND	[BX+79H],DL
		INSB
		INSB
		IMUL	SP,WORD PTR [DI+20H],520H
		ADD	[BX+DI],CH
		INC	BP
		INC	SP
LOC_2319:
		DB	'o you really want to quit? Type '
		DB	'y or nBlock mar'
LOC_2320:
		IMUL	SP,WORD PTR [BX+SI],72H
		DB	'equiredColo'
LOC_2321:
		JC	SHORT LOC_2325
		IMUL	SI,WORD PTR FS:[BP+DI+70H],616CH
		JNS	SHORT LOC_2326
		OUTSB
		OUTSW
		JZ	SHORT LOC_2327
		IMUL	BP,WORD PTR [BP+73H],6174H
LOC_2323:
		INSB
		INSB
		DB	'edUnknown c'
LOC_2324:
		OUTSW
		INSW
LOC_2325:
		INSW
		POPA
		OUTSB
		DB	 64H, 43H, 61H, 6EH, 6EH
LOC_2326:
		OUTSW
		JZ	SHORT LOC_2328
		OUTSB
LOC_2327:
		POPA
		INSW
���� ��ɀjɀji<�����o����p�0�( v��+�u���v��8�G ���}��o�i0�p� � v��}����������	���`Ϊ����o�i �p�+�u���v�
��FL�襇H)�&  �� �h�& `��H)�&   �h�& `      (  <  �  x  d  P       (  <  �  x  d d P  ( P x ( P x ( P x ( P x ( P x ( P x ( P x ( P x ( P x ( P x  < d	 �  < d	 �  < d	 �  < d	 �  < d	 �  < d	 �  < d	 �  < dd �( xx xP xP xP xP ( xx xP xP xP xP 
 F 2� ( P 2x 
 F 2� ( P �x 
 F 2� ( P 2x 
 F 2� ( P �x  (<Pdx� (<Pdx� (<Pdx�(F  > (N  6  F (V  .  >  N (^  &  6  F  V (f    .  >  N  ^ (n    &  6  F  V  f �v (F  > (N  6  F (V  .  >  N (^  &  6  F  V (f    .  >  N  ^ (n    &  6  F  V  f �v (F  > (N  6  F (V  .  >  N (^  &  6  F  V (f    .  >  N  ^ (n    &  6  F  V  f �v P 
  2 F Z n � �� �P      �2��d�d(�d<�dP�dd�dx�d��
P 
P 
P 
P 
P 
P 
P ( �(��   " 3 D U f w ( �(��
( 
( 
( 
( 
( 
( 
( ( �(��
x 
x 
x 
x 
x 
x 
x ( �(��  
   ( 2 < F P Z d n x � �   
   ( 2 < F P Z d n x � �   #�   #�   #�   #�   #�   #�   #�   #�    ( < P d x �P   
   ( 2 < F P Z d n x � � 
  

 
 
 
( 
2 
< 
F 
P 
Z 
d 
n 
x 
� 
�   
   ( 2 < F P Z d n x � � d  d d, dB dX dn d�  P      - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x �     - < K Z i x � -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix�
 


-
<
K
Z
i
x
� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix�< <<<-<<<K<Z<i<x<��	 �	�	�	-�	<�	K�	Z�	i�	x�	�d	 d	d	d	-d	<d	Kd	Zd	id	xd	�<	 <	<	<	-<	<<	K<	Z<	i<	x<	�	 			-	<	K	Z	i	x	�d ddd-d<dKdZdidxd�d ddd-d<dKdZdidxd�d ddd-d<dKdZdidxd�2 222-2<2K2Z2i2x2�2 222-2<2K2Z2i2x2�2 222-2<2K2Z2i2x2�2 222-2<2K2Z2i2x2�2 222-2<2K2Z2i2x2� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix� -<KZix�
 


-
<
K
Z
i
x
�
 


-
<
K
Z
i
x
�
 


-
<
K
Z
i
x
�
 


-
<
K
Z
i
x
�
 


-
<
K
Z
i
x
�
 


-
<
K
Z
i
x
�
 


-
<
K
Z
i
x
�
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  �Hژ��,
�h� h�`�;�<� �;H
��0׍\	�1׍]	� -����`l\	6�D�Rע �;� �����`� �;� �����`� �;�( ��������;`� ��	� ���)�� ���:	� ����"�� � � �( ����`d �ע!�:	�����(�	���` �ץ��`�(t���!����L�ל��'�(� � �'���������,� �)������/�0�1�`��`�/��L����0��0�`� �/�1m��0�,�
�)�	�)�� L�ٽtڪ��%� �&�/� �%0L�����L�����L������ �,����� |ڱ%�1m��0 |�LC���� |ڱ%�	�%8�	�%�&� �&LC����L�����������}xڨ���%���& |�LC����- |ڱ%H |ڱ%H��}xڨ�%���&������h�&h�%LC����' |ڤ/�pڠ �%�	������%i�%� e&�&�/LC���� |ڱ%Hȱ%�&h�%LC����2�pڹ	)��	:�	� �	� ��%��1ۦ/�)L�� |� |�LC�����/�p�)��	)�	�	�	 |ڦ/LC�ɀ�(逼p�

��:ۙ	�;ۙ	�<ۙ	�=ۙ	 |ڦ/LCؤ/����pڨ��ڝ ��ڝ �	� �	�  |ڠ �%��1ۦ/�) |ڥ/
��%��&� �/��������`�.��+��+�L�٠ �#���� �.L���� �ڱ#�	�#8�	�#�$� �$L�

� �ڱ#��1ۅ+ �ڽۍ( �ۍ) ��)�* 	�* L��   �%��&`�#��$`H���	
�	hJH��m	�	hn	n	��	�	`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   �=�>� 8�=H� �>�h`H�=E=�=�I�i�hI�i ��$=� 8�EH� �F�h`H���E
�FhJH��eF�FhfFfE��E�F`�>EBH$>� 8�=�=� �>�>$B� 8�A�A� �B�B �h� 8�E�E� �F�F� �G�G� �H�H`� �H�G�E���FF>f=��GeA�G�HeB�HfHfGfFfE��`�=�>E>�>I�i��=I�i i�(I�i`�=�>� �H=�*�>��>�h*��`�>EAH�AI�i�A$>� 8�=�=� �>�> ��h� 8�E�E� �F�F`��EJ�F�?=&>&?�?8�A��?&E&F��`�@EBH$B� 8�A�A� �B�B$@� 8�=�=� �>�>� �?�?� �@�@ )�h� 8�E�E� �F�F� �G�G� �H�H`��EJ�F�G�H�C�D=&>&?&@&C&D�C8�A��D�B��C�D&E&F&G&H��`���lݐ��lݘ` 	$1@Qdy����=�>��A��B�F�E�=&>&E&F=&>&E&F8�E�A��F�B��F�E��**EA*�A&B���FBjFBj`��8��
��i
�=�



=`�=�>��=��ݥ>� ސ
�>�=��݅=8&E&F���E�F`    
  ( P d � � ���@�E�=�Oޥ>�Pޥ?�Qސ�?�=�Oޅ=�>�Pޅ>8&E&F&G����`        
    (  P  d  �  �   � � � @ '  N @� �8��@� 5�I �߅A�I ~߅B�N�A �ۅg�h�MH�B ��8�g�g��hg*�M�N�B �ۅg�hh�A ��eg�g�ehg*�N`�J �߅A�J ~߅B�L�A �ۅg�h�NH�B ��8�g�g��hg*�N�L�B �ۅg�hh�A ��eg�g�ehg*�L`�K �߅A�K ~߅B�M�A �ۅg�h�LH�B ��8�g�g��hg*�L�M�B �ۅg�hh�A ��eg�g�ehg*�M`I�8i@�@�$���%

JJ(�I�i )?����(�I�i ��`� `�� `����` 	"%(+.0369<?ADGILNQSUXZ\^`bdfhjlmoprsuvwxyz{||}~~8�S�O�W�T�P�X8�U�Q�Y�V�R�Z� �[�\�]�^�\�h�[FhjFhjFhjeO�S�\)�heP�T�^�h�]FhjFhjFhjeQ�U�^)�heR�VL��\�h�[FhjFhjFhjFhjeO�S�\)�heP�T�^�h�]FhjFhjFhjFhjeQ�U�^)�heR�V�We[�[�Xe\�\�Ye]�]�Ze^�^`�)�A�JJJJ�B�i)


8�A�=�i)�J8�B�>�j)


�?�j)�J�@�ge=fE8�o�jEE.�=e?8�A�E�E� �he>fE8�p�jEE�>e@8�B�E�E�8``H�ZE����e����充��  E��� �� O��s��tz�h@���+� ��� ������m���͖�� � � � ��`
��
m��� ��ᙑ������`�,
� � 8� � 
�@@ 
��<� ( �   �S����P�  ���� ��z�@�X�����>l���?�  �����  � � � � � � � � � � � �Ʌ��& ���d��O���n	���^�N��OL�ש �u�@�v�����_�'�u���0eu�u� ev�v���` U���p


 w�o
ey�y��z`����y�#�z` 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]H� ��hHJJJJ ��h)	0�:���H�Z�uZ�vZ ��z�vz�uz�h`8� dv
&v
&v
&vi��u��ev�v� Z�u�i @��y @� �y�0ey�y� ez�zz����8�y�~�y�z��z`���s�g���s�hFi�	Fh*Fh*La�Fg*Fg*Fi�	Fh*Fh*Lt�Fg*Fg*Fi�	Fh*Fh*L��Fg*Fg*Fi�	Fh*Fh*L��Fg*Fg*`        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d�  �U�L|��p c� �u�����u��v������� ��L�`dodp� Z�{ ��z���Z�|�{�| ��z�����`H c��o�oI��o�phdvi��v
&v
&v
&v
&ve{�u�|ev�v� �u� �y��u��y��u�0�y��u�1�y��u�`�y��u�a�y��u���y��u���y��u���y�	�u���y�
�u��y��u��y�z��u� �y��u�!�y��u�P�y��u�Q�y�z`�{�u�|�v� dg�C�h��� �u�g��(���'eu�u��v�0eg�g��h���`�
��^
�o�n	�p��	�u��
�v��
`�g�h c� �u�y��g���eu�u��v�0ey�y��z�h��`�O ����`���n	`� �P�p�P�p�P�p�P�P�P���P�p�P�� �� n� q� �PI�=p�p�PI�=p�p�PI�=p�p��ܽPI�=p�p�� ��L��lN�O�n	��� ����`�
���^
����
�u��
�v��	 w�n	JJey�y��z�n	)
���ꅌ��ꅍ��	d�
&�
&�}�	�����Pe����e����n	JJHJJJe����扼
�n	)�ȹ�ꅎ��ꅏ��ꅐd�h)���&�&�&����iv����� i녗��� e�����ڥ��������������� �� �����ȥ����ȥ����ȥ������eu�u��v�0ey�y��z�e�����ƋЫ�` ?�����������������         ?���������                 ?������@�l� � �u g��Ċ��`� dk�kdk)�l�u
&k
&kl g��Ċ��k) g�`� dk�kdk)�l�u
&k
&k
&k
&kl g��Ċ��k) g�`� dk�kdk)?�l�ujj�kj)�l g��Ċ��k)? g�`��y`�����5���`�����߿�����߿�����߿�����߿        �p�k��l� �u�@�v�{�w�|�x�L���  �� �� �� �� ���0eu�u��v�ek�k��l��΢�� �k� c��k�� c��k�� c��k�� c��k��  c��0eu�u��v�(ew�w��x�ek�k��l�Ч`�gFg��w�u�Fg��w�u�Fg��w�u�Fg��w�u�Fg��w�u�Fg��w�u�Fg��w�u�Fg��w�u`�k��H�


�hL�� �k� ��k�� ��k�� ��k�� ��k��  ��0eu�u��v�ek�k��l�в`�g� Fg��u�Fg��u�Fg��u�Fg��u�Fg��u�Fg��u�Fg��u�Fg��u` K�s�s��`�sEtM  e�*��E���e���&�E���`�|�=٬�>���?���@����@�=���=�>���>�?���?8&E&F&G&H�����`            
      (   P   d   �   �     �  �  �  @  '   N  @�  �8 �� @ �  5 @B ��  	=  z ���  -1 Zb ��2�������  60  0  0  0  0  0  0  0  0  0  0  0  0 & 0 & 0 & 0 & 0 
 0 
 0 
 0 
 0 	 0 	 0 	 0 	 0  0  0  0  0 $ 0 $ 0 $ 0 $ 0  0  0  0  0 % 0 % 0 % 0 % ��  #0�9������	���  :	!	 ���  50�����������  6 0 0 0 0 0  0  0  0  0 0 0 0 0 00 0  0  0  0 0 0 0 0  0  0  0 000 0  0  0  0  0  0  0  0  0  0 000��  #0������������  :
) ' )  ,���  '0�����q�����  :�����0000&(0(00(0&(00   & 000&&0��  %#0#000#0#00000#00#0#000#0#000#0#000	0	000#00#00�q�     ��������  60  0 ' 0  0 ' 0  0 ' 0  0 ' 0  0  0  0  0  0  0  0  0  0 ' 0  0 ' 0  0 ' 0  0 ' 0  0  0  0  0  0  0  0 * 0  0 ) 0  0 ) 0  0 ( 0  0 ( ��  #0�����I�S���  60 0 0 0 00 0 0 0 0 0 0 0 00 0  0  0  0  0 0 0 00 0  0  0  0 0��  #0����Z�������  6 0  0  0  0   0   0  0  0  0  0  0  0   0   0  0  0  0  0  0  0   0   0  0  0  0  0 ! 0 ! 0  0  0  0  0   0   0  0  0 ��  #0�a���������  60 0  0  0  0  0  0  0 000 0  0  0  0 # 0 # 0  0  0 000 0  0  0  0 0 0  0  0 ( 0  0  0 0 0  0  0  0  0  0 0 0  0 0000��  #0�
��0  0   0   0  0  0  0  0 ! 0 ! 0  0  PTR FS:[SI]
		JA	SHORT $+70H
		POP	BP
		POP	BX
LOC_2515:
		DB	'fn][mb][el][we][mb][u'
LOC_2516:
		JO	SHORT $+5FH
		POP	BX
		DB	'el][we][right][cm'

SEG_A		ENDS



;------------------------------------------------------  STACK_SEG_B   ----

STACK_SEG_B	SEGMENT	WORD STACK 'STACK'

		DB	256 DUP (1)
		DB	 02H, 01H,0B9H, 10H, 00H, 00H
		DB	 1AH, 0FH,0FEH, 02H, 00H, 00H
		DB	 00H, 00H, 00H, 00H, 8CH,0C3H
		DB	 8BH

STACK_SEG_B	ENDS



		END	START

		POP	BP
		POP	BX
		OUTS	DX,WORD                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                
                  �����������������������������������������
                          SOURCER DEFINITION FILE
                  �����������������������������������������

 ������������������ Section 1: CONTROL INFORMATION   ������������������

Analysis Options = a b c d e f g h i j k l m n o p q r s t u v w x y z
uP               = 386
File format      = ASM
Word style UPPER
Label type       = Decimal
Remarks          = Interrupt & I/O only
Segment display  = Name
Target Assembler = TASM-3.0
Input filename   = PE.EXE
Code style       = Exe
Drive (output)   = C
Output filename  = PE.ASM
Passes           = 2
Xref             = OFF



 ������������������ Section 2: RANGE DEFINITION      ������������������

 ���� Segments ��������������������������

  begin      end      default	   seg	 seg          seg
 seg:off     off     ds     es	   type	 size         value
 -------     ----    ----   ----   ----- -----        -----
SEG_A:0000   FEFF    SEG_A  SEG_A  AUTO	 USE16       ; 8E2E
SEG_B:0000   0112    0000   0000   STACK USE16       ; 9FCE

 ������������������ Section 3: REFERENCE DEFINITIONS ������������������

 ���� Subroutines �����������������������
  seg:off    type & options	labels & comments
  -------    --------------	----------------------------------------------
0000:0001    SUB, FAR			       ; SUB_1
0000:0003    SUB, FAR			       ; SUB_2
0000:0005    SUB, FAR			       ; SUB_3
0000:0007    SUB, FAR			       ; SUB_4
0000:000D    SUB, FAR			       ; SUB_5
0000:002B����  :�����0000&(0(00(0&(00   & 000&&0��  %#0#000#0#00000#00#0#000#0#000#0#000	0	000#00#00�q�     ��������  60  0 ' 0  0 ' 0  0 ' 0  0 ' 0  0  0  0  0  0  0  0  0  0 ' 0  0 ' 0  0 ' 0  0 ' 0  0  0  0  0  0  0  0 * 0  0 ) 0  0 ) 0  0 ( 0  0 ( ��  #0�����I�S���  60 0 0 0 00 0 0�ɍ& LV�'�����