����|�<�����|�<�����<�|�����<�|�����<�|�����<�|���������4�P�l���؇8����؈�؉X����X�j���(�h����R�����(�8�H�X�h�x���������Ȍ؊،�����(�8�H�X�����������������"�2�B�R�b�r�����������TUU���z���oyUUmy��my֖myV�my^�myz�my֕my��my��myUUm���o���zTUU���?���߯�����������j������������o������������������������?     ��  �� �U � � _U �U�� ���_���_��  ��p?�pp�� ��  �� �U � � _U �U ��  �_  � � �  �?  0?  \  ��      ��  �� �U � � _U� �U� ��� �� �?  �? �?� �< \ ��  �� ���U �� _U �U� �Ր ��� �� �  �  �?  <    <?      �/ ��� �U� �W� pW� @U� �U7  W������? �?��� �?�P@�� �/ ��� �U� �W� pW� @U� �U�  W  �? @�? @�?  �  �  �  5  ?      �/ ��� �U� �W� pW� BU� �U� ��? ��?  ��  ��  �� <� �@5 ?� �/ ���0�U���W� pW��@U� �U� W ��? ��?  �?  �  �3  �<  P�  �<          �?  ��  |� _U_U�\U�_U�� � _�����?�                �  � �W= �U� �U��U5�U��W���� W� �����  �     (�(P  ����?�_��W��W��W� W�  _�  � �W������ �      (�(P  ����?�_��W��W��W� W�  _�  � �_���� �  �           �?���� _� ����_U�\U_U _U |� ��  �?               � �����W� ��� �W��U��U5�U��U� �W=  �  �             �  �� ����W� �  _�  W� �W��W��W��_���?��P  (�(      � �����_� �  _�  W� �W��W��W��_���?��P  (�(              "       ��� ��"�u� |U |U @U  �� ����4���
��7       "       "        �? ��  ~� _]  WU  W  �� ����4���
��7�0�?�����w�?|w�=������� ��  �?  �?  ��  ?� ��P��  ?UUUU�������������j��������������UUUU�j���j���ik��j���ik��j���o�� � �?  3��� �*�3�
� ��� �0 �?� ��? �?| �?P ��  ?� @p�� � 0�?  � �0�����0�� ��3 �?� �� �? �? ��  ?� @p�� �  �?  �� �W�@w�  �  ��  0 �������?�� ?� ��P��  ?�  �" " �  �      �
�"  �      �* �"   "      ����� � ������?���� ��� �?� �� �0� ��� ����� �����"   ��
 @U  �� �� 9 @ �  �  �  �  �  �  �  �  �  � � 	�@ l� ��  �? @U T T��)�)���~�~�������PU� � ��>  > ��>  > > >  > > >  > ~U>  > ��>  > ��>  >  P T@A� ����@�o��o������V���� ��W��  ��:�  ����  ��P�  ��W��  � ���  � ��                              �  �                             ���?���?�����  �  �  ���?���?  �?  �?  �?��?��?���������?���? �  �  �  �  �  �  �  �  �  �  �          ��������?��?��?��?��?��?��?���?���?��?��?��?� �� ���������?��?�  �  �  �  ��?��?��?��?��?��?���������?���?�  �  �  �  �  �������  �  �  �  �  ���?���?�  �  �  �  �  �  �  �  �  �  �  �  �  �  ���?���?��������?��?�  �  �  �  �  �  �  �  ��?��?���������?����?  �? �?��?��?��?��?��?��?��?��?�?�?  ��������?  ? � ?     <  ?<� �<�??<�<��                                    �������?���?���?���?���?���?���?���?���?���?���?��?< �< ����?���?��?��?��?��?��?��?��?��?��?��?��?��?������������?��?��?��?��?��?��?������ ��  ��  ��  �  � ��������?��?��?��?��?��?�������? �? �?<�?<< �< ��<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�        �?          � ����<0< � <<�  �?< < �< < �?  < < < < < < �?  �<0< < < <0�  �?������  �<<<<�<<<0  �0<<<<�?<<<<  �����������������������������������������������Վ����? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                           0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____8xHxXxhxxx0$)@$+P$.`$'P</`<0p<'�<1,"*<"'L"0\"'l"*0H8H@HHHPH`HhHpHxH�H�H(d 0d@d HdXd `dpd xd�d �d(| 0|@| H|X| `|p| x|	�|�| HAPAXA`AhApAxAHWPWXW`WhWpW@A�  � 
� � � � F�В?���;�є@�ĕB�󖘗(���9�ək����*�؜h��O�������L�ʡQ��J�ԣX�����ŦR�觫����y�'���;�ˬU�� 0@P` `p�� (@( `(�( 8�8 H0H@HPH`H �H XpX�X#�X h@h Phph�h#�h xpx�x#�x �0�@�P�`�p������8�8�  0 @ P ` p �  000#@0#P0`0�0�0 @0@#@@ `@ p@ �@ P0PPP �P `0`#``p`�`�` p0p@pPp`pp0p0�HXhxH x 0(080H0X0 x0�0�0@8@ X@#h@#x@ �@PXPhP#�P`(`8`H`x`�`�`HpxpH�X�h�x��@�@� 0@P`p��( (0(#@(#P(�(808#@8#P8p8 �8�8HPH �H �HX X0X @XPX`X�X h�h�h�h x0x@xPx`xpx�x0H0H�  0 @  0#@  0 #@ P ` p � �  000#`0 �0�0 @0@#@@ P@ �@ P0P#PP`P �P `@`P`p`�`�` p`p �p �0�@���@�P�`�p����������(8HXhx�((8(X(#�((8H8 h8 �8(H8H#XHxH#�H(XHX hX �X(hXh#xh�h(x8xHxXxhxxx�x8h8h� 0@P (P(`(p(�(�(�(8 8@8 `8 �8#�8#�8HPH pH �H#�H#�HX X@XPX`X �X#�X�X hph�h�h x0x@xPx`xpx H H�(8HX((X(h(x(�(�(8(888#H8#X8#x8 �8H8H#HH#XH#hH �HX8X HX XX hX xX�X�Xhxhx(x8xHxXxhxxx�H�H�(8HXhx�� � 0�0(0 80 H0 X0 h0 x0 �0 @X@�@(@#8@#H@#h@#x@#�@#P�P(P#8P#HP#XP#hP#xP#�P#`�`(` 8` H` h` x` �` p�p�(�8�H�X�h�x�����X X �(8HXhxx((x(((8(H(X(h88x8(#88#8H#8X#8h#HHxH(H8HHHXHhXXxhhxxxxx( x8 xH xX xh ��x��h�x��(�8�H�X�h�xHH�(8HXXhx��(8( H( X(h(�(888 �8H(H8HHHXH�H8XHXxX�X�X8hHhXh�h8x�xHx#Xx#hx#8�H�X�h�x���((�P`p�0 @ P � 00`0 �0�0 @0@P@p@�@�@ PPPpP�P#�P `@`p` �`#�` p@p �p#�p �0�@�P�`�p�����p p �(8HXhx��(X( x(#�(888 X8 h8#x8 �8H(H#8HHH#XHhH#xH�H#�HX8X HX#XX xX �Xh8h#Xh �hx(x8xHxXxhxxx�x�x�h�h�@P`p�   0 @ � � � 0@0 `0 �0@@@ �@ �@P P0P@PPP`P pP �P�P�P0`@`#P`#�`0p@p#Pp#`p#pp#�p0�@�P�`�p��� 0 0� 0@@P`p���(`(�(808 `8 �8H H@HPH `HpH�H�HX X#0X@X`X �Xh h#0h#@h#Ph �h�hx0x#@x�x� �0�@�P�`�p���  �0@P`p   0 p � � � 0P0�0@0@ @@p@ �@ �@P0P PP `PpP �P` `0`@` P`#``#p`#�`�`�`0pPp#`p#pp#�p#�p0�@�P�`�p�����P P �(8HXXhx��(8(H(#X(#x( �(888 H8#X8#h8�8H8H HH#XH#hH�H�HXHXXX xX �Xhhh �hx(x8xHxXx�xX�h�x������x�x�(8HXhx�� X h #� 0(0#80H0 h0 �0@8@X@h@x@ �@PXP�P`(`X`x`�`(p8pXp#�p�p8�H�X�h�x���( ( �0@P`0@#`p���( (0(@( `(p(�(�(#�(8@8#P8 `8#�8HPH`HpH �H �HX0X @X PX#`X�Xh@h Ph#`hph�h�h�hx x0xpx#�x0�@�P�`�p����X�X�(8HXhx��(H(X(#h(#�(�(888 H8#h8 x8�8HHH hH �HX8XHX hX#xX �Xh(hHh#Xh#hh�hx(x8xHxXxhxxx�x�xXHXH�(8HXhx��(�(888 H8#X8#�8�8H(H8HHH#XH#hH�H8XHXXX hX xX �X8h�h8xHxXxhxxx�x�x�(�(� 0@P`p (p(�(�( 808P8#`8 �8 H@H#PH `H#�H X@X PXpX�X�X h0hph0x@xPx`xpx0(0(� ( 8 H X (#Xhx�� 8 X h � 080 x0 �0@(@ 8@X@�@�@P8PHP XPhP�P�P`8` h` x`#�`#�`pXpxp�p#�p�X�x�#��#���(�8�H�X�h�x������0�0�(8HXhx� H X #h x #� � 080 H0#X0 h0#�0#�0@X@#h@x@ �@�@P(P8PHP�PH`X` h` x` �`Hp�pH�X�h�x���hphp�(8HXh h 080 h0x0�0�0@8@ H@X@#h@#x@�@P8PHP#XP#hPxP �P`(`8`H`x` �`Hp�pH�X�h�x�����(P(P�(8HXh ( X #h x � � 0H0#X0 h0#x0 �0@8@ H@h@x@ �@PHP#hP#xP �P`8` H`X` h`x`�`�`pHp#hp#xp�(�8�H�X�h�x��0�0�8 H X h 8H#X#h8 H #X #h x � � 0(080H0#X0#�0@H@ h@ x@ �@P8PHPXP �P`H` h`�`p8p hp�p�p�H����(�8�H�X�h�x���8�8��(8HXhx�( � (0H0 X0 h0 �0(@8@H@#X@#h@#x@�@(PHP#XPhP#�P(`H` h` �`(pXp�p(�8�H�X�h�x���8080�(8HXhx��(((#8(#H(#�(8(8#88H8#X8h8 x8�8H8H HH xH �HXXX hXhX�X�Xh(h8hHh�hHxXxhxxx�x�(�(�Xhx���((((8(H(X(�(8(8 H8#X8h8#�8 �8H(H 8H#HHhHxH#�H �HX(X HX#XXhX#�X �Xhhhxh�h�h�hxx(x8xHxXxhx88�( 8 H X h x � (0�0(@H@ h@ x@�@(P8PHP XP �P8`H`#X`#h`#x`#�`8pHpXphpxp�px0x0�   0 @ P ` p � � � 0�0�0@0@ @@P@ `@�@P P#0P @P#pP �P �P` `#0`#@`#P```p`�`p p0p@pPp`ppp�p�p�p�`�`�(8HXhx��((�(8(#H(#X(#h(#x(#�(#8(8H8h8 �8H8H XHxH �HX8X XX xX �X�Xh�hx(x8xHxXxhxxx�x(h(h�  ( 8 H HXhx��� ( 8  H x � 0(0 x0 �0 �0@@(@H@X@h@ x@�@PHPhP#xP�P�P`H` X`#h`#�`pHpXp#hp#xp�p�p�(�8�H�X�h�#��X�h�x�������� 0@P`p��  �  0@0P0 `0p0�0 @@@ p@ �@ P0P@PpP �P�P0`@`#`` p`#�`0p@p#`p#pp#�p0�@�P�`�p���� � �(8HXhx�((8(#X(#x(#�((8H8 X8 h8 �8(H8H#HH hH xH#�H(XHX XX hX �X(h8h#Xh#xh#�h(x8xHxXxhxxx�xXHXH� ( 8 H HXhx� 8  H � 0X0 �0@8@ H@X@h@ x@�@P(P#8P#HPXPxP�P�P`(`#8`#H`#h` �`p(p8p#Hpxp �p(�8�H�x�����H�X�h�x�hPhP�(8HXh( h x � � 0(0H0X0#h0 �0@X@ �@P(P#8PHPXP#hPxP�P#�P`H` X` h` �`pXp#hpxp�p�p�(�8�H�X�h�(p(p�(8HXh(8(#h(x(�(�(8(8 88#H8 h8 �8H8H#HHXHhHxH�H#�H�HX8X XX xX �X#�Xhh(h8h�h#�h8xHxXxhxxx�x�x�x�h�h�(8HHXhx���((( H(h(#x( �(8(888#H8X8#h8x8#�8�8H(H HH hH �H �HX(X8X#HXXX#hXxX#�X�Xh8h Hh#hh�h �hxx(xhx�x(�8�H�X�h�x�������XHXH�@P`p�� (0(@(�( 808#`8 p8�8 H0H#@H#PH pH �H X0X@XPX#pX �X@hPh`h�h`xpx�x�xphph�(8HXhx��(X(#�(8888 H8X8 h8x8�8H8H HH#XH#xH#�H �H�HXHXXX hXxX�Xhh(hXh#�h(x8xHxXxhxxx�x�x�x�h�h� ( 8 H X h Xhx��� 8  H #X h � 0(080 H0#X0#h0#x0 �0@@(@H@#X@ h@#�@�@�@P(P HP XP hPxP�P`(` H`#X`#h`x`�`p(p Xp#�p��(�8�H���H�X�h�x���pp� 0@P``p���(0( @(P(#`(#�( �(8@8 P8#`8#p8�8H0H @HpH�H �HX@XPX#`X#pX �Xh0h Ph#`h#ph�h �hx x0x@xPx�xP�`�p�������  �(8HXhx��(X(�(888 H8#X8 h8#x8 �8H8H#HH XH#hH xH#�HX8X HX#XX hX#�XhXh�hx(x8xHxXxhxxx�x�x�h�h�(8HXh ( h x � � 0X0 x0 �0@8@H@#X@h@#x@�@P8PHP#XPhP#xP�P`8` X` �`p(p8pHp�p�pH�X�h�x���xpxp�(8HXhx��(8(#�(888 H8#X8 x8 �8H(H#8H#HHXHhH#xH�H�HX(X HX#XX xX �Xh8h#Hh �hx(x8xHxXxhxxx�x�x�(�(�(8HXhx�( 8 #H #X  h #x #� (080#H0#X0h0#x0#�0(@H@ X@ h@ �@(PXP �P(`H` X` h` �`(pXp�p(�8�H�X�h�x���xpxp�(8HXhx��(X(#h( �(888 H8 X8#h8 �8 �8H(H#8H#HHXHhHxH#�H#�HX8X HX XX#hX �XhXh#�hx(x8xHxXxhxxx�x�x�h�h� 0@P`p���   #�  � #� 000@0P0`0�0�0#�0@ @#@@ `@p@ �@P@P `P�P �P`P` �` �`�`p p0p@pPp`ppp#�p#�p#�p`�p�������````� �� q� d� _� d� q�    K� T� _� d� q� d� _� d�    K� q$� 8� K$� G� K� T� d� _� qH�   \�����}�����   .�T�}�������}���   .��$� ��.$��.�T���}��H�    �	� �	� �	� �	� �� �	� �	� �	� �	� �	� �	� �$� 	� �	� 	� �	� � q	� 	� �	� �	� �	� �	� �$� �� �	�    �	� �� �	� �	� �� �	� �	� �$� _� _� _� q	� 	� _	� _	� q	� 	� _$� �    � � �	� �	� 	� 	� �	� �	� $� �� �	� �	� �$� �� �	� �	� $� 	� �	� �	� �	� �	� �	� �	� �	� �	� �	� �	� �	� �$� _� _� _$�    q	� _	� T	� d	� _$� _� _� $� �	� 	� �	� �	� �$� �	� �	� �	� �	� �	� �	� �	�    �	� �� �	� 	� �$� 	� �	� �	� 	� q� T	� _	� 	� 	� q	� 	� �	� �	� �� 	� _	� T	� K	� _	� q	� � 	� �	� 	� d	� _$�   }� �	�T	�}��	��	�}	��	��	��	�}�.	�T	�    �� d� T� Y� d� d� j� j� � � �� �� ��    �� �� �� �� � �� �� �� �� �� �� �� ��    �0�    �� �� �� �� �0�   � �� �� �� �� �� �� �� �� ����.�   .�T�h�.� ���.�.�T�T�h�T�.�   0�   T�h�h����0�    �� /2�   �





		�
	�

		�
	�L�V�`�l�p�~�����������ܮ  �2�2�]�  ���y�!���  &�  j����j�����  �Z����Z���  j����j�����  �Z����Z���  ³  ϳҳ���1�ƴʴȴ2�h���Թ
�      �
  ���
�
�
����      8     888        �     ���  >>      �     ���  >>      �   �������>>      �   �������?>      �   �������?>      �   � ���  >      �   �� ���* >      �    ��� � >      �    ��� �>      �   ������>      �   ������>      �   ������>      �   � �
��  >      ��* ��
(������
      �   8� ��    8      �#  ����  >  �      �#  � 
�?  >  �    ���꣪�� �����>����    �������� �����?����    ������� �� ���?����                                                                                                                                                                          ����� *������
���
��* 
 
�� �#��8 �#8 �  8�� �#��8 �#8 �*�*8�⨊����( �#8���/��8
�������� �#8����8(� �����"�#8 ���8�� ���� *�#8 �  �8��� ����(�#8�
�  �8�� ����( �#8 8�  �8�
� ����� �#8�:�  �8�+� ������#8�?�  �8��� �����
�#8 ���8��� ����8+�#8 � �*8��� ����8,�*8�*�* 8�� � ��8  8 � 
 :�� � ��8 
 : પ��>�� ����:���>��������� ���?�������� �� �� �� �� �� �� �� �� �� �� �� �� ����, ��������> :�*8��8?�8 �8�+8�8�?��? �?��;�:+ 8��>������> 8��8��8 �8�8��80 8��8�8 �8��8��8 8��>��    |  �  � �5 �5 p p�\s\s�p�=WU5�= p p p p �����: 8��:��� ����: 8��8��8 �8��8��8��8 8��:��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���ة�� ���  ��� �� � � � � �ߍ& ��"  � t ���� �� �� � ����� ��� ��XL �H�Z�r � � �P0� � � � ��  ��z�(h@H�' )�	� � �# �$ �% h@                                                                                                                                                                                                                                                                                                                                                                       ���  �� W� |� ,� �ũ�w  Ré �$  `� g� �� �� �� � �� �ѩ�S  n�r �s �  ��� z�������%�  � }�l ���L�®  ���LG©��h L[����"�  � b�l ���h�  ���LG©��h L������  � G�l ���B������  � #�l ���,LG���� �$  `� g� �Ьt ���L�L0���� Y�LG© �$  `� g� ,� 6�v ��� �� � 9� ,�L� K�w �� �� d� ,Ǯ  �� ,� �� �� ,�L� 5�L�H�Z� �u �x �y �z �{ �| �} �~ � �� �� z�h`H�Z� �c ��� ��� ��� ���� �� �	 �� �  �Ĭ� �r� 4ɭ� 8��� �ܩx�� ���� �� 8��� �	 �� � � �c ��� ���  �ĭ� 8��� �	 �� � ��� ��� ��c  �Ĭ� �D� 4�L�� 4� 4ɭ� �	 ��� �� � � �c ���  �ɭ� i�� �  �ĭ� � ��� ��c  �ɭ� 8��� �  �ĭ� �l� 4�L,� W� �� ��z�h`xH�Z�c 
����� 轎�� �� �
 �� � �	 ���� �i�� � JJ��- �� i� � i � � � � �Ȁ��
 �
 � �
�� � �L��z�hX`H�Z��S  n� �ȩ�d � ��"�� �"��	 �"��c  r�����z�h`H�Z��S  n� �Ĝ_ �X� �`�	  � ��_ �_ �
� ,�L�ũ�c  rˬ  ���) ɬ  ��� ɬ  ��� ɬ  �����c  rˬ  ��L�����5 ɬ  ���� ɬ  ���� ɬ  ���� ɬ  ���� ɬ  ����LV� 4� �ȩ �$  `� g�z�h`H�Z�  ɩ �S  n� �� UǮ ��)�r �s � �k �  ��� ���� GƬk ���� �L� � � �z�h`H�Z�r �=Ll��s �r �s ��Ll� pƩ��k z�h`H�Z Ré�w ��u  �� �ќm � �  �� v� J� H� v� J� �� v� J� �� v� J� �� v� J� {� v� J� �� v� J� �� v� J� �� v� J� �� v� Jɩ�  �� v� Jɩ �  {� v� J� {� v� J� w� v� J� w� v� J� w� v� �z�h`H�Z�r �s �r �=���s �s ���r ��r �s z�h`H�Z���g ��� �(�	 ��d � �c  r˜ � i�  � ɩ �  ��� � ���  ��� L�Ȭ  ��� L�Ȝ �H� ���	 ��d � �c  r˩ �  4� 4� r˩�� �	 8��	  r�� � �%��  ��Ќ L�Ȭ  ��� L�Ȝ �X� ���	 �!�c  �ʭ i � �"�c  �ʭ 8� �  4� 4� 4ɩ � �!�c  �ʭ i � �"�c  �ʩ�� � 8� � �	 8��	 �!�c  �ʭ i � �"�c  �ʭ 8� � � � �8��  �Џ� L�Ȭ  ��� L�ȩ�d � ���� ���	 ���c  r����
�  ��݌ z�h`H�  ����h`H�Z� �@� � � � ����� ���z�h`H�Z������ ���� ��z�h`H�Z�/���� ���� ��z�h`H�Z����� ���� ��z�h`H�Z�?���� ���� ��z�h`xH�Z �ɭ i�  �ɭ 8�� z�hX`H� �  �ĩ�� h`xH�Z� �  r˩�� z�hX`H�Z�  ���� �� 4� 4� 4� 4����I� �  nѩ�� � �0�&�	 ������ �n�	  nр���� ���	  n�L�ɭ 8��  n�L�����J� �  nѩ�� � ���'�	 �n����	 �0�  n�L�ɩn�	 �0�  n�L�ɭ i�  n�L����L�ɭ	 �n�L�ʭ �0���u L���H���u L���`���u L���x���u L�ʩ�u L�ʭ �0���u L���H���u L���`���u L���x��	�u L�ʩ
�u z�h`xH�Z�` ��
 �c 
�� �� � �� �	 ���� �i�� � �b Nb Nb �b �- �� i� � i � �` �` ��Ȁ���
 �
 � ��` L�z�hX`xH�Z�` �c 
�� �� � �� �
 �d �
 �	 ���� �i�� � �b Nb Nb �b �- �� i� � i � �` �` ��Ȁ���
 �
 � ��` L��z�hX`xH�Z� �� �c 
�� �� � �� ��� ��� �	 ���� �i�� � JJ���� �� N� N� N� N� � � � � �� � - �� i� � i � Ά �� � �	ȭ� �� ��N� N� N� N� ȭ� - �΅ �� � �	��� �L�z�hX`H�Z��c �f � �!�A�	 � �  nѩ�� �W�	  nѩ��f ��W�	 � �  nѩ�� �A�	  nѩ �f z�h`H�Z��d � ��I�� �I��	 �I��c  n���!���d � ��:�� �:��	 �:��c  r����䩄� �"�	  �� r� � � ɩ�d � ��j�� �j��	 �j��c  n���<�� ��z�h`H�Z�w ����c L������c L�����2�c L�����3�c L�����4�c z�h`H�Z�u � ��0� �n�	 ��c  n�L�Ϭx ����$� �c�	  �Ϭy ����<� �c�	  �Ϭz ����T� �c�	  �Ϭ{ ����l� �c�	  �Ϭ| ������ �c�	  �Ϭ} ����$� �{�	  �Ϭ~ ����<� �{�	  �Ϭ ����T� �{�	  �Ϭ� ����l� �{�	  �Ϭ� ������ �{�	  �Ϯx ����0� �n�	 ��c  n�L�Ϯy ����H� �n�	 ��c  n�L�Ϯz ����`� �n�	 ��c  n�L�Ϯ{ ����x� �n�	 ��c  n�L�Ϯ| ������ �n�	 ��c  n�L�Ϯ} ����0� ���	 ��c  n�L�Ϯ~ ����H� ���	 ��c  n�L�Ϯ ����`� ���	 ��c  n�L�Ϯ� ����x� ���	 ��c  n�L�Ϯ� ������ ���	 ��c  n�z�h`xH�Z�` �	�d ��c �c 
��j�� �j�� �
 �d �
 �	 ���� �i�� � �b Nb Nb �b �Q�� i� � i � ȲQ�� i� � i � ��
 а� i� �,�c �c 
�� �� � �� �
 �d �
 �	 ���� �i�� � �b Nb Nb �b �Q�� i� � i � �` �` ��Ȁ���
 �
 � ��` LxЩ�d z�hX`H�Z �ȩ�d � ���� ���	 ���c  n���l�� ����� 车��	 车��c  n���*�� �f ���t �  ���� �� 4� 4� 4� 4���� �̀��� �̀���Ҭ	 �A����t L%ѩ �t L%�z�h`xH�Z�c 
��j�� �j�� �
 �d �
 �	 ���� �i�� � �b Nb Nb �b �- �� i� � i � Ȳ- �� i� � i � ��
 Юz�hX`H�Z � �Ӯw �� '�L#��� n�L#��� ��L#��� ��L#��� C�z�h`H�Z�u 8�
��⑍ �⑍ ��d � ��� ȱ�	 ȱ�c ����#��j  r��LG�z�h`H�Z�u 8�
����� ���� ��d � ��� ȱ�	 ȱ�c ����#��j  r��L��z�h`H�Z�u 8�
��
�� �
�� ��d � ��� ȱ�	 ȱ�c ����#��j  r��L��z�h`H�Z�u 8�
���� ��� ��d � ��� ȱ�	 ȱ�c ����#��j  r��L�z�h`H�Z�u 8�
��2�� �2�� ��d � ��� ȱ�	 ȱ�c ����#��j  r��Lc�z�h`H�Z� ��Б� �Б�	 �Б�c  n�����x� � �	 ��d �$�c  rˬu �
���� � �c  nѩ�� �u �c  n�Lԩ�� ��c  nѩ�� � �c  nѭw �c ���  n�z�h`H�Z� �l ���i �g � �m �n �o �p �q �r �s �j �  �! z�h`H�Z�a ��d �h ��� ��L�ԭg ���D��c  4� 4� �ɭ 8��  �� `ɩ �  �˩��  r��a �a �� `ɀϩ��g L�ԩ�c  4� 4� �ɭ 8��  �� `ɩ �  �˩��  r��a �a �� `ɀϩ �g �m z�h`H�Z�a ��c  4� �ɭ 8��  �� `ɩ �  �˩��  r��a �a ��L�Ԝa ��c  4� `� �ɭ 8��  �� `ɩ �  �˩��  r��a �a ��L;թ��g � �h z�h`H�Z�a ��d �h ��� &�L֭g � �D��c  4� 4� �� �� `ɩ �  �˩�� � i�  r��a �a �� `ɀϩ �g L֩�c  4� 4� �� �� `ɩ �  �˩�� � i�  r��a �a �� `ɀϩ��g �m z�h`H�Z�a ��c  4� �� �� `ɩ �  �˩�� � i�  r��a �a ��L1֜a ��c  4� `� �� �� `ɩ �  �˩�� � i�  r��a �a ��Ln֩ �g � �h z�h`H�Z�a ��d �g ���1�
�c  4� 4� �ɭ	 8��	  r��a �a �� `ɀ���g Lש�c  4� 4� �ɭ	 8��	  r��a �a �� `ɀ� �g �m z�h`H�Z�a ��d �g ���1��c  4� 4� �ɭ	 i�	  r��a �a �� `ɀ���g L�ש�c  4� 4� �ɭ	 i�	  r��a �a �� `ɀ� �g �m z�h`H�Z�a ��d �h ��� p�Liحg ���Lح 8��  4� 4� vɭ 8�� � �c  r˭ i� ��c  r��a �a ��� 8��  J�L�ש��g Liح 8��  4� 4� vɭ 8�� � �c  r˭ i� �	�c  r��a �a ��� 8��  J�L%ة �g �m z�h`H�Z� 8��  4� 4� vɭ 8�� � �c  r˭ i� �	�c  r˭ 8��  J� vɭ 8�� � �c  r˭ i� �	�c  r˭ 8��  J� 4� 4� vɭ 8�� � �c  r˭ i� ��c  r˭ 8��  J� vɭ 8�� � �c  r˭ i� ��c  r˩��g � �h z�h`H�Z�a ��d �h ���  �L�٭g � �L�� 4� 4� vɭ i� � �c  r˭ 8�� ��c  r��a �a �� J�Lz٩ �g L�� 4� 4� vɭ i� � �c  r˭ 8�� ��c  r��a �a �� J�L�٩��g �m z�h`H�Z 4� 4� vɭ i� � �c  r˭ 8�� ��c  r� J� vɭ i� � �c  r˭ 8�� ��c  r� J� 4� 4� vɭ i� � �c  r˭ 8�� ��c  r� J� vɭ i� � �c  r˭ 8�� ��c  r˩ �g � �h z�h`H�Z�a ��d �g ���L#� 4� 4� �ɭ	 8��	  �ɭ	 8��	 � �c  r˭	 i�	 ��c  r��a �a �� `�L�ک��g Lp� 4� 4� �ɭ	 8��	  �ɭ	 8��	 � �c  r˭	 i�	 ��c  r��a �a �� `�L)۩ �g �m z�h`H�Z�a ��d �g ���L�� 4� 4� �ɭ	 i�	  �ɭ	 i�	 � �c  r˭	 8��	 ��c  r��a �a �� `�L�۩��g L)� 4� 4� �ɭ	 i�	  �ɭ	 i�	 � �c  r˭	 8��	 ��c  r��a �a �� `�L�۩ �g �m z�h`H�Z� ��� ����� ����� ����� s� � �r �s z�h`H�Z��d �g ���l� 8��  � vɭ i� �	�c  r˭ 8�� � �c  r� � vɭ i� ��c  r˭ 8�� � �c  r˭ i� ���g LKݭ 8��  � vɭ i� ��c  r˭ 8�� � �c  r� � vɭ i� �	�c  r˭ 8�� � �c  r˭ i� � �g z�h`H�Z��d �g ���l � vɭ 8�� ��c  r˭ i� � �c  r˭ 8��  � vɭ 8�� ��c  r˭ i� � �c  r˭ 8�� ���g L3� � vɭ 8�� ��c  r˭ i� � �c  r˭ 8��  � vɭ 8�� ��c  r˭ i� � �c  r˭ 8�� � �g z�h`H�Z��d �g ���{ � �ɭ	 8��	  �ɭ	 i�	 ��c  r˭	 8��	 � �c  r� � �ɭ	 i�	  �ɭ	 i�	 ��c  r˭	 8��	 � �c  r˭	 i�	 ���g L9� � �ɭ	 8��	  �ɭ	 i�	 ��c  r˭	 8��	 � �c  r� � �ɭ	 i�	  �ɭ	 i�	 ��c  r˭	 8��	 � �c  r˭	 i�	 � �g z�h`H�Z��d �g ���{ � �ɭ	 i�	  �ɭ	 8��	 ��c  r˭	 i�	 � �c  r� � �ɭ	 8��	  �ɭ	 8��	 ��c  r˭	 i�	 � �c  r˭	 8��	 ���g L?� � �ɭ	 i�	  �ɭ	 8��	 ��c  r˭	 i�	 � �c  r� � �ɭ	 8��	  �ɭ	 8��	 ��c  r˭	 i�	 � �c  r˭	 8��	 � �g z�h`H�Z�	 ���� �i�� � �b Nb Nb �b �� � � i � �� z�h`H�Z��� � � �] �	 �^ � 8�� �	 i�	  C� �� E�] � �^ �	 � ��� ,�L*��� ,�L*�� ��	�c  r� � ɩ�c  r�L*���0� ��� &�L*��� &�L*�	�c  r� � ɩ�c  r�L*���L���r �s  �l ��� ��L^� � ������� � ����� z�h`H�Z��� � � �] �	 �^ � i� �	 i�	  C� �� E�] � �^ �	 � ��� ,�L��� ,�L�� ���c  r� � ɩ�c  r�L���0� ��� &�L��� &�L��c  r� � ɩ�c  r�L���L��r �s  �l ��� ��LC� � ������� � ����� z�h`H�Z��� � � �] �	 �^ �	 8��	  C� �� E�] � �^ �	 � ��� ,�L���� ,�L��� ���c  r� � ɩ�c  r�L����0� ��� &�L���� &�L���c  r� � ɩ�c  r�L����L��r �s  �l ��� ��L� � ������� � ����� z�h`H�Z��� � � �] �	 �^ �	 i�	  C� �� E�] � �^ �	 � ��� ,�L���� ,�L��� ���c  r� � ɩ�c  r�L����0� ��� &�L���� &�L���c  r� � ɩ�c  r�L����L��r �s  �l ��� ��L�� � ������� � ����� z�h`H�Z� �U�� � �1�y��� �&����� �� �� ����� �	� ���� z�h`H�Z� ���k� �g��c����[� ���� 8��  C� ��C���� i�  C� ��.����	 8��	  C� ������] � �	 i�	  C� ��z�h`H�Z� �U�� � �1�y��� �&����� �� �� ����� �	� ���� z�h`H�Z�j � �L(�i � � ,ǩ�c  r˩��l z�h`H�Z�i ���Ld� ��� H�L����� {�L����� ��L����� &�L�� ���  Hԭ i� �#�c  r˭ 8�� L�����  {խ 8�� �#�c  r˭ i� L�����  �֭	 i�	 �#�c  r˭	 8��	 L����� &׭	 8��	 �#�c  r˭	 i�	 � ����i ����j ���i ����i ����j � �i  v�z�h`H�Z�i � � � �i ���L�� ���Ly� � � ��� ��L@���� R�L@���� ��L@���� w�L@���L@�� LN�� �L@� ���L1� � � ���  �׭ i� �#�c  r˭ 8�� L@����  R٭ 8�� �#�c  r˭ i� L@����  �ڭ	 i�	 �#�c  r˭	 8��	 L@���� wۭ	 8��	 �#�c  r˭	 i�	 L@���L@�� L��i ���Lh� ��La� ��2�j L����(LT�� �L�� ��L�� ����j L����Ly� ��� �i ����i  v� �  �	 �! � �" ���# z�h`H�Z� ���L/� ��L�i ���L� �  gܭ 8� � �#�c  r˭ i � �j L��� L��i ���L$� �  g�L���  g�L�� ��Lp�i ���Lh� �  gܭ 8� � �#�c  r˭ i � L��� LH�i ���L�� �  g��j L���  g��j L����i L�� �i z�h`H�Z� ���L� ��L��i ���L�� �  Oݭ i � �#�c  r˭ 8� � �j L|�� L��i ���L� �  O�L|��  O�L|� ��&�i ���L7� �  O��j L���  O��j L��i ���Lt� �  Oݭ i � �#�c  r˭ 8� � L��� LT���i L�� �i z�h`H�Z� ���L�� ��L��i ���L�� �  7ޭ	 8� �	 �#�c  r˭	 i �	 �j Lb�� L��i ���L�� �  7�Lb��  7�Lb� ��&�i ���L� �  7��j Lj��  7��j Lj�i ���LZ� �  7ޭ	 8� �	 �#�c  r˭	 i �	 Lj�� L:���i Lo� �i z�h`H�Z� ���L�� ��L��i ���L�� �  =߭	 i �	 �#�c  r˭	 8� �	 �j LH�� L��i ���L�� �  =�LH��  =�LH� ��&�i ���L� �  =��j LP��  =��j LP�i ���L@� �  =߭	 i �	 �#�c  r˭	 8� �	 LP�� L ���i LU� �i z�h`H�Z�# ���L�� �  ��	 �! ��" �  0� �� �# z�h`H�Z� �] �	 �^ ��d ��	 �m � �LP�n � �$�n �n �c ���  nѩ�� �	�c �m  n�La�o � �/�o �o �c ���  nѩ	�c �m �n ���  nѩ��  n�La�p � �K�p �c �c ���  nѩ�� �	�c �m �n �o  nѩ��  nѩ��  n�La��m �m �c ���  nѭ] � �^ �	 ��d z�h`H�Z� �] �	 �^ ��d ��	 �m �
L$�m ��� � �c  n��n �n �
L5�n ��� � �c  n��o �o �
LF�o ��� � �c  n��p �p �
LW�m �n �o �p � �c ���  nѩ��  nѩ��  nѩ��  n�Le�m �c ���  n�Le�n �c ���  n�Le�o �c ���  n�Le�p �c ���  nѭ] � �^ �	 ��d z�h`H�Z�r �=L���s �r �s ��L���c  � � r� � ɩ�c  r˜r �s �  ���ש�c  r�z�h`H�Z�u �����x LG������y LG������z LG������{ LG������| LG������} LG������~ LG������ LG��	����� LG��
����� z�h`H�w i�w h`H�Z� �$ �%  `� g� � � � � � � � �O �P �ߍ& z�h`�$ ���Q�% ���.�0 � `�) �* � �  W�= � g�6 �7 � �  ���0 �0 �+ � ��= �= �8 � ��% ���.�J � `� g�C �D � � � �  ��J �J �E � ��`�& �'�) ȱ'�* ȱ'�+ ȱ'�, ȱ'�- )
�����. 转��/ Ȍ& �0 �1 �+ � �'�2 �T�' ȱT�( � ��' � ��2 ��Ȍ2 �& ��`�@ �A�C ȱA�D ȱA�E ȱA�F ȱA�G )
�����H 转��I Ȍ@ �J �K �E � �#� �%  `� g�) �* � � �6 �7 � � `�3 �4�6 ȱ4�7 ȱ4�8 ȱ4�9 ȱ4�: )
�����; 转��< Ȍ3 �= �> �8 � �'�? �V�4 ȱV�5 � ��4 � ��? ��Ȍ? �3 ��`H�Z�, )?	@�M �, 4��-M �M �1 �.��- )@��J��M �M Ȍ1 �.����1 �- �1 �M �O �� �O z�h`H�Z�9 )?	@�M �9 4��-M �M �> �;��: )@��J��M �M Ȍ> �;����> �: �> �M �P �� �P z�h`H�Z�F )?	@�M �F 4��-M �M �K �H��G )@��J��M �M ȌK �H����K �G �K �M � �O � �P z�h`� �O `� �P `�S 

��<��T ȹ<��U ȹ<��V ȹ<��W � �T�' �V�4 ȱT�( �V�5 �& �3 ��2 �?  � �� W� ����$ `����A ����B �@ ��L  �� ���% `�X 
�����A 轨��B �@ ��L  �� ���% `� � � � � � � � � � � �( �) �* `Hڮx ���F�y ���?�z ���8�{ ���1�| ���*�} ���#�~ ���� ����� ����� ������v �� �v �h`H�Z�� � �
�0� � ��  ���� �(�	 ���  �� 4ɩ �  ��� �ɭ �%�. ���� � 8i(�	 �
� ���  �� 4ɩ �  ��� �˩	� � � �2 ���� �(m �	 � � ���  �� 4ɩ �  ��� � �ǩ� � �
�2 ���� �(m �	 � � ���  �� 4ɩ �  ��� � �ǭ � �) ���� � 8i(�	 ���  �� 4ɩ �  ��� �Щ
� � � �+ ���� �(�	 � � ���  �� 4ɩ �  ��� �� ɩ(�	 �� �� �/� �
����� 轶�	�)�� � �
 �	 ���m � �i�i � � ���� 0� 4��� m � � i � �
 �ǭw i
����� 轶�	�)�� �d�	 �� �� �� ���  �� �z�h`H�Z�
����� 轶�	�)�� � � �� i� � i � ʀ�z�h`H�Z� �
 �	 ���m � �i�i � � �- ��� 0��� m � � i � �
 ��z�h`H�Z��d � ��~�� �~��	 �~��c  n������z�h`H�Z��d � ���� ���	 ���c  n���?��z�h`H�Z��d  �� ��M�� �M��	 �M��c  n���l��z�h`       ��  �        * � 
      ��  �       
� *           ��  ��            <<<<<<<<<0�   <<<<<<0���  <<<<�<�?<?<<<<  <<<<0�0<<<<  �<0< <?<0<0�  �<<<<<<<<<<�  <<<�� �<<<  < < < <   < <   <0<0<0<3<3<3�  �<<0<0<0<�  <<<<<<<<<<<<�  �������  �<<<<�< < <   <<<<<<�?<<<<<<   �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  � ��� ���   �  �  �  �  �  ��  �� �  �  �  �  ����������� ���   �  �  �  �  � �� ��  �  �  �  �  ���� ��� �� �� �� �� �� �� �� �� �� ������  �   �   �   �   ?  ��������  �  �  �  ������  �  �  �  �  �������0181@1H1P1X1`1h1p1x1�1�109�90A�A0I�I0Q�Q0Y�Y0a�a0i8i@iHiPiXi`ihipixi�i�i,$,,,4,<,D,L,T,\,d,l,t,|,�,�,�,�,4�4<�<D�DL�LT�T\�\d�dl$l,l4l<lDlLlTl\ldllltl|l�l�l�l�l8@#@@H@P@`@$h@ p@x@�@"(X0X8XHXPXXX`XpXxX�X�X�X$<,< 4<<<D<L<T<$\<%d<l<t<|<&�< �<�<"8L'@LHL PLXL`LhL$xL�L ,\(4\&<\D\(L\T\d\l\t\|\�\�\"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 W� ���