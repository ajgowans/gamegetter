���  � � � � � � � � � � � ��" ��d`� ��@����'� ����0e�� e����`�


 n��
e�� e�`d
&
&
&
&��
&e��e��@e�`H� ��hHJJJJ ��h)	0�:���H�Z�Z�Z z�z�z�h`8� d
&
&
&i����e�� Z�� ��� �� ��0e�� e�z����8��~����`����������N�N*N*L9�N*N*N�N*N*LQ�N*N*N�N*N*Li�N*N*N�N*N*L��N*N*`        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l���  �U�L��� V�� ��������������� ��L��`

����� ���6����C����,0)�*��,��)��+����i�nL��ȩ �)�*�+�,L愭��e�nL������������  I�� �
>��`�	H�
H�H�H� �� � � � � � � � � 	� 
� � � � � � � � � � � � � � � � � � � � � �Сh�h�h�
h�	`��	e	�	E
�
���&E�m `��L����� ����������� ���L��`�	�+� �
� �����
m�
��� � � � �	`
�
m�� �b��
������	`� 8� � 8� � 
�@@ 
��<� ( �$� ���@ ��H���)����� �������i��i ��i��i ���ة)������ � �����ɨ��`�Z��J� �JJ��͇e �!�·i �"�H� �!hz��#�$�



e��i ��JJJJe�� ���m��� ��ȱ��i�� e��i0��i ���� t��$�#`�����0�� iɪ�骍�`H)�����hJJJJ�
ei@}���` 0`��� P���@p��      )AYq�����1Iay������@ � � �Z�	�)��
�*���+���,�L�)
��	�%�
�&��'��(Z ��z�)�	�*�
�+��,��+)*� y�z������Љ`�)�%�*�&�+�'�,�(�')i��')Ji� �0�d�%�'m:H���E�h ���(JJe��i ��&�



e��i ��'J�jJJJe��()�#� � �,'p�����0�� �ڪ�������#�!........��߬ �Q����e��e��m ��i ���L�` @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��H��
���


�h 놭���`��Ջ����  <  0       � 0         � 00�  <�8��  �  �8��  �  ��  �  �  �  �    �    �        �  �  �  ��  $0   0       � 0         � 00� �  $
�B�  �B�  �    0    ��  �    �'������  6�<�        
    
    �<�        
    
    �"    "    "    "    
 $  $ 
 $  $ 
 $  $ 
 $  $                 ��  "�� 0 ') 0 ) 0 '��) 0 ) 0 ') 0 )) 0 0 ''0 �"    "    "    "    
 $  $ 
 $  $ 
 $  $ 
 $  $                         
    
    �         �#��7�����  :
�؎�؎�1��  %
�W�
�W�
	�		
	


	
	
��Hژ��1
�h�%h�$`�@�A� �@H
��ȏ���ɏ��� ŏ��G`l�Ώ܏ꏢ �@� �����`� �@� �����`� �@�( ��������@`� �#�Y� �#��)�� �+��� �+��"�� � � �( ����`d# ��!���+���(�Y�#��` d��#��`�(t#���!�+��L��+�,�-� � �,�$��������1� �.�G�,��4�5�6�#`�#�`�4��L�����5��5�`� �4�6m+�5�1�
�.�	�.�� L������$�*�%�+�4� �*0LO����LR����Lk����� �1����� ��*�6m+�5 �Lې��� ��*�K�*8�K�*�+� �+Lې���Lr�����,�,�,}���/�*�0�+ �Lې���- ��*H ��*H�,}���*�/�+�0�,�,h�+h�*Lې���' ��4��� �*�M������*i�*� e+�+�4Lې��� ��*Hȱ*�+h�*Lې���2���O)��O:�O� �P� ��*��ɓ�4�.L�� � �Lې����4��)��O)�O�O�O ��4Lېɀ�(逼�

��ғ�M�ӓ�N�ԓ�O�Փ�P ��4Lې�4�G�����I�� �}�� �O� �P�  �� �*��ɓ�4�. ��4
��*�$�+�%�4��G��G��`�3��0��0�L��� �(���� �3L����� ��(�W�(8�W�(�)� �)L��

� ��(��ɓ�0 �����( ����) ���)�* 	�* L��   �*��+`�(��)`H���K
�LhJH��mL�LhnLnK��L�K`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   � ���������  ��� ���[��/���� 2�� Z�h�Iw� z������� ��� ��L��`�������������_^FNNEzz#W4W2Yw� ��� V��S���� ���
��� V������ ���L���(H� � Z� ��z�����e����������C��������`e����h:м`��� ���Jjj(**HJ~�~�~�~�J~�~�~�~�hJ~�~�~�~�J~�~�~�~��ж����`            x   �   ?�  ��   ��   �� ��� ��?� ��� aÁ� aÃ� aÃ� Ã� �Ç� ���� ���� ���  ��  ��� ��� ���  ?�  �   �        �   �  �               � ��������  0�                   p   | |  | >  ><>  <><  80  ?0  ? g�� ����� � |p 0w� 8�����~s�  s�  � 8��������g   w   �   �  ��` /�p x<x |x|~ <x|g <y�g�s�c��`��`� � �?  �   �   �    @                                                                    ��             ��                                                                                                                                                                                                                                                                                                                                         {|      {|          ��      ��        {|  {|  {|  {|      ��  ��  ��  ��            {|    {|          ��   ��                 {|               ��                                        34                  GH                              ��                ��                                                                        �  ��  ��  ����  ����  ����  ����                                            {|  {|  {|  {|      ��  ��  ��  ��                                                   {|  {|  {|  34      ��  ��  ��  GH                                                   ��              ��                                   34                 GH                                                     �        �    ��  34��34  ��  �  �GH��GH�  ���  ��    ��  ��  �  34 34 34  �    ��  GH GH GH  ��  �  �  ��  �  ���  ��  ����  ��  ��  �  ����  �    ��  ��������  ��  ���  ��  ���������  ����  ������  �  ����  �    ��  ��������  ��  ���  ��  ���������  ����  ������                                                                                34���  �����GH������  ��������34�������GH��������������343434�������GHGHGH�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ������������������                                            ��  ��  ��      ��  ��  ��    ����  ��  ��  34  ����  ��  ��  GH    ��  ��    [\  �  ��  ��     op  ��������    34  34�������     GH  GH����  ��      ����  ��        ����            ���             ������      ��      ���      ��      ������        ��    ���        ��    ������              ���              ������                                        ������������        ������������        ����  ������    ����  ������  ��  ����  ������  ��  ����  ������    ����  ������        ����  ������        ����  ����    34  �����  ����    GH  ������  ��    34  �  ����  ��    GH  ��  ������    34  �  �������    GH  ��  ��        34        GH                                                                                                                                    ��    ��        ����    ����        �[\+,+,[\�      ���op?@?@op���    ���+,+,���  ����?@��?@���������+,��+,�����  ���?@?@���    ���[\+,+,[\���      ��op?@?@op��        ��    ��        ����    ����                                                                                            LM�                �������������T��7����������Q]!H�H@!��!H @ 0 @ 0 p@0s        3      0</ī    3�0� 4          ����*          �3     A¡����Z      >: `  `hkkk   
:::8      ���k    � @
��       �  ��       � ��
  4 � p�7@      >��� �2�¡8���P� 0�	 �2(ʩ2��Q�
�**�ʣʣ*��*�
kkkhU`T `8:::
BL AZ�� �(���  P  >@TA  Q�*�� �   UUTPQ��3     @UA�k�<0T UUTP  7�p�  s0@pU0U@T0 @3 C@C  @7�p�P4P  �>@UA  E��   �T UUTP  T�
��  UA  ����T UUTP  �� 
��               � � �    �</ + �0�>   � � < � / k P��%(%J(*�2�<"   �@���T� � ^ ^^^^ �   U@UPT�T�T��  U�	`�    U@UPU������QU  U UU�?�j   T�B`���Zk  U UPO>��    @������ P ������   U@UPT�T���k   � @
��   U@UPUTUTU�?�*  U UU����UE  U�T`R�	&T@  U UTSO>� < o����� > ���          ���9m��x  ��            ����H�  �� 
�����!P� kZ���� J�  ��>CP!U � ������  H  U�  ��? TUU!U � ��T�P�H U�  � �`�	 � T T�T�P�H� ŀ� 
P^^!^� @T&�	`�P  ��>CP!U � �? TPPHP U�  ����
�    U � ��T�P�H U�  ���@�   �        � �0<+�X  ���  � �      0 < <�,��bT�COLLOA   p q@qPpT ll    W WP^^   T@UPUPT�T�C   �a�  N   T@UPU�3�"�"Q   U UUO�?E   B@ � ����K   T SC<
1   p@ kkk k   @ zzz@z   T@�P�P�T/T`K   � J���   T@UPUPUT<�(U   U U���2Q   T�T`R����/   U UUWp8�R��K%�P���    � �         ?B�#j�Z)F�ʠ�	 �� ?      k  kk k�  p@z@zz:� # 0
�$��`<  �N@PPT� * �"�"�3    T�  ��? @PU� * �<P�PH T�  ���c�	    llP Hq p�p r@^^TW� # ����`2� $P   �@PU� * �( < P H T�  ��2��  @� * T@P�P<H� Ā  ����V 	�
      @ p � o��̦@Ujj���a��Zhoh         ?����� < ����+� ��     ��VP���d�X�     � jWk�@    D�"PP�`   @ a X	�@ P�j�Z�j�����^     Q�j�n�o�+   � $@�  @ ��
      @ �   � �@UPWh�d��} V ZR	a	��U     `'          @   	3�      � *���������J   � ��
�
 (�"   � � � � *(*�h  
 �  �
�
�*�*��O���&`���� ����� >      <b��������(����: : > ?       ��P�P�xV藠��� 
VYef�
�� ( X^ ��xa�g���� 
@ "� Q��� ( @Րڐf�n���+��
Z_�j�k�o���� �@�$!�"H� �  
X(b� )�Pc����T�Q>�  i9Q9�3�,��  � @� $         A	 
@@    �j( ������ �    �
�*�
�
�� 
   �B�����* � � �  )*�(��� � 
   UUUUUUUUUUUUUUUUUUWUWUWUWUWUWUWUUU_U_U_U_U_U_U_UUUUUUUUUUUU�U�U�U�U�U�U�UUU�W�W�W�W�W�W�WUU�_�_�_�_�_�_�_UU�������UU��������������      �� � �<77�6�6�6�7  �<����\�p?�   �
`'X�X�X�`%�
���������������������������?�?���� ?   ? �������?����?��� ��< � � � � �����������0�0����00�� ?��������������?��< ���  �00 �����?��� ? 3 3 0 0 �?�? � ����������?  �  0 � ?����� � � ���?��� ? � ? � �����������              ? � ���?� ? 3   3   3  ?�� ����������������� � � ������������� ����0���3����0�0�����������������?��<������� � �������������� <�0�3�3�0<��� ������������?�   <   �  � � � ������������?0�����0��������������������� �� � ���������������������� � � � � � � � � � � �����������0� � � � � � � � � �0������������?�  ?  0?�  ?  ��������� ? ? ? ?�?�? ? ?  00������?�  ?  �?0  ?  �������� ? ? 3 3�3�3 ? ?  00���� � � ������� ���� ���� ����������0000000����������3  �         �        ��00   �0000�   ����         �        �  �300   0�3 0 0 3 0�   �������� � � � ��� � � � ���������00 � � �� � �� � � ��0�0�������� � � � ��� � � � ���������00 � � �� � �� � � ��0�0���� � � �������?� ���?� ���?� �������������?     ? �����������  ?�     �  0 0�    �     ���0�0 � � �  �   �  � � �00�   �     � 0 0�     �  ?  ���0�0 � � ������� � � �00����0?0??�?�? 0 ? 0 ������0�0���? ? ?�?�?�?�?�?�? ? ������������0 ? 0 ? ?�?�?0?0����0�0���? ��  ��  ��? �����������????0� �? ����0?������������< ? 3  �� ?0   �3�������?�?�� < ?�<�<�< < � ������� ������ 3 3 3�3�3 3 � ������������ < ? <�<�<�< � ��?�?��� ������ ? ?���?�? � �����������������?� �   ��������? ��� 0 000 0 0�� ��?33���� �   �?����������������? � ������� � ��?33��������� � �� � � �����������?�����0� 0�� ��� � �0������3�3�3�� 3 <<<� < < 3�3?3���30��?0�� � ����� � ���?�� �3�3?3�� 3 < <<�< < 3�3�3���30��?0�� � � ��� � � ���?�� ��������?�?�?������������������?�?�?��������������  �?�������?�������?��  �?�?�?�����?�����������  �����?���������������0�0�00�0�?�?�?�?�?�?�?�?���������������  ��  ������������ � ������������� ��3 30303?3 �� ��� � �<� � �����3�3����?3������0��<�������������?������������� ������� ?��������������?�������������0�������������?�����������������  ������������ � ���3 30303?3 �� ��<� � �<� ��� ���3�3�?3?�??��?��?������0���?���                                                                                                                                �������?�?������������?�<������   �  ? �       �������������?�� ? �� � � ����� ��?   � � � ��� � � ���?��� � � � � � �    ������ � ��             � � � � ����� � � � �          ? ? ? ? < 0     �3��?�?������������3�?������������?����       � � � �� � � �   � � � � � � � ������� � � ��  ? ������ � � ���   � � � � � � � ��������                 � ����� � � � �      < � � � �            ?                            � � � < o����� >    � � < � / k P ���9m��x         � �0<+�X�R��K%�P���        0 < <�,��b?B�#j�Z)F�ʠ�     @ p � o��̦��O���&`���� �         ?�����<b��������(����  (
�)�*�*�
��  P �@Z��Z@� � � � � � � � � � P�
�*����������X�h�`����� j � � � ��h�j�j�j�j�j���������( �          �</ + �0�>���         ��%(%J(*�2�<"��              ���  � �  � �         T�COLLOA	 �� ?     @Ujj���a��Zhoh���� >       < ����+� ��: : > ?         i ��j           ��
�*�*�*�*�*�
�
��� * 
    ? � ���������� ?        P� �j�j�V�V�F�&���V�����      QQ�����V���&�&���V����EQEQ    � �����V���&�F�V�V�j�j�  P   QQ�����V��DD���V����EQEQ   � � � � l `    Z X  Z X  Z X        (���EQEQEQEQ���(        D�V��e�e�e�e�a�a��U�U�U���� EQEQ����hUhh�hEhEh�hhU����QQ �����U�U�U��a�a�e�e�e�e��VDEQEQ����hUE��EUEU��EhU����QQ   ����������     EQEQ�
���UU����
EE      ����������    EQEQ�
���������
EE  & � � � 9 	   � � % � � % � � %         *���nP�P��n��*        P�Z�
YZYZY
YZIZI
PZUZU
UZ�Z�
 PEE�*�*U)TY�UQUQ�TYU)�*�*EQEQ P�Z�
UZUZU
PZIZI
YZYZY
YZ�Z�
PEE�*�*U)T)R)Q)Q)R)T)U)�*�*EQEQ�  ؅؀؅؀؀����U�U��    EE �����%�%�%�%�%�%����     ���U�U�����؅؀؅� � �EE ��  ��QU�?�?QU��  ��      @@@�� _ �@u  � M@s        3|A�}�V�ep� $���O�uP��w4�    @@���[����V�[� �� U   � ��[�V���V�[ � �Q  Q  ����[�V����[� �@@ U   � ��[�����[ � �Q  Q'T  'P''R'R'$�jURUR� P   TQQ @�  ��UE����UE��  � @PDPD T   P�URURj�$''R'R''P  'TQQ @�VXXXXXXV� @PDPD     Q � �b� m�0       �014O]O��XU��d] }1�10 DDD? �D�C�C�C��C�C�D?D�D*  DQE  @E? � ������� ? @T  UT D*D�D? �D�C�C�C��C�C�D?DD  DQE  @E? ��#�#�#�#�#�#�? @T  UT       �	�	�	          � T�     ���`	`	`	`	        �T�T��@ p`ll`p@       ��:UU�:�@ @ ````@ �        �
VU�
   �	  �9�9  �9�9      ��"EQ�"�@ @ @ @ @ @ @ @               UU  ��\U    �?U5 4(44 4(4  �� LULJLJL@LU  �? 0U1i1A1U1i1  �� LL
 
 @L  � 0E0hA1 )        �	`�      ( 
`X� %   p ��&�9`�         �	`� &     �`!K	� �      @      \U��  4 4(44 4U5�?  LULJLJL@LU ��  A1U1i1A1U1 0�?  LL @H@ @@ ��  @T0)11E   �  ���^U^���^���jUW�^�^yy���^�Ve]�~����^�^�^�Ve���j^U��Z^U���j���^�^�^�^���Z^�^�yyyy�^�^�WUU���^���^^y^�V�UUUUUUUUUUUUUUUU     � 
� ��       ( � �  UP��_����@� �UU�UU          @ � �@���T������� T@����_���� _ ����@  U������U��P������� UP�����������U���U    UU�����������@U@@@AG�� � ��  
 �    � � (       � � @    UU��UU ������U ���W�����U�������P�����_��@� T  P����_  �U������U�������P������������UU�U    U��U�������A���U�������@U��                     	
         !"#$%&'()*+,-./012  3456789:;<=>?@ABCD EFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������                                                                                                                                                                                                                                                 � < 3 3 �     ��    CՌ�    ��   A@� �    � � ����    ��LLA�T C    �� DD�Y    ��L�\���     � 0A�UW     � � � ��    ��  D@_p�    ?�0�0�0�?�     ��  A@CU<U    � T D0    �����D�_p    �� A�U5            ? � � � � � � ���������0 0 0�  0 ���      ��S�\�     �0������0�0�0�0.� � � � � � � � 0 0 0 0 0 0 0\֜j������<��3 � ??< 00�5�5�7�?�?�<�0�0 �         � � ���Us��?�?���5U7_������3              �        ]���� � � � � p�� ��0�p�q�q�p�p�WT ��?         �            � � ��0�0�0�004\PW�T� � � � � UUU� 0 0 0 0 0�� ��W4U�� 00T�D S \L�0�0�0�015U4U1U4 0 0 0  ���|�W�  ��� 5 5 �?     � �U0S0\�_  < 1 1 � ?U5     ��p�OWUU�D ��\�L�\0LW�PU? 5 1 5 1 5 1 4 �� O �        UUUUUU��        � � � �          � �            LULUOT��        UEUAU ��        �\�\_�        UQUUUE��        0��         U5T5P1�?        sUsU<��        UU�        �U��A��        U5U51�?        �Q�U� ��        AUT ��        UDUA��        5 4 4 ?              � � ��p0\    ��@UAUU��0     < �G5\1       � < ���0p    �� AU=��     < � AS    ��|D3 3DsAsU     0 0 � U     �  L C�0T    �?Q0 0D40U    ��< 33 �L    �� D��4    ? �5@�G�       � 0 0 0 0    �� U�T    �P4@04�     � < s 3 3 s    ��    QD��    ��  @ TDQW�    �? 0 0 01O0o����s�3�303030��� � �      p5p5p5p5�?      0|������ � � ?0?0��    \5�?������ � � �W�?����0�0�0�0U�?�������0<0W�����?�?� 0 <U� � � � � � � 0?p�������0�0�050?0=0?03��    �\����?��  0 �              WW�������?303T�U������33�  s sss�� =  W��335�1�5�5�?�  30s0����WS0S�\         = ��UU       0 <�75U5�@�G0L0p��  ��5050��T}�� 0�p�\5\1GT�0�0�0�0�0<0\�<��03��0�� 3 3�0�00000� p� � � � � � DQ=�0�0�0�000L�D��0000�4�4�501��p 0p0Qp\� � ��0<�3�0_0�  \�� � U�     �0W�L�p04 0 � � � U<U5     ��GQ�                _ \ �          UUUQWU��        U5U=�           < �          UWT\U��        U� 5          �E�T���        QUU�         L \ \ �        U5T5U5�?        3sT<Q��        ��UUUU��        S�U5U�         0W0W� �        UU@�        0W0W0��        U5T54�?        W0C��        UEU@@��                    xH�Z� ��  � �� ��� �� � E	�	�e
�
�E*�z�hX@@�s����#���C�ӡ���؎	� �d  R�  �� �� �� M������х��� �)��� �� 2� Ȇ�e � ���������	 ��� )��������)�S����L��Ѝ�������И _Ѭ���Ѝ�� ���јi _���L	�@@@@@@8  0@P`8@@@@@@p�����Т �*�	�,8��,�����p��*�	�,i�,���������i����ɀ�L��d � ɴ�
������Lu�

���ѝ*��ѝ.��ѝ2��ѝ6���)�-i�1�5���,�4i�0�8� �+�/�3�7`	
+,)*78'(56%&34#$12!"/0 -.                     � �              �     D3�L0�L3@� 1DD33DD            � 1@L�03D1���1 D 1��0�1� 1  � 1�@  D 1� 1� 1�D13@���3 D3��03��13�L13D3�3D    D 1�13��13��13@D 3@L 3@L3�L33 �  �           �          �  @    ��L 3�1�1� ��0� 1� 1� �1���� 1� 0�L3@�   �0�3L  �D1� 1� 1� ������13�L13��13���    D3���13��1� 1� �L33�L33�L03�L          ��           �    @�03�03�� 3 ��L           @  � 3��L���� @�3�L0� 1�  L 3�0�  � 1� 1� 1������ @�03��13�L13���3�    D�1�L13��13�� @L 3@L3DL3�L     �   �        �          0 �      DD13DD3 � 3�0�3D 03�D1� 1� 1D 3���@1� 1�0�� 1 D  @�1�   1� 1� 1� 1D ���@13��13�L13��13DD3D    �3D13��1�@1� 1D 33�L33�L13�L3@D  �� �)��� �� 2�����c �� ȅdT oߩ���W��������W���f�����������&�����T
��=о>� �� �� �� �� �� *� �ک �� Ȇ������ �������� �������� �������c ���袌 d� �� �� � �� �� �� � �� �� m� � u� >� �� �� �� �� ,� M� � X� �� 5� ��������ة ��� )�)��� -�������� ��� )?������L2֥T
�������� ��Zȱ�[ȱ�\ȱ�]���p ���q ����������������%�)�-�9�=�A�M�Q�U�a�e�i�r�y������������������������������������$�8�L�`�����"�6�J�^��v�}������������������������������U�����Ȟ���� �� �P���s Y������������������T
�������� �


���


� h��$P����H�i
�h�����$P0�H���h���`H 	� 	h 	� 	`� ���V��`)�  �ة�EP�P�)� �ة�EP�P`� ��V��`�$P0JJJJ
���R��S��R�ȱR�L��L����%�����L���Lu��L/��L��`��
��e�t��R�u��S��R)
�����2�f��gLٹ*�f�+�g����
i���r i�w `�����T��


����`�]������`�����t��K�u��L�K)�������`�����K��T
���M��N ȅJJ)��M


� �K ȅ)����T

m��C���K���K`
� �)��� ������� �٬�������� ������`��������� Tڥ`������`��������������P����b R�������)H��JJJ����� ������h����L�������`��������������P����b R�������)H��L:ڤd�� �	� �� ���d`��N�N�#��V�$��W� � �V��V�N�N�T
��Q�X�R�Y� �X�U��
�N�N�#��V�$��W� ���V�ȑV�N�N�`��
��#��V�$��W`���U�� �ڠ �VI)��V�B���ܱX


�MȱX


�N��8�M�M� � JfM��8�N�N� � JfN jۅJ� �V)�J�V`�M
.�N
.�MI�i�M�NI�i�N�M�N.�)����` � �V)��V�`8�V)���V�)�VL�۱Vi)�V����ܱX�ȱX�ȱX
��I��J����e���L� $*
"%(+.147:=@ȱVi�ȱVi� h�I���I�V)	`�V8`����VHȱV�JȱV�K���L���M��h)0JJJ �I�`�Ii���8�V�� ��L9ܥU
H��#��V�$��W��I�V "ܰ ��h8��L�ڤI�VH)8��)ݍ�*ݍ�+ݍ�,ݍh) ����qV�V��qV�V`���9��E��F��G��H�Em��Fm��Gm��Hm����`   �a �� K�� ��   � a � � a �    ��� K�� �a  �  ���K�K���� �]�� �V)��V�`��V8��V0`� �V ȅjjj)c��Ui�V��V0O)`�K��V
�O

	���V���܄M�X


�Oy�ݠ�V�M�M�X


�Oy�ݠ�V�U����ȱX��ޠ�V`������  
�U
H��#��V�$��W�J����ȱX��
޽���M����N��I�V/)8J��M�ȱM��IȱVɟ�� �ȱV����hHJi0 ��h8��L�ڥ_)�`�U
H��#��R�$��ShHJi0�r � �F� h�h8��L��  ? @��_�]�`��]�^J����^�_9����^�_9�ޤ^�
L����J�L�ި���������Z��[�L���h� �]�2�`��a R���)	`��������������%�)�-�9�=�A�M�Q�U�a�e�i`STAGE��TANKS�� ��� �)��� �� 2����	��b��߅ ������ V��c ��d ���	� V��T ����� ����`���`�\��]�`��ލ��ލ��ޅH��ޥZ


�L�L�[


�M�M���H�I�Ry-JJJHȱR�JȱR�Kh �b�Ii��R)�JJJJ��]8��]��LZ�I�R��&)	`�Rh`�������Z��[��T���� �Lߪ)��JJ)	`�Rh`�IeH�h:0L�`         �TIMES OUT ! �����������b�`�_)���b�` R�� �)��� �� 2���� ���������� ����e � ��dc�c0Lm�(�E���F���E��F�������� �  �� ���F�F�H� ��L�ȅG�_)�	� �
�G� ��L;� �)��� ����� �������Luխ�


����������� oߢ��L�ե]�`�_)���`�*�`)��a`�ai
��t���u����)��`��` R�� �)��� �� 2��T��L;� ��������T oߢ��L��YOU HAVE COMPLETE ��ATTACK IN THIS GAM��E.��  BUT NEXT SECTOR ....�� �)��� �� 2���������� ������ d���e � ��� ��� �����Lu�PRESS START BUTTON Copyright 1991,1992�  Thin Chen Enter.��&Ņ�'Ņ�(�� ������ d������~��� ��� �������� ��� ��� �� ���� R�L2��� ��` ����� ���_ �� I����� /�� �)��� ��L^� )�`�y���� )��s�������L��     �PAUSE� GO!��\�`�_)�`�����_)��s�������L��	�  ���R)��R $�����Lb�����Lb���T��Tٳ�����H��Tٸ�����I����$I&$H0*�h 0 8��h ��`$H�_)?�����Lb��h ��R�8�R��R�  ����R�qR��RLb�`���� �� )��L��  ���R)�	�R $�����L�����L���T��Tٳ�����H��Tٸ�����I����$I&$H0*�h 0 8��h ��`$H�_)?�����L��h ��R�qR��R�  ����R�8�R��RL�`���� �� )��L�� ���R)�	�R $�����L������L����T��Tٳ�����H��Tٸ�����I����$I&$H0*�h 0 8��h ��`$H�_)?�����L���h � �R�8�R� �R�  ��� �R�qR� �RL��`���� �� )��L�� ���R)�	�R $�����L������L����T��Tٳ�����H��Tٸ�����I����$I&$H0*�h 0 8��h ��`$H�_)?�����L���h � �R�qR� �R�  ��� �R�8�R� �RL��`���� �� )���R)���R)��i�R`�]����R)����R�:ȱR8��R�6 ȅ)?	 i� ȅ)��Rȭ�R ȅ)���R)��R`8��R`��R)��L����L/���Lu�L���R)
�E
�F 9��F�F�E�F�X� qR��F�Y�qR� h�E��` �� � � ���=���9�)��dP
&P
&Pm��PFPjFPj��JJJJfPm���$P0JJJJ`)`�`�N��G��
���G�2�G�t��E�u��F��E)���N�ȱR�JȱR�K� �E�LȱE�M ���G�G�`��N����N��N�R)JJJL��R)��!�L8�J���M8�K��w�K8�M��mL����!�J8�L��Z�M8�K��R�K8�M��HL����!�M8�K��5�L8�J��-�J8�L��#L��K8�M���L8�J���J8�L��`8`��R)�������
�R)

�L�����R)

��C���D���e�L��R)

��_)��ȱf�ȱf��e�� �R�ȱR���������_)JJ�N�)�N��L����R)��+���*����������Ly��R�:�R`���`Ly�]����R�:�R` ȅ)�`��F���R)��
�i��F�`�����(�RL���R��R)
�E

	����R)�R� �R�Ey �G��R�Ey�H�ȥG�RȥH�RȄB��R)�C�T

eC��C��B�R`� ��F��E�R,)JJ��p�ȱp��EȱRɟ�� �ȱR�����r ���Ei��r�F�`��H��I�R0�Ii��H�`���?�NȱR�JȱR�K���L���M ��L��Ii��R)���8����� ��L��I ��(��EH)�8���Nh)N�EL���\�\h���EL��I :����I�R)	`�RLY�I�R�)��)������&�ȱR8��RLY��ȱRm�RLY�ȱR8��RLY�ȱRm�RLY�ȱRi�ȱRi� h��`�����L\�8`��`�L������	� ����� ���8�
 ����� ���� ����� ��EP�P�$P��)�	��8�
 ����� �)�	i���`�T
�����s����t`��s$P0JJJJ`)`�K�
���M��N��)���M)���i
�L��������9��	��L��
��u��Q��� �uLj���M��u�=� ���	���	��U���ܱX��ȱX������0���L�L��a���`ɀ�� G�L��	
��������� G�L�� G��K�L �� �M��E��MJ�L�<8��L�5��M�ݪ����L?�N��M}����� ���	���	� ⅥL�a�u�G� ���	���	��U���ܱX��ȱX���
��#���$��� ��L���Ϣ��	)�� ��L��8����	�8`!"2	�	���	� �K�
��8�
L��
$Pi��8�ȝ�	���	���	`�E�P�B�C�D���)�JJJJ�F�)�G�F��P�J�E$P0



H�$P��9���h�����EP�P$P0���ХJ�P�F��i
��Gо�B�C�D�P`�_)�` ٩�F��E�R�)�G�)�)���)`�H ��h8� � �EG�R�Ei��r�F�`� �� ���JJJJH��������E�R)�JJ�Ȍ�R�y��� �� ���h����L��R�y������r

��  �i��w

���ɟ�� L��*��,��)��+`�_)�`������	)���8���`��	)��	LJ���	0��	
�� �����	


���	


�ڠ���> �����	�LJ�ڽ�	)�JJJJ�L�M�)�N��	���	�� �)��� ����ȩ ��	�M��ȩ���	�L�M�N�����	�����ԅ�	� ��`�_)�`�����R�&)��#`��������R�)��R8��RJJJL9�`�R:�R
H�� ���� �R�hH��� G��h�����RLg�R�����eL���� 4H\
�"�.���������������
��������"�%�(�+�.�1�4�7������������������������ ���	��������!�$�'�v� v��w�@w� v�  � ��  � w�  ����� ��v�� ����� ��w�@ �@��@ �@x�  � ��  � y�  ����� ��x�� ����� ��y�@ �@��@ �@z�  � ��  � {�  ����� ��z�� ����� ��{�@ �@��@ �@|�  � ��  � }�  ����� ��|�� ����� ��}�@ �@��@ �@~�  � ��  � �  ����� ��~�� ����� ���@ �@��@ �@��  � ��  � ��  ����� ����� ����� ����@ �@��@ �@B�R�b�B�r�v�z�~������������������������������������������Zn�nZ�HZn��nZ��p\�Hp\��\p�\p��  � &:�:&�H&:��:&��<(�H<(��(<�(<��Nb�bN�HNb��bN��dP�HdP��Pd�Pd��2F�F2�H2F��F2��H4�HH4��4H�4H��
�
����
�
����  �Vj�Xl�Xl��8�8�=�D�K�K�Z�i�x�x������ �����"{|����}~����"�����������"������������"+,�?@�-.�AB�/0�CD�12�EF�34�GH�56�IJ�78�KL�9:�MN�"����	��
��� ��!"��#$��%&�"ST�gh�UV�ij�WX�kl�YZ�mn�[\�op�]^�qr�_`�st�ab�uv�
  )�-�1�5�9�=�A�E�
 {�{����a�h�{����������
	
		  




	
	
��������	


		pw~�������������                        00  000 000 000 @@0 @@@ @P@ @P@������������������k�3�������S��                        33     � 0  �  � 0  �     33                                                                                                                                                             o   o     �   �    o o o o   � � � �      o  �o     � ���      ��  o    ��   �   ��        �        �         �       33        0        0        33                               � �� �� ��                      o o o o   � � � �                         ���
�  ����                  30 �      0 �      0       30         
�        �                            DD    � �@� �  �@� � � DD � �  �
�   � ��� �     � � �� � �     � ���� �   ��� �� ���     � ���� �   ��� �� ���                                        DD� @���� ���@�DD����������������������������������������������������������������������� ���������                      � � �  DD � � �  @� � � � @� � � � DD � � � �  � � � � ���� � � ���� � � ��� �  � �� �  � ���      �      F���   �      �   ���    �      �  ���              ���                    ������    ������    �� ��� DD �� ��� @ �� ��� @ �� ��� DD �� ���    �� ���    �� ��  � �� ��  � ��� �  �  �� �  � � ���  �  ���  � � �    �DDDDD    �DDDDD                                                              DDDDDD          ��  ��    ϯ��   ������  ��DD�� ��@�����@��� ��DD��  �ϯ���   ������    f      ��  ��    DDDDDD                                           2����	�[��	��	��	d ��	� ��	����	 ?� ����	�����	���� i<� ��`

�� �7�� � �����`� �/ ���	���	`���	��	�@�]�<��8��	 ���i0��i ���	����������i0���i �����	���  ����	�a�1�]�-�D ������ȑ�� ��� ��i0��i ���ߩ��	� ��	�_��a�Ș "���	�a�����	`��	`��	���	`��	�M�]�I��8��	 ���i��i ��i0��i ���	����������i0���i �����	��� ����	�a�1�]�-�D ����ȱ����'��� ��i0��i ���ߩ��	��	�a�����	`��	`



}������i ��J��� �����e��i ������`���� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?��������� ?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                           ?������I�& LM����<�