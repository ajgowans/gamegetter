  �� � ��P�u�u ���䁅F�偅G���& �P��� �F�H��w���Few�F��G�x� ��LP��u�u��	 ��� �P�˩��&  �� �����& ��'� �P�P���'��)������-���`��x� �w�x�	�
8�	�x�wL���w�x`� �u�v�u�w��I�z��H�}����I�G�H�F�v����� ���v�H�Hƙ���u�u��˥w��A�G���F ���
��A�G���F ���x��A�G���F ���w��A�G���F ��� �u�C�G�u
iхF�u���� ���u�u���F�G��F� �u���w�w�
�
8�
�w�uLN��u��� ���F�G��F�w�� ��`ACF��  
 �u�́�I�؁�H����w����x`



IJKLMNOQRTVWb�9��ɫͬ+���pp\5\5W�W��UU�UUpUUpUU\UU5\UU5WUU�WUU�  �UUUU  � �UUUU <     � �_UU� 3�    � �UU�? 3|    � |�UU= 3���  � _�W�_� 3 7�=? � _���W� 3 ��� � _�W�� �� �����W@�W�0 |;� ��}  @}�����:� ��    �� 0 ��0���p    @LU]��?��      4\U��*8��      �p���*<���  ������0���?  �@�T������0?  �@��������U��|�p 0?  � WUUUUU�\�P�/\�p �?  � WUU�_U5p5U�?_� �?  � _U�W�u���W� �?  � 4w��P\����W� 00   ����TU�\}U?WW 00   t���TU1p���ܥ 00   tZ�TWQ�U��ܩ �?  � �j�TW� W�_� �?  � �jW�U \5��� �?  � �jW�U p�<�� �?  � �j�� �U � �  ����5��  Wu �       ��?�W  \��      � �v��WWpU_�^      < �v�(���U��z0    � � �_5 WU�z�  �� �@�� \U�z0< ��� @�T�   pUU������ @�}�   �UU� ��5 P�  WUU �_W �UU�\UU ���  �UU5pUU]  �  uUU�UUu�    ?]UUpUU��  ��WUUpUUUW�  ��UUU\UU�U�W�UWUU\U���_�_��_U5W�_U�����_U�W5Wu����UU��V]��U]����W�U���z� �U]����Wթ���zUpU�z���Wե���zUpU�zZ��UU����^U\U�^��]UUuU��WU\UU�j}]UUu���UU5WUU���zUU]��zUU5WUU���zUU]Z��UU��UUU���zUU]j��UU� �UUU���zUU]���UUUpUUU���zUU]���UUUpUUե��zUU]���WUU\UUե��zUU]���WUU\UU�W��zUU]���WUU5WUU����zUU]���WUU5WUU}U��zUU]���UU��UU՗�ժzUU]��^�UU� �UU}��j�zUU]����_UUpU՗�j��zUU]�Z��WUpU}��j��zUU]��~��~U\�W�����zUU]������W\u������zUU]������^5W]������zUU]������z5W�������zUU]�������������������_UUU�������������?  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � ������&   � f�� �'�C������������[������& � �P�P���')�� ����������� ^�涥���� ϘLT�` <V� �'��� �P�P���)���')��淥��(��`��������4淥�i�����汥�������L���𥲅F���G ��淥�i����` � � 
 � �� 
  ���
  � ���
  �������������������������������������������������������������������������������������������������������������������������������������������������������������������                ����_U_U_U_U_U_U����UUUUUUUUUUUU�?��U�U�U�U�U�U� � � � � � � � ��U�f���f������?UUUUff��ff������U_U_U��of������        UUUUUUUUWU�_<p p � �            UUUUWU\UpU�U�UpU��               3��0 ��0 �D0WU\Up�p=�      �33�30�30DD��  u���������UUUUUUU_��5 5 � 5 5     � �P�<�C\]Ww\wWw\wq]��  �U_�zu�W|U�UUU�U]UU�W?| �        3 �U1W�|��7Ww\ww��]w��  }��W�u���UUU�U_WWUU�UW\\�         �<p�UUU]�wUwuw�]��3  WU|��_�^���UUU�U=U_�                � �@�\eq�q��9��ww��  U��u����U�UU_Up��5 7 L � � ���0�L�9dN���S�>eC�Tf���q�q�q<�  }�˫J�J��UUU����? @UUUU�8�8�8���䩣���c���c�����U{U����V3�  U�_?�:[:|��UUUUU}��=  9 6 � � �d�9N�N�9e��Ow0}sw��}sqsq��  �ի�j�k|U�U�U=U3U�U�U�U�U�UUUUWU\U\UpU�U W W | �       � �f��_�p���3�q�q?�  ���������Uw���< �\�WUUUUUUUUUUUUU��]_UWWU|_��     � ���=CUTWuUuUuu��  ��/o*e+e<��=\| � 7 ��U|UWUWUU�� 5 5         � 0 � U� <�տ߹��;|U�}U�U�U|UWUUUUUUUUU��u}U]UUUUUUU�U�U5W5|�       @DDDt��U�00           U�U��=��g������UUWU|eÛ>|ٛ������ W��V�v���U  DGD<�G<O ODOD�O�PD��D��D��|���_U_U_��    U�W�]�U�U���� �����UUWU|����=W����UUU��5 ��w�����UU�U W W W�UU�U�U�U�U�U�U�U�����  � \\� 3 UUUUUUUUUUUUUUUU?^�^^U~U��|��W��뵮���k�[�����z _ \ W W ����5�5�5w5u}���� W�             � ��������C���WUUUUUUUjuo����?                   0        �?�� � � � � � �� �W�?=0C� � � � � � ����?            ����      ����        ����      =CU��鿫�����PU_U_�_u_u_u_�_W�]���u�uon��of���j���j����  7������ 7 �� PUUUUVWU]UuVuUuU]UWU_UuU]]uU�W_�VM�~]��fu����           � �P?U�W|U�UUU�]�U�U�UՕUYUUUUUUUU]��DD��^���������������
����?     ���T_�UuUuUu]u{�~W�{�z�^�_�^�W�UU�U_ե��DD=��h�h�������f�����������b�   � < � ��������  ? ���  5 5��]W=��u^u�թu�u��������             � ���� ���?��� � � ��?��� � ���?�?   � \\�_z}z�ީ^���W֥j�������U�U� ���U�0 0 � 0��0�0���æé�^�zU�W���<p p \W�U_��W�^�_�z�ꪪ������             � �PU�UW��]W�W�W�WWW�]U]Uu�uU�UUuUUUUUUU�UWU^U^U0 � � � 0 ��T]UUWUU_U�uUWU]�_���W{~�魗�~��ժժU�e�U�V�UՕUUU             <��3LUqU�UUUUuUUUW��W��W����~��~�ꩪ�맾���������� ppp���<PCUTUUUU�UUuUUUUU��U������������������������������        ? ��UUUUUWuUUUU�UUUUUU��jݪv�ڪڪڪj�j�j�j�����C���cD��$�C`S�����                1 1 � ��?�@USUTUTWUUUUU�UU�UWUWUWUU��5 Of`�YU��_�U]�]W���� 7�70L�S �UUU��(��`j��������U_�p�STV��ff��               �� UTUUU]]UU_UpU�UWWU�U�U��5U5Տ5POUP�Ue��ff��U�T\W�W�\0�? � �� �U�U�U�]�U�U�U����P���d���f�   ��\W_Cu<p� �  ��UUUU��0    ��UUUU ��}   �U5UP1��?��U�U�U�U��D�����UUUUUUUUDD����_U_U_UU� �����UUUUU��D����UUA�<L�3�DD�����U_W�WU] �G  � 0 �             �       �00��  �     ���� ?    ����    < �� 0 �0��         � � � � | s�t0}pw������ W | � � \ � � \ �����     0 0 � �3�< � ���3�N�^���^����5�5�5�5���uw�]�]�uUwW�W�                ��_UUUUU�U���������               � <�C0T�� W��?TW��  UU��_Ujկ���0+L�\�\�q�ׯ]�]k��?�@�W | � �yp^��p}������������շ����������      �� _\��_���P=UC�T��4M�S5�����������������?��?�@�U]�w_��U��5 �]�� �� � ���� ��������         �=��?�W�UQ��  WW�U�����Zo�ׯ}U���������UU? ��@U? ��TUT�CU=U��]\��w��WW��W\�\U��pup]�������������������������]    uV    ����]   qv{����� �]cglrw|���������`dhmsx}���������aeinty~��������pbfjojojojoj����k^�������ʼL����X]  �����˯�R   ]    ����_�    ]   �����zNSV  ]   ����ΠOTW  ]    ����YPU   \[[[����ИQ[[[[ZIHJF	MMMMMMMMM-27;K
M!%).3M<G?"&*/48=?#'+059?DCB $(,16:>E@A@A@A@A��
���������� �����P���$������������������3���9� �8 �����?���> Π淥�i����Ƹ�ӥ�i�����汥��p��`�C����������������������F���G��� ����i����Ʒ�⥰i������ƶ��`�C���F���������_���G���F��� �����G���F��� �������_��`� ������t�C���F�������� �P�P���')�򥱅G���F���(������ ����i�����Ll�涩 �P�P���')�򥳅G���F���_������ ����i�����L��� �� ��t�L^�� ���G������� �P�P���')�򥱅G���F��� �0�� �����L� ��`��� � ��� � �
�		 � � �� �'� �P�P���'����`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �$ :� � ��� ��'������& � �P�P�� =��)��
�'����ƭ�婀�& `�')�;������I����H�����G� �F�')����F� �F�H�����Fi�F ��Ƭ��`���������	�
8�	���L��� �L�M�L�d��I�g��H�j��N�M�m���I�G�H�F ���M �� ���N���L�L��ɥ���W�G�T�F ��������W�G�X�F ��� �������Y�I���H���	�
8�	���L������I�G�H�F ���H�H����I�G�H�F ���[�I�ԅH� �L�L����I�G�H�F ���H�H�L�L���ƨ`WY[H�� 
 ������I����H���� � �H� =����������� ��Ƭ��`MJGFA����      <   �  �� ����?<��?��������� ��? �� �� �� ��?     ������ ��? �� �� ��          �   �   �   �  ��  ��  ��   �   ��$
�����6����7����8����9� �:�@�;���0��1��2� �6�3 ���:�>�;�? Π�6��7�:i�:��;�2���2�:iX�:��;�;�0�0��о�1�1��ж`�3JJJJe9�=�3)



e8�<��=`� �������<�>�>��?�����>i.�>��?����`��                 �  ����  -"IWes���������   .<JXft���������  ""=KYgu���������  "0>LZhv���������  "1?M[iw������"��  $2@N\jx���������  %3AO]ky���������  &4BP^lz������"��  '5CQ_m{������"��  ""DR`n|���������  ))ESao}���������  **F"bp~���������  99GUcq99999999�                                                                                                     ��                           ���pլ�lի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի�kի������������������    ���������������������������������Z���Z�������������������������������������������������������j�گu�����������������������������������j�گu�����������������������������������������������������ꯪ��������������������������    ��������������������������Z���]��v�ڪj������  < � ���?�?�������������������������������������]���Z��������������j��j����������������]���Z���������������       � ��<�������������j�ڧv��v�کj���������� � � ������� � �    ��������������������������j�ڟvu�ڧj��������������������������������z�z�z�^���z�^�^�^�W�W���W�g�W�W�W�g�W��ZW�W]��z�^Ɦ_��y�y�y����k�n�n�n�z�ꪪ������������������������������j�ڧv��v�کj��������������������������    ��������������������������  ������������z�^���^�[�ezUzV^��[�ה�V5UU�eVUU�eU��� ����[�[�k��U�fu�ZU]�}Y�U[YkU�Y�uUUU��W5��_u]�gUUUUYfUUW�����r�_�V�U�e�W�g�^�v����ꆪ������ꪪ�������������������������������j��j����    �����������������������������_�zU^e�UUՕ=YC�T5UMUS���W \�>�CTUU_�p5����u�uW_�U_YuUv}^�^�Wו}U}U�o�_5�7������Y{U{Y{U]�eW\o�]mWm�nW�}W�� ���~f�U�V�e�V�UUefUUWV_�wV�UGoG�G:G:N:�:�?���� ?    ?   ��Z_��_Z��������    ���������������������Y_UU�eYU��5TM�O���U|�^�W��|���%7�L�c�h���U���UYUU��]V]UueuUՕUUe�W5�v]՗�g\U\VWe�UU�YeUV��W�_�]]W]�]W�UUYY�e5W-�-WcYcUc�Rْ�ꝺ������������խ�߭������﫺��������������j��e}ߗu�������    �����������������ozU{�_U]�m��?�0�0GW��m�k�[��TPUUUUUUU���TfWU\�pU�e�U]U]�WU��U�e�V�U�Y�յ5�-�-�+{+{��������������U�Y�U�ի����k�f�i���z�^���W�U{Yz�^V^U^V^U{U{f{U{�{��ջ[�^���n���^�^�^�^�^��ꪪ����}�֧j�������    ��������������eeUUU�YYUe�W?��s�p3� �(X�hX�X�X�Y5�6���U�U�UE��WU|YA�UՕ�Y�U�ٛ�ٽy�]藸U\U�e\UWU[YWU�UU�YUUYUU�UWe\UlYx���ڵ۵{m{m{m{�_՗YUU�uU�Y�UU��\�p�q����ͽ����V�V�s�]UUYVU��������������������������������    ��������������UՕUVeUUUYeUU�� USUTUZU[���P5V�ZVkV�VUZY�U}U��U�C{S�^^C�P�T�UՕy%v	uՀ٠U+�Ue�UU�YUUUU�5W5g-�m�[�l�l̰����r_���5W6�-\m\[�[�l�l��l�o�mƵ�77�5-Um�[U[U[�-U�Y���������������������������������    ����������������U�UU�UYeUUUUoU�eWU\UqWU|U�g\U�UUV��UV��C?PTUA�P%T	u̀��+�
�� ( 
�0  � 0���UUeYUU]UsesU�U�eW��˵{����YWW\V\g���s[s���ưű1�1�,�oqm_kW[gkWm��\Up�qVpe\U���U�]���}���]�U��������������������    ��������������������߯_�WVUUVeUVUUUU�UVUUYUUUUeUUYUU�_U�%�	(
��@(P
@@       � L�_�Z��]�CU�Y�UU�UUUYYUUUVWU\U\YpUq]_sUs���ƶ�����s�s��m�mƭ�������ư���\WUY�U{U��{�{��UU��u�u���w�UU��������������������    ���������Z���]Z���Z�������������U�UUVVUUe�UUUYYUUUY�UV_U�W@}P��5��(�	TP@(P_�0�0�?�jU�f@�d  �g�UUUYe�UVUUVU�V�Uuuu�m�m���V\ss���ư�����qU_YUUU�YVWUWUU�e�V���������UU_WuW_WuWWUU��������������������    ��������������v�گj�����z�n�^�W�U{e]UUU�eUU�UUUUUeYUUe�UUUU�����������?���e^UpUЙ�U[W]@^��dW�U�W W�U�epUpU�eWW��\�p�qm�m�wqܟ\UpUq��U�Y��p�_�UUe�UUYeUUWVW�g�V�U��ݫ߭׵׵׽׷׷׷׷�������������UUu�uWu}u�uUU��������������������    ��������������������~�WU�YYUUU�YUUU��UV�U{e�V�����틭����������������ժ�j��e�U�U�U�Y�U�U�٫U�U�Y�U�Y�U�e�U�V^e�U]e�U�U�Y�U�e�չ߹z�j�o�u�ͭͭ˭˫ʫʫʫʪʪ�����j�֫~��������������������UU]�]]]]]��]UU��������������������    �������������������������U�V�կ5�-�+�)�)�髹���������������������������ww��                ����������Z���]��}�֪j������������ � � � �     ������?���     �Z���]W���V�������������������UUu�����w�w�UU��������������������    ��������������������������������������������������������������������������������������������������������������������������]���Z���������������U�_�u�u�u�_�U�����ꪪ����������          � WW:W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W���UUUUUUUUUUUUUUUU��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ����� ����� ��� �0�[�I��H�H�F�I�G�0�`��� ���H�H�0�0��� �P�P���)�� �� r� ��LE�` �')�
��R�I��H�� �HI��H��
�� �����`�')���') JJJJJi�� ��`�')��'JJJJ��8���\��� ��� �P`����������������&   �� � ������ �� a����& ��� ���P���)��)������ ���)���)?�?��v0 Q�� �P�ʩ������ �������`�K�G�[�F�v�� ��`�K�I�I�H� �u�I�G�H�F�u���0�� ���H�H�uLm��	�v Q�`���쁅I��H�܁�(�䁅)�
�����F����G� �F�H��(�� ���Fe(�F��G�)��`
((

FOORBBOO��ZZ�̃ԅ܇��؈T�|� �? ?�� ���?   ��������? �����gWW/"�  ��GtDWU���������W�U���  0  1WU�������ff�UUU-"�    LtDWU���:���Ù��UUU���    WU��:����ff�UUU-��  � pL�U�?��:�� �ٛ�UUU��� 00�UU5�:�:�: �6l�UWW-"" pL�UU5���:�:��9�yUWW��� 0�UU5���:�:�~6lvUWW3"" 0pL4WU5����:��ٛyUWW��� � 01W�?�����~ffvUWW3""   LD4WUժ�� ������yUWW���   WUժ�����n�g�UWW3"" 0  sDWUժު����9��U�U��� ��0WUժ^�: ���?�?�����  �����?�_�?  �           _          �u5          ��5          �u�          ���          ���          ���          ���   <     ����  �    ���� ��    ����� ��   �����  ��   ����� ��?   ����� ���   ����� ���   �����? ��<  ������ � 0   ������� �   �������  �������3   ��������  �����  \W������  \������  � \�������0 � \���������� p���������� p����������? �����������? �����������  ����������?  ����������?  ����������?  ����������� ��������?   ��������   �������    ? ���?�        ��                  �           W�          _�          ���          ���         ���          ��?          ���    ?    �������   �����?���    �����? ��   ����� ��   ��������?   �����?����   �����?����  0����� ���   �������<?   �������? �   ���������   �������<�   ���������  ����� �\W������ �\�������  � \����������� \����������� p����������� p����������? �����������? �����������  ����������?  ����������?  ����������? �����������  ��������?   ��������   ��������    ?  ���?0        ��    �?�?���?�?�?��?�? �<<� �<<�? �<<�� �<�?���<����<�� ?��?�� ?��?��?�<?���<<�����0000��00����������              00���?  0�  }? L�� �0�t�}]��q �q�:� �5 p  p   �  < ���p<0�S�� �>� �s1 ��1 ��1���1�5�p5 p  ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � Ð���& � �P�P���)���P�����&  ^����& ���� ��`�W�I�V�H ���P�R� �<�Hȩ �H�����<�H ���R�� � �� Ñ ��`����R���	�
8�	���RL���H�G� JJi��F ���R��H�G� JJi��F ��� �R�R����T� JJ}���U��T����a���S�U�H�T�I � ���S���R�R��ȩT�T� JJi}�U� �R�R����� �����a�T�I�U�H � ���R�R���`OR�=/ .12�Ui�U��T`���*�J�I� JJi��H� ��� ����H�Ď�� ��晥����`��������� ���N�I� JJiM�H������I�G�H�F ���H�H晥���� ����������I� JJ}���H������������I�G�H�F ���H�H�ƛ��晥���ƥI�G�H�F� ���������
�
8�
���Lx������ �� �� �åI�G�H�F���� ��`HJL��m 
 � ��H���� ����R� ���Hȩ��H�����?�H ���R��`��R� ���Hȩ��H�����?�H ���R�� ��H����`�G�W�I� JJi��V�H� �F��G�V�R��S�I�T�H�U� �H�F �� ��S��T�I�U�H ���R��`� �F��G�V�R�W�I�V�H��S�I�T�H�U� �F�H �� ��S��T�I�U�H ���R��`��������������������������������������������������������������������������������������������������                                                                                                      �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������(�L�p�����ܚ �$�H�l�����؛��h��� �D���Ԝ���@�d������<�Н��`�����̞��8�\�ȟ쟀����4�X�|���Ġ��x���0�T�����,�P�t�����(�L���p�����ܣ �$�H�l�ؤ������ �D�h�����ԥ�������@�d�Ц���<�`�����̧8�\�������Ȩ��4�X�|�����ĩ0�T�x�������,�����P�t���(�L�p���p���p���p�����ܬ �$�H�l����� �D�ح��h�����Ԯ���@�d�Я�������<�`�����̰��̰��̰��̰��8�\�����ȱ�X�|��4���Ĳ��0�T�x����,����P�t�������(�L���ܵp��� �$�H�l�����ض��h��� �D���Է���@�d������<�и��`�����̹ � �UpU5pU��u��u��u�WU�WU5WU5\U�� � �U\U\U5wW5wW�wW�WU�\U5\U5�U � � �UpU5pU�\��\��W��WU5WU5WU\U��  � �U\U\U5W�=W��W��WU�\U5\U5�U �    � �U\U5WU�WU�WU�WU�\U5\U5pU�� � �U\U5WU�WU�WU�\U5\U5\U5pU�U �     � �U\U5WU�W��W��W��\U5\U5pU�� � �U\U5WU�W��W��\�5\U5\U5pU�U �     � ���<0�<�<�<����\U5\U5pU�� � ��<?<7�����\U=�� < � p��U �  � �U\U5WU�\�5�7     ��\}5�U � ��p}\U5\�5�       � \�5\U5p}��   ��0W�\7�\=W����\U?pU5������?��0W�\5�\5w=�u=\u=p��� �  � �� ��p�\57\5?|�0|]?|]5�W�� ?  � �   ��p��57|5?W�0W]?�W5\U��?���?   ��pU\�5\7|37��5|U5pU��?����    ��pU\5��5��=\�\U=pU����? ��   ��pU\U5\U5|U5�U5|U5pU��?����    ��pU\U5\U5\U=\U�\U=pU����? ����p��<7�<7� 7\�5W}�wU�|U=����?�����0  0<0<0< <���wU�|U=����?   ��0  0 0<0<0 � �0 ����?���   < <� 30���      ��0�� 3< <   <<<���WU���5�<7�<����\U5��5WU����<<<���\U�\U���7�<7���\U���5W_5���<?<<<���WU���5<�77�����\U5��5WU����<<<���\U�\U���?�<?\��\U���5W_5���<?<<<���WU���?<<<������\U5��5WU����<<<���\U����7007??���\U���5W_5���<?<<<���WU�\U5\U5WU�WU�\U5\U5WU����<<<���\U�\U�WU5WU5\U�\U�WU5WU5���<?���\_����7<<7<<���\_�WU5WU5���<?   <<<��7pUp�\�5\U5p}p}��7<<<         �� p]pU�� pUp]��             3  3  3 � ��00 � 3  3  3    � �]p�\?0\?0�< �7�W�U �  � ��     � �]p�\?<\?<\�7�W5_U�U���?�  � �u���5�5<p?�� p��U �  �  �    � �u��<�5<�5�5\�?U��U���?�     � �]p]��0��0��?\U5|�?��?��? �    � �u�u�333��?\U5��=�W?��?�     � �UpU\U5\U5\U5\U5|U?��?��? �    � �UpU\U5\U5\U5\U5�U=�W?��?�     � �UpU��?�<3��?\�5|�=�U?��?���    � �<0��0<<<��7\}5|�=�}?��?���   � ?W��W��� �<<< � <<<� �W��W��� ?   < <� 7�   ��3  0 �0� 7< <   �� \UWUWUWU5wW5WU7W���_�\U�pU5����pU5�]��]��]�W��W5�_5�W5WU5\U���� \UWUWuWu7Wu7W]5W��\U�\U�pU5����pU5\��\��W��W]�W�5WU?WU5WU5\U����pU\U5\�5\�5\�5wU�wU��U�W��\U5��   ��pU\U5\�5\�5W��wU����\�5\U5����pU\U5\U5\U5\U5WU�WU�WU�WU�\U5��   ��pU\U5\U5\U5WU�WU�WU�\U5\U5����pU\_5��7<0<<�<7�����W_�WU���7����pU\_5��7<0<�� ����WU�W}�\}5�� � �U\U5�U? �        � �U?\U5�U � ��\}5���< < <  �  �  < < <���\}5���� \UWU�UWu�w5\�5\�5|Upu5\������ \U�U�UWu�w7�_7_]7w�5��5p���?< ��U5pU�pU�p]�\]�\W5\W5�U=\]W_5��? ��U5pU�pU�p]�������u�\_�\W7�W<���pU\�5\�5\U5w���U�\W=�Up�?��?  ��pU\�5\�5\U5W��w}�|U7�U���?�  ��p]\]5\W5\W5wW��U�\W=�Up�?��?  ��pu\u5\u5\�5W��wU�|�5�U���?�  ��0<��3<0�0�U�WU�W����7��7\}5�����0<��3�0�U�W}�W����7��7\}5\�5� ��0< ��0<00������7�?<��0p}��   < <� 7�  <  �  �  < � � 7< <   �� ����:��:����:��:����pw��<3�� ����:��:����:��:����pwpw�� �� ����:��:����:��:����pw��<3�� ����:��:����:��:����pwpw�� �� ����:��:����:��:����pw�} � �� ����:��:����:��:����pwp� �0 �� ����:��:����:��:����pw�} � �� ����:��:����:��:����pwp� �0 �� ����:; ;<; ;��:����pw��<3����:��:< 0< ��:��:��p��<3< ��:��:<?�� 00�� <?��:��:<           <  � � �0 �  <           ? �� pWpW\W\U\U�_pUpU��  ?  �  W�]�]p]5pU5p}5�W5pUpU�� ?  ? �� pupu\u\U\U\�pUpU��  ?  �  W�U��p�5p�5pU5p�p�pU�U �  ? �� pWpw\u\U��\wp]pU��  ?  �  W����p]5pU5pW5p�5pupU�� ?  ? �� pUpU\U\U\U\UpUpU��  ?  �  W�U�UpU5pU5pU5pU5pUpU�� ?  ? �� 0?03<?��\w\Up]p]��  ?  3 �� 0303<3��\s\spsps��  3       0 0 < ������0 0                   0 ����0              ��� p�<\]�\��wW�wW�w��W�=\�pU��  ��� p�\}\U5W]5ww7ww7Wu7\u7p����?  �<_�U5WW5w��w��w��|W�pW5�U ��?  ��_p}5\U5\U��������]��]5pW��  7<77����wU�\w�\w�\w=\U\UpU��  0 <�0���WW��U�w�5w�5|�5pU5pU5�U �  7<77����wU�\��\��\��\U7\UpU��  0 <�0���WW�wU�wW5wW5wW5�U5pU5�U � < �07���U����|3��3�=0��?\U5p}�� <  � ��T��� 3�3�00<�0U@}�� <  � � �7 � 0� 0 0  T  }�� <  �       � 0 0       |  � � �UE5 ��0�E�\U5pw��   pw��  � �UE5�0��0�E�\U5pw�� pw��     � �U\E1W�W1�WE�\U5p��3   �� � � �U\E1W1�W1�WE�\U5�� w�� �    ? ��\D 535 5\Dpw��    pw��  ? ��\D353535\Dpw�� pw��     ? ��\UWU5WU5W5������    pw��  ? ��\UWU5WU5W5������ pw��     ? ��\D353535\D   �� pw��     ? ��\D3535            pw��       ��\@5 5�0   �    pL��       ��  4 4        0       �� T�P5�P5�pUsu5�5WU�W����5 ��� T�P5�P7tpupu7p�5�U �����  ��0\�\�p4�U\]�\W��U�W��\?� ��|0W�w�\W4|WwW�W|U�� �U��<�<�U�\5�4��W4�wU=UpU=|}�W�?� <�<�U�\5 4��W�|U�pU�|UW}=�s� �?<�<�U�\U5\U5W��W]�w]?�pU=|}�W�?� <�<�U�\U5\U5W_��u��u�p_�|UW}=�s� �?<�<�U�\5�4��W4�U�p�p�|U=W}���?�L0��W4�U�p�0LD1��           D�31@�0                           �            � ��0��:�U��U��U��U��:0��� �  � �~����5� �� �� �� ׬�5���~ �  � �=p�\�0ת�ת�ת�ת�\�0p��= �  � �� ��2�T����E����80��� �  � �� � 0 �� �� � �0 � �� �  �  �       � � � �      �  � �? 0� L�ӝc�1h0ԃţA�lP0�� ��ap8pw:\w�l��h�ԃţA�lP0���? 0� T���cd1h0ԃţA�lP0�� ��d09pv7�t�l��h�ԃţA�lP0����p�a0L�1L�5�Aţ@�+P���L6��   ��p�i0LU5L�5lU1+Q���L2����p��0(0
4�ţ@�+P���L6��   ��p�(0
4�5�@1+P���L2����p�a0L�1L�5�Aţ@�+|�<�=�      ��p�a0L�1L�5�Aţ@�               ��p�a0L�1                        ��p�                              ��pU_W\W5_U5�]=_=w=�7�U�W�?����pU_W_W5pU5�]=_7_7�5�_�pU?�� ��pUp��\�5\U�\u|�0|�0��0WU?�������pU\��\��\U|u��0��0\�0W��U ���pU\�5\}5\�5�<�� �7 ?���\��W= � ��p�\�5\}5\�5�<�� �� �W���= |� ����pU\U5\U5\U5WU�wU�wW?������W � ��pU\U5\U5\U5WU��U��u�W����= |� ����pU\�5\�5�}�W}����< <� 7\�5W}������pU\�5\�5�}�W}����< <� 7L�1�����pU\�5\�5013DL�              3@D1L�                        �� <?�<������5U�W�|U=pU\]5���< ?��<7�7�7���5|U=W�]�\U5\]5\�5��?��<7�7?�7���5|�=����}���7\]5\s5��?   ��?������� ?             ��?������                  �� 00?�� ����             0��� wuw]5�W3���\�w5|��? �� �� 0��� wuw]5�W���3\�w5|��:�<��� W7�]�\u���7_7��5�\�7�W= �3 � ��� W7�]�\u���7_7��5�\�7�W=������<<?��5\ww]7��5<7?7��5\w���� �<?��5\ww]7��5<7?7��5\w�����  <?��5\ww]7��5��Ww5��7\]���� �<?��5\ww]7��5��Ww5��7\]�����  <?��5\w��777<?77��7\w����   <?��1Lw7?777<3777?7Lw����   <?��0@777 7<07 77@7�� ��   0? �    4 7<  7 4  � ��    ��?\U��U�<W=���:W�:��;p��� ��� ��?\U��U�<W=���W���>{5��?;<�   ��WU5WU|�<��0�^��~���?0W0���  ���WU5WU|�<��0�z��zռ�?�\����0<    < ��p}\�5\�5w�=�U7���W3��3� �  < ��p}\�5\�5|���U�|�?s�:��:��  < ��pU\}5\�5w�=׾7���W3��3� �  < ��pU\}5\�5|��ܾ�|�?s�:��:��  < ��p}\�5�<7�<��������U3��3����  ��pM\�5�7��   ����E3��3����   � p \ 5� 7         � 3� 3� �       0  4                00     � ���:+��'�����{U�\U5p��� ��� � ���:K��K�����{U�_U�\U5�U����: � ���?��������{U�\U5p���� �� � ���?��������{U�_U�\U5�U����: � ���;{"�{"����{U�\U5\�?����?�  � ���;�a�a����{U�\U5�W5��?��� �? � ���:��ꫪ����{U�\U5\�?����?�  � ���:��ꫪ����{U�\U5�W5��?��� �? � ���;{"�{"����{U�\U5\U5��?�����?    � ������:��:�U?pUpU����:��    � ������:��:� ?      ����:��    � ������:            ����:��0 � ;� ;� ۖ�WU3�L=�4p�5ph�� ?  � ��j3�U�lU�s3�_314��\hp� � 0 � ;� ;� ۖ�WU3\�=�4p�5ph�� ?  � ��j3�U�lU�s0�_034��5\hp��?  <  � �Õ��U��U�gE��4D4\P���?  0  �  ��3W>�U�g���4D8\ �R � <  � �Õ��U��U�gE�E4D4\P���?  0  �  ��3W>�U�gE�E4D8\ �R � <  � �Õ��U����7?���7L4\\���?  0  �  � <� ���V7p�D�� ?          0 07 � �p��� �4                           7 � �  7    0    �?p�;\�:ܵ�uW_0W�\�0\Up� �?     ?��\�W��u�W]�W�\5�\55p��?       0��W�W5p]7p]���p�_5�U5 W �   �� �WpW53]�o\�y�Gv5�\5�W �    ����U�wU�wU�|�=|U=�U�s]�|]=�U �    �0�U3wU�w��|�=|U=�U�|U=p}�U �  ����U�wU�wU�|U=|U=�U�s_�|U=�U �    �0�U3wU�wU�|U=|U=�U�|_=pU�U �  ����U�w��w��|�=|}=��óiμ�>�� �    �0�U3w���}�|�=p}���i���U �     � �Up��}p�pU�}p}p}�} �       0 4      �       040    pU���߳�5�������밪:�� � � � �Up��ܪߴ�5�������밪:������� <pU���߷�5�������밮:�� � � � �Up��ܪߴ�5�������밮:�����?� |U5���p�������꬯?��:�� � �  ��W|�7ܫ�p�������꬯���:������� <|U5���p�������꬯?��:�� � �  ��U|�7ܫ�p�{�����꬯?��:�����?� ��<����޼����ꬪꬪꬪ갪:�>��?�?��<�����ܺ���껪껪꼪��?�?��?  ?0�00�3��޼����ꬪꬪꬪ갪:�>��?�??0��<��7��7��>�������  ��<����޼������ꬪ����:�>��?�?��<|��{������뻺뻪����?�?��?  ?��<����޼����묪ꬪ��갫;�>��?�?�0�=<��7��7�����>�������  � ��?���ì����אַ���7�������  �� ;��>��ì�ì�>��ﯮ���7���<��   � ?? �� �� � �        � � �� �? �� ?      0��    ��   �� 0         ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  � ��� �'�R��S s�������& � �P�P���)��'�)@�� � `��R�R��� �R��')� s�L��R


eR���X`�R����I���H� �a �`�R����I���H�S�a ȥSI�S`HKNQT� �R�S�R���I���H�I�G�H�F�S� �0�� ���H�H�SL���S�R�R��ͩ �R� �S�R���I��H�S� ���I�G�H�F ���H�H�S�S���R����I�G�H�F ���R�R���`ILORUDX[�
 � � ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������$
�����6����7�Q��8�R��9� �:�@�;���0��1��2� �6�3 w��:�>�;�? ���6��7�:i�:��;�2���2�:iX�:��;�;�0�0��о�1�1��ж`�3JJJJe9�=�3)



e8�<��=`� �������<�>�>��?�����>i.�>��?����`��                                             '0:LWaml �       (1;MXbn|���      )2<NYco}����    !*3=OZdp~����    	"+4>P[eq����    
#,5?Q\fr�����  $-6@R]gs�����  %.7AS^ht�����  &/8BT_iuI�����            jvJ�����            kw�����              x�����              y�����                        ���CC�����9{V�GF    ��Ϡ���U�Kz`�HED                                          S�                           � � � 0�000000000�� �   �                    ��    ?�� ����?�    ��                       � � � l l [ [�V�V�U�U�V�UlV��lf���j�f���� � �                ��    000000�    ��                         � � k�V�UlU[UVUVUUUUUUUUUUU�VUV�i��e���e���j����������������� � � �        ��    �?��� � � � ���?    ��               � ��k��o=�5 5 5 � � U�U�U5UU5U5U�U�U�U�U����f��nf��zf��zf��f��f��f��������      ��     �         �    ��                           ��V��5����� � �                   � ? :   ;�;�;g��g���z������g���g������      ��    <�    ��                     ��??@@DDU��5�7p7�0 ? �         � � � � ���<� �    ��9f��f���f���f���f��f晹f�������      ��    0 0 0 0 3 < 0 0     ��                  ��?  DUUUUUUUWU�U�����������_���7�5�5}5W5_5�:�;������pf��of��~f��f��f��f���g��������      ��    ���� � � � � ��    ��          �?�?�?                ��  DDTU��<00        � ��� � � � �        < � � � ���������������~晙ff��f晽������      ��    �3 00000�0 3��    ��              ��?<<�?�?? ? ? <         ?�?�? ?         ? ? ? ? ? ? ? ?  ? � ���??�?�  �?�?�?        �s s             �?�?�?�?�              ��  DDUU_�p�� 0 0          �0          �   ; ;;;�����n���n���g���f��fꙪg������      ��     � 0 0   � ?    ��          ��?�?�        ?�?�?�?�?�?�?�?�      ��  DDUUU�W?_?_?_?|?|�|�|?|?_?�?�?�?�?����|=�?�?�?�?�?�?����ff��ffٟ�z��ff��ff���g���g������      ��    030�?00    �     �  ? ? ? ?               ��  DDQUU�W �        � p p p �          � p p p �       �����z�����������z��z���z�ꫪ����      ��    �?��� � � � ���?    ��   0 �              � W � � p p �                 ��        � �D UUUU�} �       �  � �      � �   ���f���f���f晙ff��ff��fg��f{�꿪����      ? �       � ?    ������\������������������������������W �                   � p \ � �  �?�?�?        ? ? ? ? ������? UUUUUWUW�\?�?�?�/�/���?����������� �n���g��f���f���f���f��f��z������             � �0<<�<33�   � � �        �?�?�?  ? � ���������_k���p� � � p � � � W�}_֕j��������???�?�?�        �?�?�?   �?�?�*? ���U�UUWU|U�W �     � � � p � � ���� � � �����of��zf��n枹n���g���ff��ff������           ����|}�}�Q�P    � � � � � � �  �0?<�?�        �_~UW��     W ~U�_��������Z�������������:�                                     > ��U�U�UUWUWUWUUUUUUUUUUUVUZU[U[UZUVUjU�Z�kf���f���n��n��f���f����������?           ?���W��          ��?<?�� <<�?�        � u�_UP@�P�}�u������Ɦ������^�^�W�����W�����               > � �UU9U�U�U�UUUUUUUUUUUUUU�V�UzU~U{UnU������꿪����Ϊ�� :                   = �P@5 � U T � � � � � �@�@�@�P�P�P��\�\�G�A�P�U���������������Zo�֭�k�ꪪ����� 9 9 � � ��UUUU9U9Y:�9f:�f���                            � � � � � � � ���p�p�p�p�s����^��<7�7�7<��^?� � � � :                       : � ���:�:�?�_]:�:�:�5���:�:�:�:\9�                             ���                � ������ � ��?�?�?�?�????????����? ?             �?�?  ? � �� ? ?�?�        �?�?����������        ��<<<<<<�?�?<<        ��?<<<�?���?<       � | W���up]p]   � U_uU5U5�u�� W | �      u_U�            ����������        ��p�3�����|�?��ŕ��K��ј��W��ݛ��c�&�鞬�o�2�����{�>��ĥ��J��Ш��V��ܫ��b�%�讫�n�1�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ��j�ֲB�����?���kYꛪ雪�Z�k�ꫩ�����������?��?0S]�_��1L��S���S߷S�_S���700   ���/�2<����0:2<� ���0   ���[U�������������ۗ��[U��������������UݗUٗU���We�We�We���U��U����   <�2,� *"   (�(�/��
   <�3 �    ��?������y�����竧߫���w�������������UT9�:Ge�G��Wf�W��Wfꗩ�\�:�� � ���:�:������< ���������;����WUէ������3����'�ۧ��WU����������������A�{��$�I�C�ۓ�����Ɠ��������3����{��0��� ?�� ���0�Ǽ�6�����WU�����(�7��7(����WU����WUի������|7S������3��w~5{�۝{���6m�7]���<  � <<<3�<  0������� � ��0� <�   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �H�@�I�/� �H�� �����`��K -��K�K� ��� �K� �J��J��������` R��@JJeH�H��I`�AH)��o��HhJJJJ)���y���I` 0`��� P���@p��@@@@@@AAAAABBBBB 	�Hi0�H��I`�I�  ��  �`�Fi0�F��G`��



���� ����F����� ������`�\�5�5�5�5\��|\|ppp��\W5�5|WW5��W5�5���5W5�0����=W5�=��W5�W|5�5W��\5W��5�5\��?W5�5�ppp��W5�5���5W5��\�5�5�5|5W�      �?�?       < � ��� <  ��?<< �  ��  ����� 0   <<0        ��H



����h��� �F����� ������`� �ÑF����� ������`��<<<�?�?<��?<��?<�?���?<  <�?���?<<<<�?��?�? �� �?�?�?�? ��   ��? ��?<�?�<<<�?�?<<<���������?�?������ ?��� � ��?< < < < < < �?�?<??�?�?�<�<�<�<<?<�<�<�?�??<��?<<<<�?���?<�?�   ��?<<�?��?�<��?<�?���?�?� ��? <�?��?�?������<<<<<<�?�<<<<<<���<�<�<�<�?�???<0<??���??<<??��� � � � ��? ?��� �?�                 ����   � �         �0�        �?�?      �H�H��I`�H�H����I`�H8�0�H��I`�F�F��G`�������� � � �* �	�
`�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`�ð9� �I� 	�H�a
���ӅF��ӅG��b� �F�H���� ���Fi�F��G�b��`�P� O� X� �� a� �ͩ �P`���'�')�Y��Z�Y��0
�a���`  ��Y�Y�Y�Y�Z��`���<� ����� ��ɀ�%�@� �ʦ�� ���@��� �L��  �L�� u�桥����`���P�Q���L��
�G�p�p)š�;�� �3 �ɦ�� ��
�0����
� �(
���H
�h
��
��
�� ��
`���`�`��J� �` �� e� �� �˦����
��)I���@

}���uɅG��ɅF �ߦ����������`�����������������8\����4X|�������(� �)�(��
8��(�)L�ɥ(� �)�0`� �𦡼@��
� ����
��0�����yШ� ���`  ���0��𦡽 ŀ�#�@���0Ł�����@ �ɥ�������@`������� �ɥ��0���,���0Ł�#�@��� ŀ�� ���@ �ɥ�������@`���P�W �ɦ�������� #� �ɥ��=�����`��������ʐ'� ������@

��������ʝ@ �ɥ���Ƥ��`���P�P��� �P�@�yН ��`    ���� ɀ���	@� � �`����}p˅� ��`���`���`�fː6� �` �� e� �˦����@
yk�}�����G���F �ߦ���I��`  ���`��)�'��JJJJJ)����)����e�����G���F �� �ߦ��`�`�p�
���  ��Ơ`  �˩ �a �`���� �I� 	�H�P��@� �È��`�� �È��`��  �  �  �  Ĉ��` �� �� �� �����`�) �[��ŋ�U������z�����}Ш� �<����� �@
�`
��
��
�� 
����
��� �e���
� � 
�揥�)����`�)�(���$��� �������)ŏ����
����
� � 
`���D��� 0=�-�9� ����ł�$��8�-��������  �̥��`� �a  �Ɨ`�����`�������Ո�����	��i����� ��`c
��ɸ�ƈ����` �� �Щ��& `摥�)��$����JJJJ}lͨ�oͅa��� I� �`���`  �`  &'&'&'&'))( *+*+*+*+))( ��� "�`�)��	�r����`�r��r�r�����s`������
���r�� P� � � �̦�����Ͱ愥�� l� ��` '�`� �� 	Υ��������͐� ����� 	�`��)�
���;� ���2�)�����)���� �)�
��������)�������� Q�`����}Ш� �� ���z�y���`���`��
���y���yݗΐ� �y�z�z)e𪽙΅a  �` "$��� �I� 	�H�z� ����� �a �`������&�����z�υ `���z�υ `�	��z�υ `�����z�υ `���z�!υ `��ɦz�$υ ` �y���y�Oϐ �� �� IХ�

ez��Qυa � ��` !#$%"���;���8�z)�1��� �I� 	�H���
�z� ������ �HI��H���� �����Ɔ`������ ɀ�����!���褂� ���ߢ � �@��ł��������� P�`����`� �y�z�z��� ������}Ѕ��й� }Й� `  ������� ��`�� ��`��  �  �  �  �` �� �� �� ��`��� �I� 	�H�z ���`� ������	�
8�	����LfЦ��ЅG��ЅF� ��� �����


��F��ȱF����ƚ������

��F��ȱF����ƚ��晥���à� ������Й������`0Tx������ `� ����&  �ҩ � ��������������s�����z�y�����r���������`�������� ��
��
��
�@
�`
�ĝ 
�� � ��� � �a�`  ���Ð� ��`� � � ���� ȩ�� ��Ðꈄ}�����& � �P *ҥP����� �ѩ��&  ��`� �{���|� �~���{i�{��|���~�{�	� ������~�~��� ����������`�
����~� �P�P�� ��ƙ��`�#�����}�8�}��L�Ѧ�� �~� ���}� � �}�#i�#`�#�����}�8�}��L.Ҧ#�} ���e#�#���}�8�}��LHҦ���� ��� � ��� `�@�I� �H����H��`���`�H��� ���H ������@�I���H��� ���H ������]�I���H� ���H��`��`�������	�
8�	����L�ҥ�� P�`���& � �0��A��@��1 A��0�H� 	�I� �0�@i�@�1��Ai�A�0�Ð�` �� rө��& �
��S��B�T��C� �0�0�`�B� �a  ��0�0�Ð� kҩ��&  ^� ^� Y� O� ���������������`� �ݘӐ����
�����F����G� �F� ��l��`	$.�$H ���%�I�mՑյ�����!�E�i֍ֱ֕Թ������A�e׉׭������=�a؅ة������9�]ف٥������5ڡ�Y�}����1���                                    ������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������@�¤�8(�,�����������������/��@�   @�2�4�"8�*<�?��?��/����@�   �����U�Q�ZA�U T UZA��E��U����       ������[UU[UU������             0� �?�j�UU�UU՚j��?0�        � ���������U�������U�����������U�������U������ �       0 ������UUUUUU������0       �������U�����������U����lQ9kE�ZQ�ATU U@DUT UZD�kQ�lE9��Ϭ�����kfe[UUKDD[UUkfe�������������:��9Vf�UU��DD�UU�Vf險9��:������>�a�[E�kQ�E:kQ�E:kQ�[E�kQ�E:kQ�E:kQ�[E�kQ�E:kQ�E:kQ�e꼪>����ϫ�����VfeUUUDDDUUUVfe���������kQ�E:kQ�[E�kQ�E:kQ�E:kQ�[E�kQ�E:ë}�8�"ër�������*��
����/��@�   ̫0�	̫��,�*=�*?��/���@�    ���U�p�5���ܵ�\�����pU5�U � � �     ���U�p�5���ܵ�\�����pU5�U����� < ���U�p�5\��ܷ�\�����pU5�U � � �     ���U�p�5���ܵ�\�����pU5�U���?� <��Wp]7�_��z��z�\_=pU5�U � �  �   <��Wp]7�_��z��z�\_�pU5�U����� <<��Wp]5�_��z��z�\_?pU5�U � �  �   <��Wp]7�_��z��z�\_=pU5�U���?�  �<���U�|U�\U�\U�\U�\U�pU5�U=��?�? �<���U��U�{U�{U�{U�|U��U?�W?��?  ?0 00�3�U�|U�\U�\U�\U�\U�pU5�U=��?�? 0��<wU7_U7WU�WU�WU�WU=�U�����   �<���U�|��\��\���U�\��p�5�U=��?�? �<���W��u�{u�{u�{W�|���U?�W?��?  ? �<���U�|U�\��\U��U�\��pU5�U=��?�? 0�?<w�7�]7�]��]�w���=�U�����     �  � ? ?�������?��?������?��<�   <  <???����?��������?���?��<�      0��    ��   �� 0         � ?? �� �� � �        � � �� �? �� ?�� 7|�=p}�\U�\�=\��_���7�U�<��   � ��?p��\u�\��\��\���7�U�����   �<�����|���U�\��\w�\w�pW7��=��?�?   ��?�^5��?�0�0�0� 0 0 0��?    0 ��*��*�+8+8,0Q0U0�/��*      ��.� /8�,8�,<�<< <8<,� +��+��/      ��*�(*��"��+8Y,L4��?L4L4��?      ��*��80#?<��0��?��?��?��/��+      ��* (��*��* 4��4 44 4��?      ��+<�<}0 0 0< <8 ,8 ,8 ,��+   �n� 
�� 
�`��� ��a  �`��	��� 
��
`��)�쥙JJ����ř�� 
����
��� �� �`�����@
�@
`���� 
��������
� � 
`�� 
`��` �ۥ�������ɀ�	�����@
`���`��� ����Ŋ��܅a  Ȧ����@
`�܅a  �`		

�n����ʊ

��� �����@
2���uܦ��� }���yܐ ��Lcܥ�}�܅��� ��� ��Lc� �ۥ�i ���暥����`  ����������������-��<��K� � 0)@�	��^��Y����`���M� �Y�Z�n�[� 
�\�[�@
��]�\�^�Z�^}Ѕ^ ���]��[i�[�Z�Z��ӦY���!�e�� ��`  
#(-27�n� 
�� 
�`��a  � ��`���0����� 
��
`��)�襙JJ��� 
��� �o o�`�n����ʊ

��� ������}�܅��`���@
�0�����&�`� ����ř��o���� ��L�ݦo��݅a  ȥ�i ���o�暥����``		

�o���`� � ���@
� � ���a  �`i-� �a� ��0����a���`��  ��`�n� 
�
�� 
�`��a  �`��	��� 
��
`��)�쥙J���8噅�� 
����o o�`�n� 
�
�� 
�`� �a�   �`���
�� �* �
�n� ��
��� 
���Ƈ`��)�ץ�J���8噅�� 
�� ��`�n����ʊ

��� �����@
ř�����}�܅`�� �a�   ȥ�i ���暥����`��n�n��
�2��
0-��
�o� 
)�� 
)��o�oi�a� 
�İ
�`  Ȧn� 
�n�`�
�� �` ߩ �n�n��
�T�����L�')�N� 
��:����
� � 
�3ɀ�	 F� U�L��Ɂ�	 F� .�L��ɂ�	 F� ,�L��Ƀ� nަn� 
�n�n���`�� �F�H���� ���Fi�F��G���`����
�
8�
����L�������X����c�戥Xi�X�
�8�
�X`��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������Ð%�
����F���G�#)��F��#ee'�#�#L2�(� �)�(��
8��(�)L8⦙�(� �)�0ƙ�`���& �#)
����F���G�
����H���I������F����H�)�@� �P����)�`�p)��ƙԩ��`��3�G�[�o������������#�7�K�_�s�������������'�;�O�c�w������������+�?�S�g�{�
&*?FJZz|��������� 
"%)>G�Z���������	!$=EJdxz������� 
#*7IZ^cw��������&5DIMe���������� 	/7;W\ex���������	$+/?EWwx|������
 '*;@HZ\dy������	+35@FIMY[d������	
!7@Ubz|������� $'>E�Z\e}������ �)5?H\ez����� #$)>FKU]d������� "'K<GYegqxy������'(9G[k|����������#,FJOY[��������� ?EGYh�������57EGdgx~���������L7;<ACKOSmqw}����&(+,9ABHZux{������� $?HKe}��������� 
<Z��������Jw� *JWcqz��������'	 *BFHMex������� (DZ]ceh���������-;ACD\~������Ziz��(7��*���,;J  -5;MWwy�������� !(-7FU|}~����-<KZix���,;JYhw� ),7Dq�|������� -����&5������	,-ACJ]cxy}������	
(*7@FKOY����� ')59WY[ms������� 
*,5FHU\dx}�����*-EHKfu�������� #,-9EZ[ch{������� GObcdefx��������	7U[e�����������ix/�$%&�b	
Uds,Jh >\��"^b�c��*u�I�-x���@|����'��,J�� Kx/\�1|�$�qF)�fJ�<K��"#
,}������������������#�/�;�G�S�_�k�w��������������������+�7�C�	  
		 		
 	 	
	  			  
		

	 	
	
	
 
		 

	 
  	
	  �
��{�F�|�G���� ���F�
���� ���ƙ�  �`������������������������ �%�*�/�4�9�>�C�H�M�R�W�\�a�f�k�p�u�z������������                            �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������& ������ � � �* �	�
� ����[�� ������& ����� \� ���������i<���`���`���>�]�:��8� ��i0��i ������������i0���i �������  ���a�.�]�*�D �����ȑ���� ��i0��i ������ ��_��a�Ș -��a����`�`���`��K�]�G��8� ��i��i ��i0��i ������������i0���i ������� ���a�0�]�,�D ���ȱ����'��� ��i0��i ���ߩ���a����`�`



}J��K�i ��J��� ��N�e��i ������`� � ��@����������`H)���hJJJJ�
ei@}�` 0`��� P���@p��      

�� �B� � �����`� �/ �P�P� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                  �����ȱ�� � ����0��� �J���� � ��� �* ���`����� �  �ܥ
��3��4�`� � � �� � �����
����`
��3��4��
���ȱ���� ��	�� k�L�� �L�� ��0]���JJJ���� ��	�Bȱ�4�

��4� �)�7� �� �"JJJJ�%�)pJJJJ	�1 �� � ��`� �.�>�����k�L��+��%8�(�%���)�+ �� )�`� �.�% �� )�`�+���(}%�%����)�+ �� )�`�.�� �� �� )�`�+�Ž%8�(�%��")�%L��")�%���ǽ)�+ �� )�`�+� �� )�`� ���)����1��)pJJJJ	�1�

��)�%�48��4��7� �4�7�4� �7� `�4e�4���7�7��ީ�7���4�ҭ �

��)�JJ%	J� `���� �.`
em ������ )�+�JJJJ�(��.`�����e`���ȱ������.�@���*����� �  `��ý
��
��L����ȱ��
�L����ȱ�L��
qm �����ȱ�� �L��0)

�������� �����)� ����� ���� �	�	�Z��M)x�IJJ�����=��9�0 �8���
�� ���� �� L��e�������� ��	�� � �0

��������( ����) �
����* �
�	�
�� �* `M�9�����+�E���]����O����S�=�2��. } � } .	}.	}�0 ���	.	.	T} . !� 	�	}.	}�
\�
\�	}.	}.	}�0  . T  .	T}	�}0  } � � }	�}	�0  } � } �	}�	��0 �  � � �	��	�T
�\
<�	��	}T . !}`   �
� 	� 
\ 	� 
� 	� 
\ 	� 
\ 
� � 
� 
\ 
� (8 
� 
\ � 
� 
� � 
� 
\ � 
� ( 
� � � 
\ 
� � 
< 
� � � 
< 
� 
< � 
< 
� � � 
� X 
� 
\ 
� 
\ 
< � 
� X8 ( � ( �   X � �   ?����	} !}T. } �	�}	�!� �	} !}T. } T	.	�!}   �
\ 
� 	� 
\ 
< � ( � 
\ 
� 	� 
\ � ( 
\8  �����@}�}T.}@�   ��	��}	�}	��	}.��	�	�1}  �
\ 
< 
\ 
� 	� 
� 
\8  1�1��@ .h�hA� K�����h 	h@ 	@ 	10 	@ � h h	}�  	.	@h	}!h �
< 
� 
� 
� 	� 
� 	� � 
< � 
< 
� 	� � 
� 
<  �����2� 
��}@0 � 
��}h0 � 
���� 
���h 	h}�}0 � 	�h�0 � ��@0 h 	h}h} 	}�}� 	����0   c�c��@  	 T� < 	 T� < 	 T�	 T�  P � "<  � !�  	� �@ < 	� �@ < 	� �@	� �@  �	@	.  !} Z	@	.  }  !�!��2!�	� 	� !}	� 	� . !T@ !�	� 	� !}	� 	� . !T@ !.� �  T }T. � �"\	� 	� !}	. 	. T}�!�    �����@T�T�}�}�� T "<  T�T�}�}�� T !�  @�@��@�@ T !�  @�@��@�@!@ !T@T@T}@}@T@ !� ���<�}@}@T}�T}0   U�U�dh�}�h�}�h�< �}�h�}�h�}�h�}@ �<��<��(X �<��<��<�<�� �}�����} � <  <0 ����} � <  0   ���@T T	@ T @	@	T}0 } }	T@ }@T	@T	}�0 � �	�� � <
\<�T  v0 } }	�}	T.}!@ "< 0 @ @	T} � !�`   ��%��!�!T! � �!.!  !�!T! � �!.T 	T.� � � �  ��@ � � � � � �0 �� �!!. � �� �T� � �!.!�AT@   �
� 
 
� 
 
� 	� 
� 
 
� 
 
� 
 
� 	� 
 
� ( 
� � � 
 
� 
 
� ( 
� � ( 
 	� 
 
� 
\ ( � 
\ 
 
� 
 ( 
� 
\ 	� 
� 
 � 
�8   ��o�ho�P o �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xة �& �� ���  �  �  � � ĩ��& � ��$  �� � P𩩍&   ����&  �  ����& �� P�  � � � �Щ��&  �ҩ��& �P�� @ȥ��3�����s���� P𩠍&  ��L_����& �� P�  ���𝩠�& �� P� ����ЙL����& �� P�  �L�H�H�H���  � � � ��  {� ��P�	 ���'��P��#e�#h�h�h(@������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ � �