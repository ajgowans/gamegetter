                                 	                                                4     4      	             5                         	  4     	    4                                      	      6      6        6   7                                7                 4                                  5      6       6       6       6   4     	        7 	        7  	          	     4                                                 4               4                              4                                                   �                            
         
          
                           > 4                    >                      3                    :   
        
        4                                               3                   :                     4              6        6        6                   >         >               4                                            3               >                                                    4                 :  3                      :                       
         4
                  > 4                       4                                                   �       "       "       "     "      "      "     "       "     "      "      "             ?                  "             8"  =    "   ?  "   >  "     "       "   "     "   ;   " =     "     "    8 "       "   >   "     8"       "       "  ?  "      "    ""     "      "      " =   "   ?   "    8"       "     8"  ;    "       "     "" =  "    "     "       "       "" =     "   >  "       "   8  "       "      "      "     "       "   =   "     8"       "       "     "  ;  ? "       "     ? "       "     ""        "       "       "       "     8"       "       "       "       "       "�                                                                      <      6<  =   6             9               @                                =  9                >         5 =          3            !  ; !!<      6<      6<             9            9            59  >             !!!      !!!!!   9           <    3<     <     !              <  @   <               !      !    ;  =                       =  >          9                         <     !<   !!<  3!!!          >        =         4    =                                        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ��  �������  �<<<< �� �?  �<< <� <<<�   �?�<<<<<�? <  �< < � < <�  �<<< �<<<<�  �?<< < <     �<<<<�<<<<�  �<<<<�? ��   � ��  ���  �   �  ��  �  �  �  �  �     � �  �  0 � � � � � 0   �������   �� � � �        �  0<�?�<�<<  ?<�<�<�??  ��  ��     ���3  ��� �  � � �  �� � � � � 0   �  ��   <�<�<�???  �� �  �� � � 0   �? ?��� ? �?                  �?���?      00��00   ��  ��  _U������ �  ,0 ?0 �  �� ��� ��� p�Wp�Wp�Wp}U��U��U ��  �� �*� ��7 ��� ���      ��  ��  _U������ �  ,0 ?0 �  ��  �� ��� ��Wp�W3��W3^UWU�WU��� �*�<��?����� �?  �?  W� ��� ���  �  �� ��� �0 ��� \��W��U�U�U3'\U3<\U�WU�����n��������?�?�?                         ��  ��  _U������ �  ,0 ?0 �  �� ��� ��W��_�U��W�������?<��?  � �� �U5 ��? ��? �
0 �3 �� �0 �� ���U|U5�}5�W5�\U5 \U5 ��?���뼪�ۼ��ڼ�����?<��  �?  �?  W� ��� ��� �����0���2�pW��W��\U\U\UpUpUUp�_����n��k����?�         �� �� |U �� �� � �� ��0 � ��? �����_��UU=�W����UU�UU�UU ��  �� �*7 �� ��? ��?      �  �? �U� ������ : �8 0� � �  ��  ��  �_��_��_���U�0�U�0�U� ��<�����?��� �  �? �U� ������ : �8 0� � �  ��  �� �_��_��_���U}�U��U� ��  /�  �� ܣ �� �� �?  ��  W�  �� �� �  3�  3� � �����5�W���U���U���U���U5��U5<�U�������p�:p�:�?�?��?                         �  �? �U� ������ : �8 0� � �  ��  �_��_��W�V?��>���>���?��/<��  �� \U ��7 ��? � ̀ �� � �� ��� p�U\�U=\�}�\���\U5?\U5 ��? ��?窪>���>��>���? ??< �?  ��  W�  �� ��?���3�Ì3��p��p���p����U�5�U�5�U�5�U��UU�����������������        �� �� pU= ��� ��� 0� 0 ? 0�? ��? ��� ��W|UU�W����UU�UU�UU ��  ?�  ܨ p� �� �����������?��������������������� �� �� �� �� �� �� �� ��������������?����������  � �� �U5 ��? ��? �
0 �3 �� �0 �� �� \ W] _�� wU� �W� W�> WU �� �� �*7 �� ��? ��?  �� �� |U �� �� � �� ��0 � ��� �����_��UU=�W����UU�UU�UU ��  �� �*7 �� ��? ��? ��  �� \U ��7 ��? � ̀ �� � �� ��? p�5 pu� �_� �U� ��� �� �U� ���  ?�  ܨ p� �� ���� �� pU= ��� ��� 0� 0 ? 0�? ��? ��� ��W|UU�W����UU�UU�UU ��  ?�  ܨ p� �� ��     6  �  `  �   7  �  p  �   7                                            (  @!   E   F @@  	  `   @���*WUU ���+     �   p  �	   '   �   p  �   7   �   p   �                         @   P      (   H  Q  ��  � @`   	    ����UU�����                                                                             @U PP� TU� T�� U��@U�*PU�RT��TT�*�U�R�U����Z��A�UZ *  ��  �� ��
 ��* ��� ���Z�����
���*���jj��j������j��Z������      ��  `U �ZQ �VP�VY ` X   X   X   X   � @�VP �UU  ��     ��*�VU�ZUUUY @                         U  U @VUUU�VU����*    �
 �U� UVUPYA	 U %  �  �   �  �@ %P %UYU	�V�*�*        �   �   �  ��  ��  `   �h  	&  �H @� �R `) ��B `$e  ��  h
   )   �   �  i
  �	  �*  f&  ��  ��  �� Y� f� e�
 ��
 e�
  bd `b H�� D�� ��Y Xb� ��� ��� `�� ���  �j   h   `   `   `   �j�
 ��
 e�
 j�
 j�
 ��
 �� i� ��  �*  �
  *   *   *   *   �   �� ���/��������������������������������������������0��?���\￣
��
�� 	���
U�pU�pU�\U��U��
U��
U~�U^}U^MUzO��������A��A��A��A��A��A��A��A��A��A��A��A��U�CU�@�U�@"U�@*U�@
U�BU�BU�H��H��`����@��@��@��C�jO�"HP�"� �N%�T� ?����� ����*<0� ��3 ��>����?� ��?�8*����J?
H%�*�j�N�^/R2�+ �Ϩ����լ*L�3<T/�������������������    UUUU������������p�� ���  ��  \�  p�  p�  ��  ��   � �  �"
 �� ��  ��� �* �   �   ��* "�
 ��
 �� �*( �


�

��
���
��
 *��( ����>����� �
;   , ��� ���  *�   �   *  �*  �  �
            0    00�  �  [��VP���Z @    * � � �h*V ���        0�   �  [ �V��P�Z�  @ � � *  ��D h*P�&�� H��      ���0  �*8�U�:�U�:LUU:�U�:�UU:LUU:�UU:�U�9���:���:���             �?  _��UU�UUp�5p5p5p5p5p5p5p�5�UU�UU _� �?      �� �i��U�6�V�լVU�W�Z�k�j�k�Z�[����\5? \5  \5  W5  W5  W5  �    <� <0�  �  � ���������  �:��: ��� ��� �� ��0� 3� �     �  \  p  p  p  p  p  p  \  W5 ��� ���������     ���* 8�BU9�BU�RUN�R�N�R������~9D�B9T�R9U�R>U�RU�CU�N�����?���?  �SUU�SUU�Se��S��S���S���S���S��S���S���S��������������?�����z������W�__^�]���]���UU��_կ����������������^����������?���UUUU@@TAQUuU]]�U��������������ꮫj��z��ڦ������j�jj�j���� 0  t U�Un����� 0 �t �V�U���� 0  t U�Un�����0 �t �V�U,�²��2�Ϻ��,��.�>(8�
����� ���Z�W�Z�W�n��������?�?������<��<  �  � �/��_-0�U�0�U�<s��s�5 s��?sU_�}��_�0OU U |U; p�; ��: �U ��       �  �? ��00��30_���U���U��s��?s�� s�� sUW]�_u L�; �U; pU� \�� W=����?  ��  0� 0{?0x�0zU�<^U��_W� \W��WW�W�U��}�pW� �U� �U0 �U= �W �W �U ��    �  �?  � �^?^��^U3�WU��WW� WW� _W���U���u� p]� �W1 �U �U �W5�:|����            �  �  ?���V��j=�zU�Z�WU�[�:���:���� �� ������0�jկΪ:�Ϊ��Z��?���ꫪ�ꫪ�ꫪ�:��������� �:  �          �< ���0���3���< ���??�������?��?�?��?����?�������
  ��UU�BU��RU��R���R�Ԓ*Pզ
U�( T�
QU�VUU�ZUVꪪ�����? �? ��������?���?k���k���k���k��������������>���?������ �?  �? �������:���:���꿪�꿪j鿪j���Z���V���V:���:���� �?     00�0 �?��30��������������>������� �?�000000   0  �   �  l  g6 �Y� �]� pVepWupWup]]�]� �u�  w7  �;   ���              � � �W�s5__}=sww3r�u#p]]�]� �u�  w7  �;   ���   � �9 0T� LY� �� ST��$U��D���HY��DU��DV��HU9�DV:�V���� �?             �� ��: ����,���뫪﫪�����ꫪ�묪�찪:���� �                      �� ��: ���0/��?쫪>���:���:���;���<��:<��0��    � ��; ��� �:� �^� �W���W���e���U���Y�������=��U: �� �� ��   � �U��WU?pe�լ�V�|�[�W�5W�5���6�j�5WU���e�ji�UZ���       � ������?���ꬊ��|��Wկ:���:\U�:��:��>�������U=  � ���?VUU�VUU�[j��l��*���:�2�>><��<0��0������ �        ���>��:���:�V�:�]u>�u]�u]�u]��UU���ʬ�����꬯����?��   �?  ��  ��  ��0�V���]u��u]��u]��u]��UU����>�� ��  �  ��  �? �/�l<+��k�:��?���?������迢��+���+�+���/��������������?            ?  ��  7[��\��5[���X�%�  7�  �������  $                                            �  ������:  ��V���� �iU�Z���?��Z�ZU�������U��������V�>�����V��?�����Z����Z���V����Y]�����<�Y]U��>  �U�UU�  pU��U�   _�� ��   W�  _  ��   �  7,   �7  7<   ��  ��   ��      �?   ������ �oj���� <�V��U�: ��U�U�: ����Z�� ����j�� <����j�� �뺪��U� ����j��� ��U�j�� \�V����� \�U���? \��_U�� |���� �� �U��  �5 ���?  �� �:�?   {�    �>     �      �	       `e        Pj)                                           �?       ������ �������?���V�jUiÀ��U�V������U������j��������j��������Z����>�����j�<����Zue  ���Uue  �kUU�U   _U��U   [� �_�  ��  ���  p>   ;�  �   8�  �   <� ��   ??  �      ������?  ����Z�� �jU�V�6< �ZUjU��� �Z������ �V������ �V�����<��U�������Z���^� ��j��UW� �뫪Z�W5 ���VU�_5 ���U��^5 ����z=  ��U? {  �� \  �� �  � ���       �;       �        `       Y	     h�                    �=<�5  ���w�  _U�y  WUU_7 �@P]�  �]u ~�^]U TU]��|UeYU���zYU���VU ��pUW ��pUW �\�W \\�U ��\_U ��_WU ��W_U ��UW� WUU� WUU]� WU��� lUi��  ��V�>  �W��  L~�  0�SU:  ��NU�   S9U�  �U�T�  \UyU�  kZ�i�  �����         <     ���5   �_�  |U�}  \UU_7  U@]�  ��]u ��{]U PU]� �U�YU= �W�YU5 [U�V]5 ���U]5 ����]5 �3�W5 ��WU5�y�^_U5�zUUWU=�]UU_� WUUW� WUU�� WUUY� WV�V� l�Z��  �UU�>  �W��  L~� �S�S�: T�SU: lU�^U: �U�WU: �V>_U9 ���UU:  �ïi:  � ��  <     ���5   �_�  |U�}  \UU_7  U@]�  ��]u ��{]U 8P_Y� �U�YU �W�YU= [U�V]5 ����]5 ����W5 �3�WU5 � �_U5��3sWU=�z�o_U���_W� ��W�� WUU]� �UUY� WZ�V� l�Z�� <�UU�> ǓW�� T^}� [U~_� [U�SU: [U�SU: k��NU9 ��SU: � NU:   �UU:   �j�:    �� �               ?��  3���  ����  𪪪� 쯮�:3 ������ �����>������ ������������3 �����  ����   ��>   ����   ���>   ����   ���>   ����   ���>    ��� ��> 0� ��> �?���� ��ê� �:���? ����i ��i����V�ڕ�.PZ`*�Ze�ր�R媪U*T�Wi�i@U��*�  ��    ���? ���� <���3 ?��? 3��:�����>  ?����  ����  ��3  |���  ����? �����  �����   ���?   ���>   ���    ��>    ���    ��>    ��    ��>    ��>    ���    ��>0 ���>�0���?��i?0���� �pe��l���Օ�.PYZ*�Z��֨�Q�Ue� VUj�U���bUih*  ?            ���           WUU?         �wU]�        p}UU�=        p}Uw]�       \UuU�W       \U��U�=       \]5��U5       �] �}�      �� |wW�      \7  �]w��?    \?  ���w�   �  ���U]��   �   ���wuw�       w���w}�      �_}u}�[=      {��ߟ]��      �uW��m�     ��u����     �߽wu�y�     ������=     ��ߵz�w�6     �{}�����6      ��W����>      ���[���      �^W�> �       ���� �        ��:  �      ���U:  �      _u�U:  �     �WUW�:  �     ���u�  �     ��m��  0     �}�:   0     ����?                               ��           WU=           �U�          �_U           |�5           ���          �uU          �U���        \U]�]�       �_U}uU�      ��|]]w��?    �?��u��w�     ��u��U]��      ���wuw�     ��w���w}�     ��_}u}�[=      {��ߟ]��      �uW��m�     ��u����     �߽wu�y�     ������     ��ߵz�w�6     �{}�����6      ��W����>      ���[��7      �^W�> ;       ���� ;      ����� ;      _u�U: �     �WUW�: �     ���u� �     ��m�� �      �}�: �      ����?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��  �������  �<<<< �� �?  �<< <� <<<�   �?�<<<<<�? <  �< < � < <�  �<<< �<<<<�  �?<< < <     �<<<<�<<<<�  �<<<<�? ��   � ��  ���  �   �  ��  �  �  �  �  �     � �  �  0 � � � � � 0   �������   �� � � �        �  0<�?�<�<<  ?<�<�<�??  ��  ��     ���3  ��� �  � � �  �� � � � � 0   �  ��   <�<�<�???  �� �  �� � � 0   �? ?��� ? �?                  �?���?          ���    d,���%��.`d1d2d3��-��6`d$������������  ����8��������% Xݤ�|� ����� ��������8������  ���������% Xݥ8���������8������ �����% Xݤ�N� ���� �� �����������  ��� �% Xݥi���  �����% Xݥ���� ��� �% Xݥ8���� �����% Xݥ�� �������� ��( 5�`d�T��Z�/���� ���� ��z�`H�
�����轟���h`dd�0����d# ��d� {���%� �R���R�����7���� �d$ Xݩ���%�b���%��R���R���$��7��)��(d&d'��� � \��)I
��R���R�����7��e�� �d$ Xݢ 5������R���R���������n�d$ Xݢ�R���R�����������d$ Xݩ����� ܢ �  ��0 !���
����������d# �ݢ �  ��
 !����񀺩��� �� �ܩ
��d����(�d# �ݩ��%d ҅������� ܭ  ���婁�� �� 5ީ �X� � `S���/����Z�'� ��e��i ���e&��i � �ަ)� �%%�����Q�����1������(���e��i ��i0��i ��жz�`���d�� ��$�� � ��� � �܅d$ Xݥ)�"�j������,�"���P������$ X�`œ	#� �X� � ���%���2����<���U���U��d$ Xݢ 5ީ��V������
�U���U���d$ X�ڢ 5�����# )�
��U���U�����=�����d$ Xݭ  ��� !� !� !ހ�d�����l������0)��m�e���o���
i��U���U�� X� !ހ���ʥ������$�-� ��2i@�2�3i �3؀��2i�2�3i �3� �ܢ 5ީ����d# ��`ٚ��!�E�E�i�ɛ)����Q�����|�����dd�,����d# ���/�/ �ܥ/������ � '� ���/�� @ީ��(�� ܩ��4�� ܩ��% ҅������� ܭ  ����` @ީ��>�� ܩ��J�� ܩ��Z�� ܩ��f�� ܩ��v�� ܩ����� ܩ
��ɪ���  !� !ހ�  ���� @ީ
� �� ` ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              �?0�?<��WeWeWeW$!eWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeWeW$!eWeWeWe���?0�?�:������<�00��Y�Y�Y�Y�H��Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�Y�H��Y�Y�Y���0000��������?                                                                                                                                                                                    ������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTEEQQTEEQQTEEQQTEEQQTEEQQTEDQDEDQDEDQDEDQDEDQDEEQQTEEQQTEEQQTEEQQTEEQQTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU                                  @                                  @                                  @  � �  � �   � �  ? ? �? ?    �@ �� � ���<� � �  ? ? �� ?�� �C��� �? ��� ?�� � �? ? ��?���C�����? ��?��?�� � �? ?����?���C������ ��?��?�� ? �? ?����?����C�������� ?��?�?� ? �? ?���������C �?����? ?����� ? �? ?�? ��? ���C ����?  ������? �?�?� �� ���C ����  �? ����? �?�?� �� ���@ ����  ��  ��� �?�?� ��? ���@ ����  �� �� � �?�?� ��� ��?@ �����  ��? �? � �?�?� ��� �@ �����  ����? � �?�?� �?� �@�����? ���� � ���?���?�? �@?����������� �? ���?���?�?�� @���������?���� �����������?���� @���������?����  ���������������? @�������?����  ��������������? @����������?  �������������� @���� �����  ��� ����� � ?� @�? �? �? � �   � ���� ?  �  @                                  @                                  @                                  @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTEEQQTEEQQTEEQQTEEQQTEEQQTEDQDEDQDEDQDEDQDEDQDEEQQTEEQQTEEQQTEEQQTEEQQTUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������                                                                                                                                                                                                                                                            ��� 3030��?�  00 30 ?����                    0�?��� �?���������� ������  � ����  3�����  � 0���  3��?��  <�?0���<�? ������  �� � ����  0����  � 0 ���  ��?���  ��0�?�� ���   � �?       �             � � 0�� ��  ?  �?����?          ����0 ��       ��            ? ����?     �  ��                             ��                              �                              �                            ��                            ��                              �   �
          �
            �  �V%     �
  �Z�            � �U$    �Z� XT*         ?��� `  %    `P	 V @�         端� �VU
    `  % X �         ����  ��     �UV
 �ZU)         ����          ��   ��        
����                           ����                       �  ����                       ?=  ����    ����          �A� ����    ����        ? �� l���    ����       ��G�� ����    �?�?�?�?       |�ϒ�� l���   ��������<      �_�?�ڿ? ����   ��������?      p�>@骿? ����   ��������?      \����j�� l���0  �>�>�>�>      w�����������/~   ����     �]�������������  � � � �      ����������� W��0�0�0�0�      |꿚����?����T�����������?�0��������?�����T����������?�<�����������?����ϰ������������VZi���������*����"�ժ������� �ji��������
���*����
����?�3��? 0���������?�����0���������� �eY�eY��� �eY�eY���8 �eY�eY���� �eY�eY������������������������8�������ꋈȯW����oU��ȼW5   lU����W5   lU����W5   lU��� W5   lU��� W5   lU��� W5   lU��� W5   lU��� W5   lU��� W5   lU��� W5   lU��� W5   lU�� W5   lU�� W5   lU�� W5   lU�� W5   lU�� W5   lU�� W����oU�����������������������������ꪪ����������\UUUUUUժ�\UUUUUUժ�\UUUUUUժ�\UUUUUUժ�\UUUUUUժ�\UUUUUUժ�\�U��Uժ�\�UW�Uժ�\W�UW�Uժ����U��Uժ����U7�Uժ�\�U7�Uժ�\��U7�Uժ����U7�Uժ��pU7�Uժ����U7�Uժ�\��W7�Uժ�W�W7�Uժ��U_��Uժ��U_W�Uժ��UsW�Uժ�'\Us��Uժ�<\U_�jUժ��WUWUUUժ����WUUUժ���nWUUUժ����]UUUժ���]UUUժ�����UUUժ����������� �  � �� �� ��  �  �  �  �  � ����������?� ?��? � � � �? � ��?��?����?� ?� ?  ? � � �?  ?� ?��?�� � � � �����������?��? � �\��W\��W\}U]\��_\��_\�\\��\\��p\�\\��\�����_��UU}�W�W��W�UUW�UUW�UUW\��U\��U�*wU��]U��U����\U�_\��_\�Uu\��\��\�
p\�s\��\�p\��_\��_\]]\W]]\_�]\wU\�W�\W��\WU\��W\��U�*wU��]U��U����\�U\�U\W�U���U���U\�U\��U���U�pU���U\��WW�W�U_�U_�Us'\Us<\U_�WUW���W��nW���]��]��������           �������V�`���������   ��� ��������j��j��������� ��: �  &����
                     ������eZ�`�fi�������� ��: �  ��? �p� �\Z��e��e�\Z�p� ��? &����
                     �����ijV�`UU�������   ��� �\��W��ȿ�?��j0������� ��6 �  &����
                     ���������`Uij������   �   �   �   �   �   �   �   �   �   �  �&����
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �� ���ߍ&  p� {� Ƀ p��ߍ&  {� �� @ީ��&  ©��& � � 5� @� Sͩ��  {�9 �r�  �� ����� �X � � �ߍ&  @�L��C �I�B ����@ 	)�@ �  )� ɀ*�  )� bɀ�  ) � mɭ  )� �ǭ  )� �� �� R� �� �� �ͭP ���0�N �(�, ���  {�P 5ީߍ& �, �� �L � v�L� �� F� �í= �t��+ ���c �� S΢ 5ޜ+ �P ����P � � ������> �- � ���  {� ڢ< 5� �����. L�L��	�B ��= ��< ���0 �H �; ����P ����< �����P  v� =ͭ0 �L� �ܭ? ��? �> ����> ��> LM��/ �0 �? �> �H �@ �A �C �B �+ �; �P �9 ���0 ��< �r�= � � � ����`Z���& �, 
���� ȹ�� �܍ ��
 �	 � ��	���)��Z��� iZ� � i � �	 iZ�	 �
 i �
 �ͩ�
 �	 � �	����c����
 �c�	 � �& z`�Z� �	�������Z���Z� �	���%�3� �© �����	�� �	 i	�	 �
 i �
 �; z�`�Z8�1�U ����{���,�=�P�\L��::
���Í轊Íl�T �8�T ����8��T �,�S ���W �V L[ÌT �8�T ����T �,�S �W L[ÌT �8�T ����T �,�S �W �V L[â��&� ����V �]�S ��T �>�W �|�U � z�`��"�=�=�=�=�=�=�=�=�=�=�=�=�=��Z�b�: �
� ���8�9 � ��� ڮ: ��������	������7 � �̩� �� �$  X��: ��	�� � g� ����Цz�`Z�

8�9 �E �< �E �L��8��E �L�Ġ �e� ȹe� �܍ �< � �= � �� �� ��$  Xݭ@ ��:�D �D ��	�A 

��A 

� �D )
m ���� ȹ�� �܍ ��A 


m@ 
��e� ȹe� �܍ �> ���? ��U�% ��$  Xݩ��% �C �Le����C �y�F �E �
8��E i��E ��`�C ���C �T�A � �i:
���� ȹ�� �܍ �C �A ��< 8���< i� �F �= � �G �� �� ��$  X�z`�Z� � �U �����L�ƹ]�V �|�W �>� �� �E ��8��E �ӭU :
���ƍ轑ƍl� LcƭW ɀ����)���LcƭW )
i
�LcƢLcƢLcƭW )
i�LcƭW �����LcƢLcƭW �����LcƭW )
i �LcƢ$LcƭW )
i*�LcƭW )
i.�LcƢ2LcƢ4LcƢ6LcƢ8Lc�L��L��L�Ž�ƍ 轻� �܍ �U ʽ�ƍ �
Ǎ ��$  X�Ls�z�`�Ż������������
��'���,�9�F�K�P�U�Z�]�`ƐR�R�R>S�S�ST^T�T�TUV�V^U�U�UW^W�W�ST�WX^V�VnX�X^X�RڭP ���V�L ��O���U�% �I �E �
8��E �6��E ��-�Q � �R � �I � �J � �, ��Ǎ ��Ǎ �$  Xݩ��% �`	$$$�< � �= � �� ��  �����7�7 ��f���7 � �  ������7 ��� � ���A� �7  �̀�; ����< ���< �#�< �$���9 � ������9 ���9  �­B �Y�= i� �< �  �������@ ��B �7�7 ��0���7 � �  ������7 ��� � ���� �7  �̀��A �B ���@ �
�@ )I�@ `�< :� �= � �� ��  �����5�7 ��8���7 � �  ������7 ��� � ���� �7  �̭< ���< �B �U�= i� �< �  �����5�7 ��8���7 � �  ������7 ��� � ���� �7  �̩�@ ��B ��A �B ���@ �
�@ )I�@ `�B ���@ `�B � �
��B ��@ `�C �w����  ���C �D ��@ �A ��< i�F �	�< 8��F �= �G �H �>� �9��H 8��H حA ��< ::���|��< i��|�= i�>�� `ک� �� �B � �L�ʽ��m= � � �= L�ʭ> ���	� �= L�ʭ �= �< �  �����d�7 ��0���7 � �  ������7 ��� � ���� �7  �̀-�B �	�� 8��= �B �@ )��@ �� i�= �	�B ��B �` ��������









�� �� � � � ��� ���c��>ڠ ��	��8�	��� �8� ����8�9 � ��� � �����ɽ���7 ���&���� �� �=� �\�  ������� `� �J�|����2::�	��.�'� ��>� �� ��  ���������  �� � ������`�C �5�� �� �F � �G �  ������7 �����8���� ��`�� �U �	���� �U�>� �� �U ʽ�ƍ �
Ǎ  �����ԭU ��������ũ� ����  ������m2 �2 �3 i �3 ة�`�> ��? �L�̭< � �� � � �@ ���= � �� ��= i� �� �� �U �	���� �?�>� �� �U ʽ�ƍ �
Ǎ  �����ԭU ��������+ �
� 8� �= `ڭ7 
���� ��� �܍ �`8������  ����9�m2 �2 �3 i �3 � ��/ i�/ ����H i	�H �	���d�? �` �������0 8��0 � ��`�� ��� � ܩ� ��� � ܩ� ��� � ܩ"� ��� � ܩ"� ��� � �`� m � �m 8� � � �7�
�3� � �+� m � �m 8� � � ���� � ����� `��Y�< � �= i� �� �� � � �=� �\� �� ��  �����������= 8��= �	�= i�= `ک���  ��< H�= H�< �C  ��h�= h�< �< �V�� �� ��$ ��e� �e� �܍ �< � �= �  X� !ޢ�e� �e� �܍ �< � �= �  X݀��`���L�Ͻ]�V ��S �>�T �|�W � �U �!�V �]�S ��T �>�W �|�U � 耸::
���ύȹ�ύl ��L�� X�L�� ��L�� ��L�� ��L�� ��L�� I�L�� v�L�� ��L��L�� [�L�� ��L�΀� )�L�� ;�L�� ��L�� c�L�� ��L�� �L�� ��L��`0�6�<�B�H�N�T�Z�`�f�i�o�u�w�}σωϏϕϛ�ڭS ���.���U LVЩ� �� �V ��W ɀ��S ��S � ��S ::� �T �  �����#�T i�  �������V � �T � �S ��W I��W �� �S �W I�W �V �`ڭW �	��W �W ���T ��T �S �S ���W ��U �`ڭW ���W �W ���S �S ��S �S �S ���W ��U �`�S 8��< ��U `Z�V ��S �)�L��V �E�V ���T i�T �T �z�.��V �'�W ���W �W �!�mT �T �W �S �S ���U z`�����W �S � ��U �W �����\8��T ��T i�T ��W `ڭW 	����,���&� ����� �S ��T i�>��]�|�S �S ���W ��U �`Z�V �_�V ��1�T i�T �T �Z�	�K )��?�T �z�8��V �1��V ��W �W ���W �W ��mT �T �W �S �S ���U z`����
Z�V �_�V ��1�T i�T �T �R�	�K )��?�T �z�8��V �1��V ��W �W �
��W �W �{�mT �T �W �S �S ���U z`�����
Z�V �_�V ��1�T i�T �T �JИ�K )��?�T �z�8��V �1��V ��W �W ���W �W ���mT �T �W �S �S ���U z`������Z�S ��U �D�W �W ��:�	��4�W �/���)� �Ȁ��� �S ��T i�>� �]�|��V z`�V ��T �z��U ��T i�T ��S 8�< ����V `��W �W ���2��.�W �)���#� ����� �S ��T 8��>�]�|�`�V ��S 8�< ����V �S ��T �z��U ��S �S �T i�T �W `ڭS ���U �$�W ���W �W �#�mS �S �/�mT �T �W �`������
������
�S �,��U ��T ���U ��S �S �T 8��T `�V ��T ɂ�i�T �W ��T �
�8��T �W ��U `�S ���U ��S �S `ڭ, �������� �Ԁ �Հ �ր &؀ ���`ڭL �L�ծK ���mI � �J � �
� ��  ��������+ �
 5�L�� ����� F�����N ��O ��L L�խK ��I �:��I �(�6�K ���mI �I �M I�M �K 
mM 
���ՍQ 轤� �܍R �2�K ���K ��L �
�O ��O ��L ��O �O ����L LJ��`��X�Y�Zf[Z�K ���f�J �M ���M �p��M �i�M ��	�K ��'�V������� ����]����]�M �4���.� ����K �f֝ �{֝>8��J �!��]�|�M �K  �����N �M ����� ������֍Q 轐� �܍R z`ZJ:JZ:JZ:ZJ:ZZJ:JZ:JZ>\:]6^�O ��O L�׭K �L���L/���L�׭J �f�Ai�J �M )��L�נ���� �Ȁ��� �I ��J i�>��]� �|L�ש�O �K �M L�׭J �:�8��J �M )��L���K �M L�׭I �����M )� �!�I �I �y�K �M �q�M )� ��I �I �`���Z� ����� �I ��J i$�>��]�|�3�I �%����M )� ��I �I ��K �M ��M )� ��I �I �M �I � �J � �� �$�  ������P  v٩��+ �
 5ހ �����N  F�����N �M )
��"؍Q �"� �܍R `2_.`�L ��L L�حK �,�IJ�I�K ���I ��I �K )��1���+� ����� �I ::��J i�>� �]�|��K �K )���؍Q ��� �܍R �K �I � �J � �� �$�  ������P  v٩��+ �
 5� F�����N `*a"c�`�� �� �� �� �< � �= �  ������� `�C �7��3�� �� �� � �I � �J � �F � �G �  ������� `� �(�� �� � � �� �>�  ������ �� `�, ��/��G��`��y�
�N �*�I �r�J ��K ��L ��O �M �Y�%�I �f�J ��M �K �L ��N �=�%�I �f�J ��N �O �L �K �M � �$�I �f�J �
�N �O �L �K �M � ��`�� �P� �	 �`�Z�. �L^� @� c�H�� �� � ܩ� �� �6  �ܭ5  �ܭ4  �ܩ� �*� � ܩ� �*� �3  �ܭ2  �ܭ1  ��h���G���  {��
 5�� �)�� �P� �J�� ܈��� �� �#  �݈�Ω �X � � �� �n� �
 ܭ. :�  Lܩ� �z� � ܜ �n� �� �� �� �#  �ݩ� � �aۍ �b�  Lܭ  ��$������� �ܩ���  �� I� � 5ހ�����  �� ���z�`nz� �X � � �6 �3 ��(�5 �2 �
��4 �1 ��3 �6 �2 �5 �1 �4 ���� `H�Z� �  ~� )��&  �ܢ 5ީ� �P� �� ��  �ݩ� �T� �  ܮ  ���� 5� �ܭ �& ���% z�h`�Z
���� ��� � ��$�-�c��b��]��:�8�0�8�7�  Lܭ8 ���� 5�Ȁ�z�`Z� �c��$��b��%��]��&���� ��� ��  �ޠ ��� Ȳ�� � i0� � i � � ��� � z`ڪ)�JJJJ�  L܊)�  L��`H� �  ���� �2��h`H�  ����h`� �� ���`H�z� h`)?	�`�� ��� �3  �ܭ2  �ܭ1  �ܩ	� ��� �/  �ܩ	� ��� �H  �ܩ%� ��� �0  �ܩ%� ��� �- : ��`�Z �ޮ � �$ � �	�-% ��!���Q�����1��	�-% ��� ��� m � � i � � i0� � i � �Сz�`�Z �ޭ � � �# � ��% ������U�% ����% �% ��� ����I���� ��� i0� � i � � Яz�`�Z�5���� ���� ��z�`� � !�ʀ�`�Z� � ��L��� � � �@� � � ��6� Z� ���%, P8. . ��. . ��. 8. ��z� ���0��� i0� � i � ��Щ� 5�LE�z�`�@� � � � �� i0� � i � ���� m � � i � `��# ���ة��  ��� �� �
� �ߍ& ��" � t ���� �� �� � ����� ���� � �0� ��� �#  ��XL �H�Zx� �� (z�hX@H�Zx�' )��! � ��! ��# �� ��� �� ��� �$ �% (z�hX@� �X �Y �Z  C� G� � � � � � � � �* �� �� � ���� �� `�Y ���%�� � C�z � �{ �  y�� �� �| � �Z ���%�� � G䭇 � �� �  ��� �� ͉ � ��X ���X�Y ����e � C�^ � �_ �  ��Z ����s � G�l � �m �  ��e �e �` � ���s �s �n � �� K� ��`�[ �\�^ ȱ\�_ ȱ\�` ȱ\�a ȱ\�b )
���c ��d �b )0�h ȱ\����� �� Ȍ[ �e �f �` � �L��g  s�� ��\ � ��g ��Ȍg �[ ���w �x�z ȱx�{ ȱx�| ȱx�} ȱx�~ )
��� �썀 �~ )0�� ȱx����� �� Ȍw �� �� �| � �� �Y � �� )�����Z ��  ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��썌 �썍 �� )0�� ȱ������ �� Ȍ� �� �� �� � Ш� �Z � �� )��@З���Y �w  ည�i �j�l ȱj�m ȱj�n ȱj�o ȱj�p )
���q ��r �p )0�v ȱj����� �� Ȍi �s �t �n � Ч�u  ��� ��j � ��u ��Ȍu �i ���� 
���덡 轛덢 ���\ ȱ��] `�� 
���덡 轣덢 ���j ȱ��k `H�Z�a )?	@�� �a I��-� �� �f �c��b )@��J��� �� �h �8��h ��b )0�h Ȍf �c����f �b �f �� � z�h`H�Z�o )?	@�� �o I��-� �� �t �q��p )@��J��� �� �v �8��v ��p )0�v Ȍt �q����t �p �t �� � z�h`H�Z�} )?	@�� �} I��-� �� �� ���~ )@��J��� �� �� �8��� ��~ )0�� Ȍ� ����΂ �~ �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����Ώ �� �� �� � z�h`� `� `H�Z�� ���%�� ���� �� �� )?
���덧 ��덨 ��  ��z�h`�� �* �� `�� ���� ȱ��� ȱ��� ȱ��� )
��썖 �썗 �� )0�� Ȍ� �� �� �� � ~䜩 `H�Z�� ���Lw孓 �� �� I�� )��� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����Θ �� �� �� )�� �� )����
�@����� �� �� �( �� ͝ ��* �� � �� ͔ � ��z�h`H�Z�  s�  ��[ �i ��g �u  �� �� �� � K���X z�h`H�Z�Y � �
�Z � ��� �� )?ͤ �Q�� �K�� 
����x ��덅 ���y ��덆 �w �� � �Y �Z �� )�����Z  �᭣ ���Y  � K�z�h` �� � �
� � �
� � �
� � �
� � �
� � �
� � i
� � |� � �� � �� � |<� � `�� u�� ��� i�� |�� ��� �(� � �� � �<� �     � �
�"8
�" �
�" �
�" �
�" �
�" �
�" �
�" �
�" �
�" ��" �
�"     � �
�" �
�" �
�" ��" ��" ��" ��" ��" ��" ��" ��" ��" ��" �
�" �
�" ��" �(�"     � ��� ��� ��� ��� ��� ���8�� ��� ��� ���  �� ��� ��� ��� ��� ��� �$�� ���     � ��� ��� ��� ��� ��� ���8�� ���8�� ���8�� ���  �� ���  �� ��� ���     �8�"�8�"�8�"�8�"�u�"�8�"�  �"�8�"�u�"� ��"� ��"�8�"�8�"� ��"�8�"� ��"�  �"�8�"�  �"�8�"�     � G�"� Y�"� u�"� Y�"� u�"� ��"� ��"� ��"� ��"�     � � �6� u �6� i �6� � �6� u@��     � ��"� ��"� ��"� ��"� ��"� |�"� ��"� ��"� �@��     � ��1� /$�1�     � u�� `�� P�� :��     � ���     �O�� �� ��� ���   ���O�� �� ��� ���   ���O�� �� ��� ���   ���     � T�1� G�1�     � ��� ��� |�� u�� |� � �� � �� � �� � �� � �� � �� � �� � �� � �� � �� � �� �     � ��  ��  ��  ��  ��  ��  ��  ��  ��  �� � � &�      � � � �~ � �} � �| � �{ � �z � �y � �x � �w � �v � �u � �t � �s �     �
�

		�
	 �
�



	�			�
�������������!�  ����  _���  =�  ��  �  ��  ��  W�i�����k��W������k�������
�쁈�   ���   �o�   ���   �?�   ��>�M�W���PAUSE$C$B$S$T$R$PUSHcSTART$BOUNScGAME$READY$GAMEcOVER$CONTINUE]$END$HIGHcSCORE$YOURcSCORE$NEWcHIGEcSCORE$PROGRAMS$SONGcQI$GRAPHICcDESIGNER$ZHANGcLI$SOUNDcCREATOR$HUcXUHUI$&�,�.�0�2�4�6�A�L�R�\�f�j�u���������J�JKPK�K�KLPL�L�LMPM�M�MNPN�N�NOPO�OPPP�P�P�O�O�O�OQPQ�Q�QRPR�J�J�J�J�J�J�J�J�J�J�J�J�J�J�J�J�J�JpB�B0C0C�CPD�C�DEpE�E�E�F�F0FPG�G�I�IJPJHpH�H0I  ��� �� $(,�zjZJ:*
  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             W���j�