�<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  ����������������������������������������                                                                                  �
      `	    P`�*     �Z�  PVUU)03  �Z�  P`�* 03  `	      �
                             �      30     �           03  �*      03       �      00      �            ���00�  300000   300�00����000030   0000<0   000000�����000   **�*�*�
� ""�  (
�                                                                                                                                                                                                                          �                                                          @           @                                            �                                                                   @        *�
    @U              P    @U        "�     P�         U   P    PU       *     PU��        UU     @UU      "��    T�� @     TU  U    E@U@   �*    T �            @      D    "�     TUTUU  @    U               *�
     TUUU   P @  A@               "        @   P T  PTQU             ���
            PPE   Q T              �""            @UU    @               ��              UU              
     �"              T                �      "                               (P      �    �                          H     �                              �     �    �           @              <�     �                @             �(     �    �                         �     �                              
     "   �                        @�     
          PQ                 @�      �          @Q            �          
   (                    �   ��     "   (                     �   ��     �   (                     �   ��     �
   (                     �   �
      
   (                     �   �
      �   (                     �   �?      "   (                     �   �?      
* (                     �   �?     ����
 (                     �  �?     ���� (                     � <�?      ��� ��                     �@T��?      ��� ��                     �CT��?     �������                    ������
     �����ww                    ������
     �������                     Z�eY�
     �������                     Z�eY�*     �������                     Z�eY�*     �������                     Z�eY�*     ����UUU       ����          Z�eY�*     ��_U���      ����:          Z�eY�*     \U�����󿪪�������?          �����*     ������������������UUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������������������������������������������������������������ ��������������������������������������� ���������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                  @@                                                                          @                                                T                                   @ @                                  P         T      @                          @                                   T                                                                                @           �                                      �                                      ���?        T  U                        �|w�        U PD  U T                  �|U�   0     P  @                  �w�                                   ���?   0                               ��                                     ���� 0                               ���U                                  ��p} 0                             0�?�p}                                0�0��U 0                             0�0���                                0�?�� 70                             0�0���7                               0�0�����0                  @          0�������                               0 ���?��0                             0 ���>���                             0 ���>���           P                p0 ���> ���                           �3 ���? 3�                           @�? ���� 3�3                          ���u= ��������                          ��su� ��������                          ����� �������?                          �� �3 �������:                          �������������:                          ��UUUUUU�U���>                          �������j�U���?                          �eUUUUe�j魪:                          諪������j���*                          諪�����Zi���/                          ��������Zi���*                          ��i]�u]�Zi魪:                          �k������Zi���?                          ��]�u]�Zi���?                          �ꫪ�����j�VU        ���������������������������������������������*������������������������������������������������������������������������������ ��������������������������������������? ��������������������������������������
 ��������������������������������������                                                                                                                                                                                                                      �                                                              @           @                                        �                                                                       @    *�
    @  @U              P    @U    "�     P  P(          U   P    PU   *     P  PU          UU     @UU  "��    T T   @     TU  U    E@U �*   T  T �            @      D "�     TUU TUTUU  @    U           *�
   PQU   TUUU   P @  A@           "           @   P T  PTQU         ���
                PPE   Q T          �""                @UU    @           ��                  UU         �     �"                  T            P*      "                               �      �                               ��     �   �                        @�     �                    @         @�      �   �               @          �< @    �                              �  @    �  �                         �� @   ��                             � @    �  �          PQ              | @   ��              @Q             @ @   �  �                        ��� @  ��                             ��� @   �  �                         ��� @  ��
                              �
 @   �
  �                          �
 @  ��
                              � @   �
  �                          � @  ��
*�                          � @   ���
�                          � @@������                         ���P@ ��� �?                          ���WP���� ��                          ���W�������                         �����������ww                         �������������                         �Z�eX����?��                         �Z�eY����?��                         �Z�eY��������                         �Z�eY��������                      @UUUUUUUUUUUUUUUUUUUUUU                 PUUUUUUUUUUUUUUUUUUUUUU                TUUUUUUUUUUUUUUUUUUUUUU     ����       UUUUUUUUUUUUUUUUUUUUUUU    ����?���������������������������������������
������������������������������������������������������������������������������ ��������������������������������������� ���������������������������������������                                                #    ¯   ���  0   0�?   <�?�  ����  / �� / ���/���/���/��?�/��?������         0 �
�
 ������     �?     �? �
  ���� �������������� ����    ���
        ? ?  ?����      �P`=P=`=`=�    <����<� ������� � 0    �  ����?�?� ���������*�

(�*�*�*�*
(�*�*
(
(
(
 
 
(
(
(
 
 �*�*
(�*�*�*�*
(�*�*
 
(
( (
 
 
(
( (
 
 
(�*�*�*
 
(�*�*�*� �� ����������/�������࿪���������/𪪪���������꯮�����������������꯮�𫪪��𫪪�/�����/���𿪪�����������;���*�? �? � � � �  ���௪�����?��������������ꯪ������ꪪ��뫢��뫪��뫪���꿪��꼪�������𪾪������ ���@   � {�����?�x�7��{�����?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�                                    ��V���                           @��Z��*
�V���                           �*��P������                         TTQ�UUUU�����                        TUUU�ViUQUU�����                        �H�ZRU��ZU�             TP     UU�TT��RU�TU��jUU�            P�Z  @�aUU���@�UU��ZUi�          @TZUUUE@PETUU��JQ�RU������          @EYU��ZQ @@�*UU���VZ�U��jU���           DT���*U AQUU����iU��j�j����           Pe����UUPRT��VJA������j����           TUUU��JUPUUU�@U�V����������           Z��fY�V $j�
Pj��T���Vi�jj��           T�Z��V�j U`YVUURP��jU��������            @UUU��V��UUUU���Z�j���V���               �jDVZ�
DUUEQjU�V�V�U�V���               ZUUUh�ZTa�U����jYUU���              �UQUUI��Ue��j�����j��Z���              PEUUUU�jeP�j���Z�j������Q        �� TTU)UU�jii�Z���UU���������U        jU% EUiU���������ZUU��j��j���UU      �PU��U�%UU��jj�����fUV��Z���U���ZU      �UUE�jUU�����VU�jUY�j�Z���j���Z�      �UUU�VPY�����VUUVj������������Z��      ��VUi�U������U���ZU������������j%��   ��*U���jU�����ZZe��������������������  ����������Z���������������������*�
     �������*������������������������������������������������������������������������fUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��iUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��n�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUﯪjUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUjUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUjUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUjUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUjVUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�YUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�ZUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�fUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��fUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�nUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���oUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUi�kUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�۩UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���eUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UYUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��_UVUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�eVUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���YUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��ߙ]UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���ZjUUUUUUUUUUUUUUUUUUUUUUUUUU��VUUUUUU���_~UUjUUUUUUUUUUUUUUUUUUUUUUU�ZjUUUUUU�ￖzU��UUUUUUUUUUUUUUUUUUUUUU��jjUUUUUU����n���VUUUUUUUUUUUUUUUUUUUUU���ZUUUUUU����k���VUUUUUUUUUUUUUUUUUUUUU����UUUUUU����]���VUUUUUUUUUUUUUUUUUUUUUe龚UUUUUU����jߪ�fUUUUUUUUUUUUUUUUUUUUUi��ZUUUUUU�������n_UUUUUUUUUUUUUUUUUUUUU����UUUUUU��������ZUUUUUUUUUUUUUUUUUUUUU��VUUUUUU����ﯾ�iUUUUUUUUUUUUUUUUUUUUU��YUUUUUUe������UUUUUUUUUUUUUUUUUUUUU���ZUUUUUUe���ﮪ�kUUUUUUUUUUUUUUUUUUUUU����UUUUUUi���믿��U�ZUUUUUUYUUUUU�e�U�����jY�jeU�����������UeUUe�VUUU�U����Z�ZY���Z�j�VU����������믪UUW]VYVUjU����jY�����ejY�����������������_UU�Z�jU�����U���﫪��������������j��j�Z���ꪪꪪ���������ꪪ��������������jeYU�����������뿾�������������������j�������������������뫯����������������������몪��������������������������������������������������������������������������������������������������                                                                                  �
      `	    P`�*     �Z�  PVUU)03  �Z�  P`�* 03  `	      �
                             �      30     �           03  �*      03       �      00      �            ���00�  300000   300�00����000030   0000<0   000000�����000   **�*�*�
� ""�  (
�         #    ¯   ���  0   0�?   <�?�  ����  / �� / ���/���/���/��?�/��?������              *        *                          �      ( �      ( �
      �
      ��   �* Ve   `% Ve  �b% ��* ���� ��/  �b����/  �b�ê�* ��Zsê��������������������                        <    ��  �W  �W `���Z	�� V%���*���������������         0 �
�
 ������   ? ? ? ?  ?������       ? ?  ?����           ?  ? "               ?                   �                 �@���        �P`=P=`=`=�      �
�/����������`��)�
� �� ����������/�������࿪���������/𪪪���������꯮�����������������꯮�𫪪��𫪪�/�����/���𿪪�����������;���*�? �? � � � �  ���௪�����?��������������ꯪ������ꪪ��뫢��뫪��뫪���꿪��꼪�������𪾪������ ���@UUUUYUUUUUU�UUUUU��UUUUU��UUUU����_[������������_U�����TUUeUUUUUUbUUUUUU�VUUUUU�VUUU�����UU�����������������_UUUUUeUUUUUfUUUUU��UUUUU�0UUUUU��FUUE���UU�������������TUYUUUUUU�UUUUUU�WUUUUUWUUUU��VUUUU���QU������U�������U��W���WU�ZU�O���_ZU�*�

(�*�*�*�*
(�*�*
(
(
(
 
 
(
(
(
 
 �*�*
(�*�*�*�*
(�*�*
 
(
( (
 
 
(
( (
 
 
(�*�*�*
 
(�*�*�*    3       ��       ��      ��      ��      ��   <�ã����UUUUUUUUU��������*��������     �?     �? �
  ���� �������������� ����    ���
 �     �     �/  �* �� ���������
�������  ���  ���*  <����<������������������������������������_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�wUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�ת���������������������������������ח                                �֗���������������������������������:֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗   �����������*   ������������   ֗                 �          �   ֗  �������������  ������������
  ֗                           ֗   *    0     *  �
        �  ֗       0        �     ?    �  ֗       �        �    ��    �  ֗       �        �    <    �  ֗       �        �   �
�   �  ֗       �        �   �*�   �  ֗       �        �   ��   �  ֗       �       �   ����   �  ֗       ��      �   ����   �  ֗        �       �   ����   �  ֗      ��       �   ����   �  ֗     � �      �   � *�   �  ֗      ��       �    "0   �  ֗        �       �        �  ֗        �      �    ��   �  ֗                �     ?    �  ֗                �          �  ֗   *          *  �
         �  ֗                           ֗  ����     ����  ����    ����
  ֗                 �          �   ֗   ���     ���*   ����    ����   ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗X}������_U�������W_�UUUUUUUUUUU%֗X}������_U�������__�UUUUUUUUUUU%֗X}�����__U����W�_�UUUUUUUUUUU%֗?<����� ����?���            ֗X}������_U����W��_�WUUUUUUUUUUU%֗X�������_U����W��_�WUUUUUUUUUUU%֗������� � ��?���            ֗X�W������WU�U��W��_�WUUUUUUUUUUU%֗X�W������_U�U������_�WUUUUUUUUUUU%֗X�W������_U�U�����W_�WUUUUUUUUUUU%֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                �          �     ֗                �         �    ֗                �        ��    ֗                �        �0,    ֗                �        �0,    ֗  �   �         ,        8 �    ֗ �� ��
        ,       � �
   ֗ ��+ �/        ,      ���
  ֗ �U� �U�        ,      �?000�  ֗ nU�kU�        ,      �� �  ֗�[U��VU�       ,      �#0��   ֗�[UU�UU�       ,      �� �
  ֗�[UUUUU�       ,      �� �  ֗�[UUUUU�       ,      �#��   ֗�[UUUUU�       ,      ����  ֗�[UUUUU�       �>      �" ��  ֗�[UUUUU�       �>      �#(�   ֗ nUUUUU�       ���      �� D�  ֗ nUUUUU�       ��^�    �*��  ֗ �VUUU�.       ���_    �#( �"  ֗ �kUUU�       @U}�     ��
�  ֗ ��VU��      �����    �    ֗  �kU�+      ������    �g�d  ֗  ��U�      �*  ��    �� `  ֗   �+       ������    ��A��
  ֗   ��        �����     $ ��  ֗    �            |�      8@	�   ֗    (            �_     �P /   ֗                  �     �> �
   ֗                          ��    ֗                          ��
    ֗                           �     ֗                                 ֗  ����     ������             ֗  ����     ������    ������  ֗  ��}��}     �W}��}    ������  ֗  ��}��     ��}���    ��}��}  ֗  ��}��     ��}���    ��}���  ֗  _�}��     @�}��}    ��}���  ֗  ����     �����}     ��}��}  ֗  ����     �����}     �����}   ֗                        �����}   ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗                                 ֗             �������            ֗             �������            ֗             � �����            ֗             �?����             ֗             �?����             ֗             � ����             ֗             ������             ֗             ������             ֗                                 ֗���������������������������������:֗                                ��ת����������������������������������wUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�������������������������������������  0<<����<<�  0<<����>������������<����  �?���������  <<��������   <<���������?  <<���������   <<��<������  <<��<�������  �?�����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���* 0 � � 0 0 0   0������                       \UUUUU          ���? ����?  \UUUUU          WUU5 pUUU5  \UUUUU5          WUU5 pUUU5  \UUUUU�          WUU5 pUUU5  �_���_U         W�5 p��5  �^���~U         W�? p5 p5  �^����U5         W   p5 p5   \� �W�         W   �? p5   \�  _�
        W      p5   \�  |�
        W��?    \5   \�  p�
        WUU5    W   \�  p�
        WUU5   �U   \�  p�
        WUU5   p�    \�  p�
        ��5   \5    \�  p�
          p5   W    \�  p�
          p5  �U    \�  p�
 �����    p5  p�     \�  p�
 WUUU�
   p5  \5     \�  p�
 WUUU�
   p5  W     \�  p�
 WUUU�
   p5 �U     \�  p�
 �����
   p5 p�      \�  \�
 �����
 �p5 p5      \�  W�
 �����
 Wp5 p5 �?   \� �U�
        W�5 p��5   \� pU�
        WUU5 pUUU5   \� \U�
        WUU5 pUUU5   \���WU�
        WUU5 pUUU5   \UUUUU�        ���? ����?   \UUUUժ                      \UUUU�*                      \UUUU�
                      \����� ������ ��������?��? \�����  ������ ��󮪪��;��: \����* �������> ��������;��: \�    ���ꪪ�� ���ꪪ��;��: \�    ���ꪪ�� ���ꪪ��;��: \�    ���ꪪ���������?�: \�    �������������? \�    ��������������   \�    ��������>����   \�    �������:��>����   \�    ��ê�:�:��>����   \�    ��Ϊ�:�:��>����� \�    ��������:������� \�    ��ꪪ���:�������� \�     �������:�������� \�     �������:�������� \�     �������:������� \�      �꯳��:������� \�      ���:�:������   \�      ���:�:������   \�      ���:�:������   \�      ���:�:������  �_��    �?����;�:�������?\UU�    ������;�:��������:\UU�
   ���ꪪ;�:���������:\UU�
   ���ꪪ;�:���������:\UU�
   ������;�:���������:����
    �����;�:���������:����
    �����?�?����������?����
                                                     ������� ����?���� ���� <� <� �������� ��������������� �?������ ��� <���� �������� ������������ �����<��<� �� ������������ �?�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�����_U�����WU�5@�\Ut�5 WU��5��\U�����WU�U5W�\UsU�UUsUU�5��\U�_�UUsUU�5��\U\�UUsUU��5��\U�_�UUsUUU�5W�\UsU�UUsUU��5���_���UsUU�5@� \t�UsUU���W�_���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������*������������*������������*������������*������������*�U  �U   ^)�W5  �U  �W+�|� �U  x�)��U= �U �_}(� _� �U �U(� �U�U ~� (�  W5�U�W (�  |��Ux� (�  �W�U�_5  (�   \�U�U  (������U�����+�UUUUUUUUUUU)�UUUUUUUUUUU)�UUUUUUUUUUU)�UUUUUUUUUUU)�UUUUUUUUUUU)�UUUUUUUUUUU)������U�����+�  �_�U_=  (�  �W�U|� (�  ��U�W/ (� �W}�U \� (� |U�U �U(� _� �U  _�(��U �U  p�*�� �U  �W+�W9  �U   |)������������*������������*������������*������������*������������*������������*������������*������������*������������*�          (�<�<�������+� � ������+�<�C<�     (� � ������+�<�C<�������+� �      (�<�C<�������+� � ������+�<�C<�     (� � ������+�<�C<�������+� �      (�     ������+������������+�           (������������+������������+�           (������������+������������+�           (������������+������������+�           (������������+������������+������������*������������*������������*������������*������������*������������*������������*������������*������������*�  �       (� ��       (� ��/       (� �>       (� ��       (����       (����       (���+�       (�  ��       (����       (��?�?       (����;       (��¿>       (�� �      (�   �       (�           (�           (�           (�           (�           (�           (�           (�           (�           (�           (�           (�           (������������*������������*������������*������������*�����������������hUUUUUUUUUUUUU�  
�_�_���������  �u]�U���]��]�Օ  ��]�U���]��]�Օ  ���W��]]w���  ��]U���]]]]]�]�  �u]U���u]]]]�u�  �_������W]��Օ  XUUUUUUUUUUUUU�               �               �              �              �              �       <       �              �              �       �       �       ��      �       ��      �   �� ��   �  �  
 � ����  �  ������� ��  ����������  ���������������  ���������������  ���������������  ���������������               �               �               �  (             �  
����������������������������������hUUUUUUUUUUUUU�  
XU��_��_��W�UU�  XUuuuWwuWu]WWU�  XUuuuWwuWuuWWU�  XUuuu��_�uuWWU�  XUuuuwuUWuuWWU�  XUuuu�uUWu]WWU�  XUu�_WwU��W�UU�  XUUUUUUUUUUUUU�               �               �               �               �               �               �               �        0      �        0      �        0      �        0      �        ��     �        ��  �  �        ��  0  �        ��? �  �      ����������   �������������  ���������������  ���������������   ������������               �               �  (             �  
����������������������������������hUUUUUUUUUUUUU�  
X�_��_��_���W�  XuuuuuWwuWwUuU�  XuuuuuWuuWwUuU�  Xuuu�_W�_W�_uU�  X�uuWWuW�wUuU�  Xuuuu]Ww]WwUuU�  Xuu�uu�uuWwUuU�  XUUUUUUUUUUUUU�    �?         �  0   ��       �  p  ��       �  \  ��      �  \U T�]     �  PU ��U    �  ST P@    �  �  U   T   �  � P @U  @   �    PQ  T  �  <   T�� @U  �  � C  �  P �  @0  @�  U �  @�p  �S P�  ��?�   WP U�  0 �W    T D�  ��0@   @ �   �
� T   PA�    ?  P��  TQ�    � @��?  р     �   � 0�      �    ���  (         0�  
����������������������������������hUUUUUUUUUUUUU�  
XUU��_W�_���U�  XUUWwuWWWWuUWW�  XUUWuuWWWWuUWW�  XUUW�_WWW��_�U�  XUUWuWWWWUwUwU�  XUUWw]WWWUwU�U�  XUU�uu��_��WW�  XUUUUUUUUUUUUU�               �               �  ���          �  ȼ�          �  ȿ�          �  ȼ��          �  ȿ��          �  ȼ��          �  ȿ��  �      �  ȼ��  ���   �  ���  �3���  �  ����  ����   �  ���������   �  ���������   �  ����� U@U����  �UU�U������ZUU�  ���j�jUUUUUUUU�  �VUUUUUUUUUUUU�  XUUUUUUUUUUUUU�  XUUUUUUUUUUUUU�  XUUUUUUUUUUUUU�  XUUUUUUUUUUUUU�  hUUUUUUUUUUUUU�  
�����������������  ? � ���?���?��� ?                         ���?��<00                                ���?��<00              ���?��<00            ���?��<00        ���?��<00      ���?��<00    ���?��<00  ���?��<00  ���?��<00  ���?��<00    �� �? � �< 00 H�Z����� ����������������� ���r� ~����h�	����������� ������ �������	��������� ���D� ~�L}� ~� ~���������� ���� p��i��� ��	������� p��	8��	�� ��	�\� ~�L˛z�h`xH�Z��
����������������d���������JJ���%�����i����i ��Ɨ��� �Ȁ�Ɩ��� �����L.�z�hX`H� �� �����h`H�Z�/���� ���� ��z�h`H�Z�R����S���dǩ�� �� �����z�h` �� /2�   Ɯ	�����? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                          ����dvdwd|d�d�dީ ��` ��������n�	�  ��x���'������8������?0�?����  ��� ~��̥	��������	���d��  ��0�ޥ��d0dީ��݀ ���斥�)�
� �� {��  � {��`�
�����轶�	�)������ ��`���� ���w }��v�� џ 4�`H�w }� [� {�  ������ ��w�x���v�;����w�w��  � ��ǩ �w  怾�����w�w� 0  � �쀪��w  �Lҟh`H�Z �����d�����@ �����L@���i����+��8󅔽E󅕊
�����	�)�� #��L@�������i� }� [� {�  ���� [��� �� �����L���"����
�  � ��å���̩ ���  �L7���м��� �
ƍ  � �쀝��� ���ƌ  �L7�z�h`�Z��

e���|z�`H�Z��
�����	�)�������+��8󅔽E� �奌i	
�����	�)���i����+��8󅔽E� ����Оz�h`HڽR󅔅�Y󅕅�����
�����	�)�� ����h`H�Z� �
�����	�)�������+��8󅔽E� �����Т ��1�w�����+��8󅔽E�ڊ
�����	�)�� #����z�h`H�Z���d�e����i �� �	����0���e��i ����z�h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���ة��� ���  ��� � �� � � �� � �ߍ& ��"  �� t ����� ��� �� � ������ ��� ��XL �H�Z�� �00�� � � �� �P0Μ Μ �� � �Ν  ��e��e� h��e(z�h@H�$ �% hX@                                                                                          � �� � B� 
� ���< {��� ���d � � ���� ����� �� � �� ���d � ����d 쭍 � � cـ�� �΀�� ]ʀ�� �é ��  � 	쀳�w �x �y �z  ��`�^�Z�_�`�a�T�U�V�W��X�Y�@�P�Q� � �{ ������ �� � �v `��d � ��O� ���� ��� �  x� S� � ,� =� �� [� {�  ����	�����O� �  � ���O�O�Ȋ	����  � �� �O���	���� ���O�O��O  怘�	���� ���O�O�0�O  �L����u�O� �q��$�X�
c�T�0\�8��T�U��X�Y ��F��#�T�0;�8��T�U�Pi�P�Q� �����T�0�8��T�U� ���V�WL��`�O
���� � 轮� � � x�`�4�� ��� �P 9�`�4�� ��� �V 9�`�@�� ��� �T 9�  9�`� ��� ��� �X� xÀ� x���
��`H�Z�
���� 轆�	�)�� ��� ��� �  �� � z�h` �� �� �� �� �� <� :� 9� R� � t� �� �� 
� =� {� �� V� � l� =� � k� ڭ� ���� �  �� {���d�`� �G�I�H0��l �G����G� ����_`� �]�H � �R�: �� �0 ��  �ĩ �� � �Ѐ i߭� ����]�� ���!� H�� � �H �0 8���: 8��$��
Т`�Z�� � i� �� � i�	 z�`� �* � �?�! �� � ��  
ѩ ��  ŭ� ���!� H��
� �* � 8���! 8��.��е`�Z� �l ��#�^ �� �T �  A� �߭� ���
�IȘ�I�����z�`ڭ� i�� � i� �` l� �� ^� |� �� �� ��`��� �(�� � �l ��*� �l �^ 8� �� � 	� 8� �� �� ͗ �� �� ���ʮ� ��l `� �l ��.� �H � � �A�0�A��H �T �0 �^ �: ��A��������`H�Z�w ��;� 8��� � �K � �)�K �	�K �L �M ��K �0�3 �� i�� �= ����z�h`� � � �(��� �$�� � )i {ɼ Ș� �0� � ����`H�Z�w ��Q� �K � �C�3 �� �= �� �K ��� {ɼ3 �����3 ���K �� {ɼ3 ��Ȕ3�y0� �K ��бz�h`�w �/� �N � �!�6 �� �@ �� �
 {ɼ6 �Ȕ6�|0� �N ����`� �H ��!�0 �� �: �� �	 {ɼ0 �Ȕ0�x0� �H ����`� �T �� �^ �� �l ����� {�����`�w ���r � ���r ��Z �X�d `�w ��6�r ��/� �N � �!�@�
��@��N �Z �6 �d �Ȕ@��@����`�w � �6�s ��/� �P � �!�@�
��@��P �[ �8 �e �ȔB��@����`�w � ��s � ���s �P�[ �*�e `�w ��4�r ��-�Z �� �d �� � {ɭ?���?�d �d �)�r ��?`�w � �4�s ��-�[ �� �e �� � {ɭ?���?�e �e �X0�s ��?`� �* ��&� �� �! �� � {�Δ Δ �� � �#� �* ����`� �* �� ���* �t� � Ș�! �����` %�` � R� ��`�=� � � �(� �H�   �`� ٩	 ٩
 �` �� r� �� ��` �� r� �� ��`� ��� �� � �� � {�`�� �� �w � ��  {ɀ��� {ɀ	��� {�`H�Z�
��� ��	�)�� �Q� �@� �0 �� ��z�h`�� �u� �� �� � � �H � ��
��� � �l �p �* �
�I�����M�N�?�@� �) �w � ��  Fʀ��� Fʀ� Fʩ� �� 
i�H�� Ȍ\�]�Z�G� �_�`�a`�� �b��^ ȹb��T �����` �� �� �� W� �� �� O� �� �� �� �� �� {� S� A� �� l� =� ,� k� ڭ� ���� �  �� {���d�`� �G�I�H0��l �G�����M�0��p �G�G� ����_` ��` �` ��`�Z� �l ��*� �&�^ 8�0�� �T �  �� �߭� ���
�IȘ�I������z�` �� �� K�`� �l ��"� ��j ���j �T �� �^ ��  ~ˀ�j �����`ڢ �H � ���H � � � � �� �0 �� �: ������`�p ��$� � �h � ���h ��p �2�X �)�b ��h `� �l ��(� �$�� )�� ̭� �l �� �C�� �T �� �^ �����`�� �� )����� ��� ��
�� �X�� �
��� �)�� �� �� �`� �* � �# �� ���� �� �  }̭� �! ��* ������`���� � � �� �`�p ��4� �0�X �� �b �� � ��  $έi �0�i �b �b �W0�p ��i `� �l ��T� �P�T �� �^ �� �l ��  $ν?�0.� �?�l �� �C��  3ͭ� �l �� �C�� �T �� �^ ��Ș�?�����`ڭ� � �Δ �� � ��� �� � � �� �20� �� �� ��Ε �� �*� �� �� �� �W0� �� �`� �H � �&�0 �� �: �� � ��� � �� �0 �x0� �H �����`ک�
��� ��	�)�� �� ��  ���`� �* � �*� �� �! �� �*  ��Δ Δ Δ �� � � � �* �����`ڭ� 
��� ȹ�	�)�� �� �� ��  ���` ��` #�`� ٩ ٩ ٩ � o�`� � � � �(� �=�   �`�� �P� �� �� � � �l �C�* �H �I�?� ������p �M� �) �j �� �� 
i�H�� Ȍ\�]�Z�G� �_�`�a` !� �� ��  � �� �� C� �� �� d� �� � {� #� �� T� l� =� ,� k� ڭ� ���� �  �� {���d�`� �G�I�H0� �l �G�� ���G� ����_`� �* � �H�! �� � ��  
ѩ �� �� �� �Ѐ ˭� ���� H�� � �* � 8���! �$�����`� �]�H � �J�: �� �0 �� �� �� 
р 'ѩ ��  �Э� ��� � H��� �H �0 8���: ���(譍 ��������`� �l � �A�^ �� �T ��  Gѩ ��  �Э� ���#� H���H�I�]� 8��� ��*�����`�Z� �l � �#�^ �� �T �  �� �߭� ���
�IȘ�I������z�`�Z� � �� �� � �  �� �߭� ����]z�`ڭ� i�� � i� �`�Z�� � i� �� � i�	 z�`�Z�� 8�0� i� �� � i�	 z�`�Z�� � i� �� � i�	 z�`� �* � �;� �� �! �� �*  �ҽ% ��� �% �*  �ѭ� �! �� ���
� �* ��% �����`� �H � �,�0 �� �: �� �H  �ҽH  �ѭ� �: �� ���� �H � �����`H��Ε �� � 0�� �� �(	� � �� ����� � h`� � � �$�� ��� �$��  Z�� �� � �0� � 譍 ���
�����`H�Z�� H�� H)�
���� ���	�)�� ��� ���  ��h�� h�� z�h`Hڨ��
��� ȹ�	�)�� �� ��  ���h`� �l � �j� �� )���T �� �^ �� �l ��  �ֽh � ���h �l ��  9ӭ� �l �� �C�&�h ���h �T �� �^ �� �C �ӭ� �T �� �^ �����`H�Z� �� )� ���� )�� ���� �L��-��� �A�� )������ ��� �+����� ��� ����� � �� ���� ���� z�h`H�Z���Δ �� �0L9ԩ�� �r��� �� �n�b�n�� �[��(�?� ��Ε �� � 0�A� �� �:� � �?�/��+�?� ��� �?� �� �"��"�� �	� � �?z�h`ڭ� ��� � � � � � � � �	� � � �`H�Z� ��� �X� � ��  � 	� [�<�� ��� �
��� ȹ�	�)�� �
� �
�  �� [�  ��� [��  
��d �z�h`H�Z� ��� �;� � ��  � 	� [�F�� ��� � {� [�  ��� [��  
��d �z�h`� � �Z0�� �  ���L���� j�LC���� ��  � 	� ��L��	����*� ��� �� � � �"L�թ"� L��� L�Պ	����*� ��� �� � � � 0L�թ � L��� L�Պ	����'� � �� ���0�.�� �'�=0�!�=� ��	����� � �n��n� � �	����5�P� �.� �0'� �) �) ���8�P��Pح� �� Dր I�`� �* � �, �� �� � �� � ��  =ԭ� � �� �! �� �* ������`Hڢ �H � � =ԭ� �0 �� �: �� �H �������h`� �l � ��T �� �^ �� �l �� �  �������`� � �� �� � �� � �� Ζ  ��`ڭ� 
���� ȹ��	�)�� �� ��� � �  ���`�� �$�T �V �T�U �W �<� ��^ �_ ��` �a �� ��l �m � ��n �o �* �+ �, �- �H �I �% �& �' �( �. �/ �I�J�K�L� ���������	� �) ��h ��i �(�j �2�k �?�@�A�B�� 
i�H�� �� Ȍ\�]�Z�G� �_�`�a`� ٩ ٩ ٩ � �`�� � � �(� �/�  0�`H� �d�m � ��i � � �U��� 0��� ��h`�  ٩ ٩ ٩ � K�`��� ���� �P 9�`��� ���� �V 9�`��� ���� �T 9�  9�`� ���� ��� �X� �؀� ����
��`� ���� ��� �X� �؀� ����
��`�i�
��`� �`�	�)�� �z� ���  ���`�
��`� �`�	�)�� �z� ��� ��� ���  ��`�� � � �(� �g�   �`� �� �� �� Z� � �� �� �� �� �� �� {�� ��� �� %� �� -� �� l� =� ,� k� ڭ� ���� �  �� {���d�`� ���� �D�� � xà �  ��
 {���d�� ��L�`�Z�\ʎ� �� 

m� ����| z�`�F�� �
�� � �� �Z� �<�� ����)����!������
 �٢��� ������� � ����� `�_���0 �٭� ���� ���w ���x ��Z�D��Z �� �� ���4�a��� ���^�^��
��Z�^���Z��`��� �ک�Z`�\ʎ� �� 

m� �����mT�T�U�`�Q�P�_����W�V�Y�X�U�T�#�V�W�T�U�a���
��X�Y��Y�X`H�\�V��8�V�8�X�]�X���X����ah`H�P� ��R�<�
�R���`��Rh`�l ���I�H0��l �G�m ���J�H0��m �G�n ���K�H0��n �G�G������_`� � ���$�  ��� � ��� �� ���%� ��������� ���&� ��������� ���'� ��������� �� �2� ��������� ��!�3� ��������� ��"�4� ��������� ��#�5� �������`H�Z�� �� )�
���� ���	�)�� ��� ���  ��z�h`H�% � �*�! �  �� �ݭ� ���� H�� �% ����ʎ��$�& � �*�" �  �� �ݭ� ���� H���& ����ʎ��%�' � �*�# �  �� �ݭ� ���� H���' ����ʎ��&�( � �*�$ �   �� �ݭ� ���� H���( ����ʎ��'h`�Z� �i� � �i�	 z�`H�Z�l � �(�^ 8�/�� i	�� �F� �Y�  �߭� ����I�\�m � �(�_ 8�/�� i�� �-� �;�  �߭� ����J�-�n � �&�` 8�/�� i�� �� �%�  �߭� ����Kz�h`H�]�H � �*�: �0  M� i߭� ���� H��]��H �g� ��2�I � �*�; �1  M� i߭� ���� H��]��I �g�!��3�J � �*�< �2  M� i߭� ���� H��]��J �g�"��4�K � �*�= �3  M� i߭� ���� H��]��K �g�#��5h`�Z� �i� �i� i�	 z�`H�Z� i0�� i�� �t� ���  ��z�h`H�Z� ͗ 0͘ 0�*� ͗ � � � 0� 0��	 � ����� �� �� � z�h`H�l ���h � �� �l �+�^ ��h �m ���i � �� �m �-�_ ��i �n ���j � �� �n �.�` ��j h`H�l � ��D �0�D �Y�^ i� ����D �m � ��E �0�E �;�_ i� ����E �n � ��F �0�F �%�` i� ����F h`�Z�G ��F�H � ��H �0 �: �4�I � ��I �1 �; �"�J � ��J �2 �< ��K � �	�K �3 �= z�`H�l � �.�^ �Y��^ �S � M��?�?�0�?�^ �
��l �2�h �m � �.�_ �Y��_ �S � M��@�@�0�@�_ �
��m �<�i �n � �.�` �Y��` �S � M��A�A�0�A�` �
��n �F�j h`�� ��S � ��l �m �n �I�J�K�H �I �J �K �% �& �' �( � �������� �) �2�h �<�i �F�j �� i�H�� Ȍ\�]�Z�G� �_�`�a�� ������ �� �� `� � �Z0�� �  ���L������ � � j�L�� ��L����� ��  � 	� ��L��	����� � �"�!�"� ��	����� � � 0�� � � �	����5�P� �.� �0'� �) �) ���8�P��Pح� � � '� ��`�  ��� ��  � 	� �� � ��L��� ��$�� �� �L��� � � �0L���� �P���� �� �
0B�� ��� �8��/� ��� �� �0#�� � � �0�� �� �20;��� ��L��P� �L��� � �0� �) �) ���8�P��P� '�`H�% � ����% ���� 0�% h`� �S �  M�`�% � �*� �� �! �� �%  ��Δ Δ �� � �� �% �) �& � �*� �� �" �� �&  ��Δ Δ �� � �� �& �) �' � �*� �� �# �� �'  ��Δ Δ �� � �� �' �) �( � �*�  �� �$ �� �(  ��Δ Δ �� �  �� �( �) `H�Z�
���� ���	�)�� ��� ���  ��z�h`H� �H � �$�0 �� �: �� �H  �䭔 �0 �x0� �H �G �����h`H�Z��
���� ���	�)�� ��� ���  ��� � z�h`� �% � � ���% �t� � Ȕ!������`H�Z�
���� 轴�	�)�� ����� ��� ��� �S ��  ��z�h`H�Z




�� ��)� �& z�h`H�Z�� �d�m� � ��i � � ���� 0��� m � � i � � ��z�h`H�Z�� �d�m� � ��i � � ���� 0��� m � � i � � ��z�h`H�Z� �d�m � ��i � � � ��� 0��� ��z�h`H�  ���� g�h`Hڭ  �����h`H�� �  ����� �0�h`�Z�P���� ���� ��z�`� � � � � � � � � � �( �) �* `H�Z�� �@�� � � � ������ ���z�h`H�Z�� � �孖 
���� ��� � ���$��a��b��c��d�8�7��  V�Ȁ�z�h`H�Z�)�JJJJ��  V�)��  V�z�h`H�Z�)�JJJJ��  ��)��  ��z�h`xH�Z�� �a��$��b��%��c��&��d��'������ ����� ��� �� �d��� ���� �� ����� Ȳ���� �Ζ ��� � z�hX`xH�Z�� ������ ����� ��� �� �d��� ���� �� ����� Ȳ���� �Ζ Б� � z�hX`H�Z� �� ��  � 	� � � � � � � � �� �� �b�c��ez�h`Hڪ�� ���b����� �b���c�h`H�Z�c���C�� 
����� ���� �b

����$�* ȱ�



�� �� ȱڍ) ȱ�� �( �b� ��z�h`�c�* `�� ���Q�� ���.�� � 쭰 �� � �  ��� � 	쭽 �� � �  Q�� �� Ͳ � N��� �� Ϳ � .꭬ ���.�� � � 	�� �� � � � �  ���� �� �� � ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��V��� �V��� Ȍ� �� �� �� � �L�鮹 �d�� ���� �� ��� ��� � ��� ��莹 �� ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��V��� �V��� Ȍ� �� �� �� � �#� ��  � 	쭰 �� � � �� �� � � `�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��V��� �V��� Ȍ� �� �� �� � �4�� �d�� ���� �� ��� ��� � ��� ���� �� ��`��퍮 轴퍯 `�&��� �&��� `��퍮 ��퍯 `��퍻 轾퍼 `�:��� �:��� `��퍻 ��퍼 `H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����θ �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� �ª�� )@��J��� �� Ȍ� ������� �� �� �� �� �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� �ͪ�� )@��J��� �� Ȍ� ������� �� �� �� � � �� �� z�h`� �� `� �� `H�Z�d�� g��� N� �윭 �� ��� ��  N� .� �� Q���� z�h`�&��� �:��� �'��� �;��� `��퍮 ��퍻 ��퍯 ��퍼 `��퍮 ��퍻 ��퍯 ��퍼 `H�Z�L��� �M��� �� ���  �� ����� z�h`H�Z�N��� �O��� �� ���  �� ����� z�h`H�Z�P��� �Q��� �� ���  �� ����� z�h` �    �� �� �� �� �    _�  d�  j�  q�  w�  �  ��  ��  ��  ��  ��  ��  ��  /�  2�  5�  8�  ;�  ?�  C�  G�  K�  O�  T�  Y�  _�    ��0�t���  �c���"�  z��a�  ��*��  ���� 

  � �� �� �� � �� �� �� �� �� �$�    � �� �� �� � �� �� �� �� j� d$� � d�    d� T� Y� q� d� d� Y� d$� � � � d� � �� �� �� �� �$�    � �� �� �� � � �� � ��  �   ��T�h�.� ���h�.�@���T�h���T�h�.� ���   h�.�@���T�h���T�h���T�h���T�h���T�h�   ��T�h���T�h���T�h���T�h�.� ���.� ����    �� ����T�h���T�h�.� ���.� ���.� ���    �� �� �� �$� � �� �� �� �� �� �� �� ��.B� �� �� ��.B� � �� � �B� K� T� _� d� q�    w� q� d� d� �� _� d� _� T� _� d� q� w� q� d� d� �� K�    T� _� d� q� w� q� d<� �� � �� �l�   .0���}����$� �.�T�}�����������\B�������\B� ��� ��.B� �� �� �� �� ��    �� �� �� ��.� �� �� �� �� �� �� �� �� �� �� ��.� ��    �� �� �� �� �� �� �<�.� ���   GAMEaOVER$YOUaWINd$aSINKINGa$NOaWEAPONd$GaTaC$����������3�#���ˎ���g�˗/�M�������$$$""""	 Ir	,Or+/Su$$$$+T}6Y|�@PEXE�PQ�QR"R� �*((((
(
H �=���  ���    ��  "$.R�R3S�S	tF-�S�S�S�SnZF2�ST+TCT�T[T�UOU�U�U/V9VCV�VW9WqW	
6�F�(D��|��� H ��<!L!===
((((
....,!,/////!/////+ /wW�k�k�k�k�$	!�}}} �� �� q� q� q� q� q� � j� �� ��    j� �� �� 5� K� K� �� �� � � � � �    �� q� �� �� q� �� �� 8� T� T� �� �� T� T� T� T� T� _� j�    q� q� j� q� q� 5� 8� 8� �� ��    _� _� _� _� _� j� j� _� _� _0�    �� �� �� �� �� �� �� �    � � � �� j� q� q� � � � � �� � q� q� � j� q� Y� q�    T� T� T� _� T0�   T�T������.�    ��}�}�}� ��T� ��T�T�T�}�}� �� ��}� ���}����:�    ����� ���� �� ���� ���� �� ���   :� ��:���� ����:��}� �����}���:��:���� ��   T���T���:� ��T���   }���}������:���}�}�����}��:� �� ��.��    �� �� ��� ��}���}���}���}���   �
	�
	�
�

		�		�		 �����4����� � �+���  ����E������� ���  ��/�  ������������ 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  W� ���