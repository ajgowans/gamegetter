�� �� �"�;�� �� ��/�� �� �
�#�� �� 0�� �� �� �� �� �� �� �� L ��� ��Ly�L��                                                                                                                                                                                                                                                                                                                                                                                                                                            �ȍ� ���� � ���	�f �(�g ��� �(�� �U�� � ��  (ũ��� ����  \� (� \�d�g ��� ��� �
�f �� iK��  (ŀ����f �� iK��  (ũ�f �� iK��  (ũ�f �� iK��  (ũ"�f �K��  (Ů   ����Ή �� � ����� ��L��Ly�          � �? �<�<�<�<� <� << ?< ?<�<�<��� �? �               <  ? � � � � �  �  <  ?   � � � �                 � �?�������  �  ? � � ? � � � ?��?��?                �? �� ?� �  �  � �? �  <  <  <�<�?����                 �  � �� �� �� << ?<���������� � � �                �� �� �  �  <  ?  �?�����  �  �  �  ?���                  � � <   � ������?�?�<� <� ?������                ��?��?�  � � � �  �  <  <  ?     � �                 � ��?�<�?�� �������� < <�����                 ��?�<� <� <� ?� ?�� � � � �  ? � ?                                                                                                                                                                                                                                                                                                                    ������  03  �  �� ������ ������  �� � � �  �  <�    ������  ��  <��?0������� ������  ��  <���� ��   ������  �� ����0�������� ������  �<�3<��0������   ������  ����0�0��3������� �� ���  �30�<<�����   ������  0�0��03�3�������� � ���  � ���� 033����<�    ������   ?���� 033������    �� ���   ����03�3���� ��� ������   ���30�<<���<�   ������  �?��0�30��3��<��� ������    ��3��0�����   ������  �������0������� ������    <<�����<3�   ������  ���<��?0��<3��� ������    < � � �  �����    ������  ��  �  �� �������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           H���� �*�� ��� ��� ��; ���< ��� �< �g �; �f  (ŭ< �u�� ��  \��< �� ���� �ө�d ���e ��� �< �< �g �; �f �*�� ���  (��e �e �e �g �d �f �� �� �+��  (ŭe �H0� ��  \� �� � ����� ��� ��  \� \�< �g ��� �; �f �*��  ŭ; i�; �f  (ŭd �f �+��  ŭd 8��d �f  (ŭd �� \��� ^� ��  ��� �� hL� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          g� n���� ����  <�(�� ��� �W�� ��f ���g  (ŭ� �1�� �g �>��g �@��  \��߮  ���L �     �                                     ���                                     ��                                   �? �                                   � �                                   �  ?                                   �   ?                                  �?   ?                                  �                                     �                                      �                                       �                                      �?                                      �?                 <                    �                 �                    �                 �    �   <          �                ��    <   �          �                ��    ?  ��          �                ��    �   ��          �                 �0   ��   �0�        �                ���  ��   �0�     ?  �     � ? �     �   ��  ���     ��  �    �<�� �<  �? <�  �<     �� �� �    ��3��?0� �� <���? <��3��  �   ����<���� �0�� � ?� ?�?<�  �   �����3�,�?�����������?�3  �   ? <0������<�< ������?�  �  �? <�<?����0<�?��� <?���?0?  �?  �< ��00��?� �?� �����  �� �?���<��<<����������<���   ����?� ������<����?����0��??���   ���  � ������� �?��?�������?             �                        �            �3                                      �?                                      ?                                     �                                     ?                                     �                                     � �                                    < �                                     ? �                                      <                                      ?                                     �                                     �                                     ��                                      �?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                      �                                 ���  �                                ����� �                                �������?                               ��������                               ���������?                           ������������                          �������������                          �������������                           ������������?                            �����������?                            �����������?                           �������������                           �������������                         ��������������                         ��������������                        ���������������                        �����?�?�������                         ��?�� ������                          ���� ������<                         ���?  �������                         ���?    ������                         �� �     ����?                         ��  �    ����?                         ��     �? ����                         ��     �� ����                          ���   �� ���?�                          ���   ?  ����?                          ��� �  ����?                          �� < �   ���                          � � ?�  ���                           �    ���                           �0 �0  ���                           <<� �<�  ?��                            0���� �?                            ����� ��                            �����  �                            �< ��  0                            �0 �0  �                            ��3 <  �                            0��0 �  0�                             0 ?<      �                             0       ?                             0  � �  �                       0     �    <  ����                       �   ��  �5  �                         � � � ��U   �?                 �   � � � �UT   <�               � �   ��? 0  < |QU                    � 0� �U� ��� WUU     0                 �  |U�    �UUE  �  �               0 0  WU�=    _UUU  �  �               0�   WUU�   �UUU  0  �         ���(
��  �WUUW �WUUU5��? ��                �   �WUU_��UUUUT� 0 �<                   �WUU}UUUUUUUU?  0<�                   �WUUuUUUUUUU�  �0�         �����"���
 �WU�UUUUUUU<   �                     W��UUUUUEU    �                     _��UUUUUU�                      0�    _� �WUUUUU|=                      0    |5 �_UUUUEE=                            �5  ~UU�UUU�                            �7  �UU�UUQ�                        �  ?  ����UUU�                            �   � pUT�                            �  ? \UDU�                            �    WQ                    �       �   �UUT                     �       �� �UUAE                    ?        �� �WU U@                    ��         �  _UA                       ��      � |�                         ��       0�E� �?     (               <�      �� �   ��� �               �"�     �� �  ��� �*               �*���
  �  � �    
 �(* *             �" �  �     ��   �  �����               �   �?
  *�   � ��*��
           � 
�
�( �

�   ��
�����*            ������* �

�   ���������            :  �*� � *2��
  ���* ���           �
  �� �� �2��*  � �*��
�           *���  �"�(( �2(�� �( *
�*�
           ���  �( 
 �3��� �*� �*(          ����0  �(��  ���ʠ� �� ��            ��
��� ��
�     �   ���  ��            �� �p3 ����   ��
�( 0�
   �
            * �� ���(    � ܌ � �            
  p �
(     0
�00 �                 7�  � �?��??ܠ
p3�                     7 �* �����?0���0 ���                    �   ���à  0�}ss                 �          �}#  � ���                  p3          �0  03 07                  ��          0�  �� �7                   0          �0  00 0           ������������� ��  0��  �����?        ������������� ��  ��  ������        � �����1 �_ ��?   � ����� �        � ���  � ��? �   �������  ?        � ���  0 �� �  ��?����  �        � ���  � �� �  ������  �        � ���  0 �� �  ������  �       � ���  � �� �  ��� ����  �       � ���  0 �� �  ��? ����  �       � ���  � �� �  �� ����  �       � ���  0 �_� �  �� ����  �       �������� �� �  ��  ����  �       ��������0���� �  ��  ����  �       � �������_� �  �� ����  �       � ���  0� � �  �� ����  �       � ���  ��� �  ��? ����  �       � ���  0��� �  ��� ����  �       � ���  � �� �  ������  �       � ���  0 �� �  ������  �       � ���  � �� �  ������  �        � ���  0 �� �  ��?����  �        � ���  � �_�? �   �������  ?        � �����1 ���?   � ����� �       ���������������  �� �������       ���������������   �� ������?                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ��
��*�     �*��
��*                   "                                 "                                 ��
��
�      �
   �                                �*"                                  �                      ��
�      �
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     H�@��  <��� ��� �@�� �
�f ��g  (ũ�� �B�� ��f  (ũ�f  (ŭ� i4�� ��f  a��� i4�� ��f  a��� i4�� �!�f  a��� i4�� �#�f  a��4�� �%�f  a���� ��� �A�� ��f �,�g  (ũ�f �� i4��  a��� i4�� ��f  a��� i4�� �!�f  a��� i4�� �#�f  a��4�� �%�f  a���� ��� �E�� ��f �K�g  (ũ
�� �G�� ��f  (ũ�f �b�g �� ���i4�� ���  a��� ���i4�� ��f  a��� ���i4�� ��f  a��� ���i4�� ��f  a��4�� ��f  a��
�� ����  \�Β �� � ��� hL �� � � � � � ��00 0  � �?�?    000�  �0�?  �?0 � 0 000� � 0 �0000��?  � � � � �0000�0000��0000�? 0 ��000<03�000��������� ��������  ����������?����� ������������������<� ���<�����<����<�����������?��� ���� ���  � ��� ���  ��  �  �� �� �� �((���������*�
��<��������� �?<��������� <<��� ��  <�������  <������� <<��?� �� �?�?������� �������� ��<<�?�?�??<<�?<<?<< �<�<<��<?<�?<<?< <�?�?<�?�?��<�� ��  �� �� �0 3 �0 �? �?� ��   �� ̪ ê � �         �   �  ��  �� �� �0 3 �0 �? �?� �?0  0�  ̪  � 0� �6 ��7 �7 �� �  �?  �? ��� �_U ��� ��� �U]  WU  T  �
  h  f  �� V� h  �5  �?  �  TT  _�  ?�                                                                                                                                                                                                                        H�L ��@�� ��� �5�� ��f �A�g  a��5�� �U�g  a��@�� �ȍ� �   ����������hΒ  \� � ��ߩ�� �T���6�� ��f �A�g  a��5�� �U�g  a��ȍ� �   �������"����Β  \� � ��߀���� �R���G�L�7�� ��f �A�g  a��5�� �U�g  a��ȍ� �   ������� ����Β  \� � ��߀i��� �R�����8�� ��f �A�g  a��5�� �U�g  a��ȍ� �   �������,����Β  \� � ��߀������ ��� �� �� �hL�©9�� ��f �A�g  a��5�� �U�g  a��ȍ� �   ����������Β  \� � ��߀���� ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �@�� ��� ��� �@�� �
�f ��g  (ŭ� i4�� ��f  a��� i4�� ��f  a��� i4�� �!�f  a��� i4�� �#�f  a��4�� �%�f  a���� ��� �B�� ��f ��g  (ũ�f  (ũ�� ��� �A�� ��f �"�g  (ũ#�f �� ���i4��  a��!�f �� ���i4��  a���f �� ���i4��  a���f �� ���i4��  a��%�f �4��  a���� ��� �>�� ��f �@�g  (ũ
�� ��� �?�� ��f �T�g  (ŭ� � �@��f �r�g �J�� ��� ���  (ŭ� 8�� ���f  (ŭ� 8�� �� �f  (ŭ� ����� ���	�� L�LG���f �A�g �� ���i4�� ����  a��U�g �� ���i4��  a����� � \�   ������ ��L��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �@��  <�� � �3�� ����� �%����� ������ ���� � �� ���� L ��� ��
�5�� �)L ����6�� ����7�� ����8�� ��9�� ��f �A�g  a��� ���5�� ����6�� ����7�� ��8�� ��f �U�g  a����� ���  \�   ����
Β �� � ��L��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �@�� �� � ��� �� �a�� � ��	�� �� �� �M�� � ��	�� �� �� �� �6�� � ��	�� �� �� �� �� ����� � \��� ���� ���L �L ��� �
0%�� �� � ��� �
0�� �� �� �
0�� �� ��f �b�g �� ���i4�� � ��  a�����  a���f �� ���i4�� � ��  a�����  a���f �� ���i4�� � ��  a�����  a���f �� ���i4�� � ��  a�����  a��#�f �,�g �� ���i4�� � ��  a�����  a��!�f �� ���i4�� � ��  a�����  a���f �� ���i4�� � ��  a�����  a���f �� ���i4�� � ��  a�����  a�L �L �                                                               H��� ��� ��f �x�g ��� �� ��H��  (�� ��� �0�I��  (�� �� hL���� ��                                                                                                                                                                                     <�� � �L �Lq� <�@�� � �  g� n��� �� �� �� ��� ��� �F�� ��f �M�g  (ũ�� �n�g �D��  (ũ�� ��� �C�� ��f �p�g � ��  (ũ��� �O�g  (ŀ��L/©��� �  ���K���GΒ �� � ��P��  \���ߩ���  \� \� \� \��� ��� ���  ^� ��L�� ����L/� �𩴍� �O�g � ��  (ũ��� �p�g  (Ů  ��������Β �� � �ƩP��  \���ũ���  \� \� \� \�L/�������� �?<��?�?���� �����<����<��� <����?<����?<��?��<��?<<�?�?�??<��??<<�?<<?<� ?<<  <�<� �<<� <?� ?<�<<?� ?< �?�?<��?<�?�?��<��?<��?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              H �� Э� ������ �� ��� �L�� �O�� �� ��  �� +� �� �� ���� �%�� ����  �� +� �� �� ���� �� �� �0��  \�h`�� ����  �� +� �� �� ���� �֭� �ʩ��  �� +� �� �� ���� ��H�� �� �� �� ��� �� ��� h`H�� �� �� ��� h`H��� �? ��; �,�{ �} � �� �C �D �E �F �G �H �i �j �k �d �Q �S �t �v �� ��� �P�� �F�| �~ �� �� ���K �M �T �=�� ��� ��� ��� ���� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �Z �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� � �� �� �� �� �� �� �� �� �� �� h`H���< �z�R h`H�r�< �d�R h`H�r�< �F�R h`H�p�< �n�R h`H���< �\�R hH���< ���M �z�R h`H���< �v�R h`H�Z�� � �m�� ��?�� �#��4��9��?��J��A�� �<�� �� �,�Q �x�R �*�� �%�� � �� ����� ������� ���"���%���� ���@ ��� ���� ���@ z�h`�� �(8�
�����9 轣��: �� 8� 
��9�� ȱ9�@ �ͭ� ��� ���@ ��H��� ���@ h`H�� ���� ���� ���� �� ��� �<�� �h�@ h`H�� ��Q�� ���� ���@ �<�� �(8�
�����9 轣��: �� 8� 
��9�� ȱ9�@ ��� ��� ���@ h`�� ���,�Q �\�R �� �� �0	�-8����� 
������ ����@ Lȃ�� 8�-
��-��� �-��@ LȃH�� ��$�� ���,�d �t�e ��� �F�
�,�Q �n�R �*�� �z�@ h`H Ƅ�� �0f ꄭ� ��\�3�� ��� ��� �� �f �� �g  (��� �<07�� �� �� � ��� i�� �Z��� 8��� �F0	���� �� �� h`H�� �f �� 8��g ��� ��� �3��  �h`H�; i�� 0C�; 8��� 8�< i�� 0-�< 8��� "�� i�� ��� �,�� ��� ���� � �h` <� �� 5��,�� �P�� ��� ���  +� �� ��R  +� ��  � �� _��R �R � ���R  3� _��R �R � �� �� �� _���R  3� _�  � +� �� _��R �0 \�R � ���� �R��  �� @� _��� � ����� ��  `�<�R   � �� _��R �R � ���� �R��  �� @� <� +� �� _��� � ��  ���R  3� _��R �R � ���R   � +� �� _��R �0��  \�R � ��`�  ��L/�`H�Z�� 8�
��鈍9 �鈍: �� 8�
��9�7 ȱ9�8 �� 
��7�9 ȱ7�: �� 

��9�c�ͥ ȱ9ͥ �� ��� �� z�h`�� ȱ9��*��,��.��0��2��4��6��8�	�:�
�<��>�H�d Lm��Q Lm��S Lm��C Lm��G Lm��H Lm��F Lm��{ Lm��} Lm��i Lm��j Lm��E Lm��������������LÆ�k Lm�� Lm��t Lm��v Lm��� Lm�H�Z�� 8�
��鈍9 �鈍: �� 8�
��9�7 ȱ9�8 �� 
��7�9 ȱ7�: �� 

��9�c�ͥ ȱ9ͥ �� ��� �� z�h`�� ȱ9������"��*��,�6ȱ9��  M�L��ȱ9��  �L��ȱ9��  2�L�� ��L��ȱ9��  ��L������"��*�	�2�
�:��B��J�Tȱ9��  ��L��ȱ9��  ��L��ȱ9��  ��L��ȱ9��  �L��ȱ9��  ^�L��ȱ9��  ��L��ȱ9��  9�L����������&�ȱ9��  l�L��ȱ9��  ��L��ȱ9��  �L��ȱ9��  S�L����������#�'�+�/�3�7�;�?�C�G�K�O�S�W�[�_�c�g�k���������ԉى����6�G�`�i����������,�9�B�O�`�m���������ދ���.�?�`�m��� "�(3�3>�>I�Yd�c HSxc ! " !,x)4 ?J�Wb c :Hnc U	U +U#.v:E
vFQvS^ c,7 c(3 2= NY
gc(3 4?xBM c" 'n&1 ,7nBM R]}U` c(3v6JxHS c U$
v)	U*U(3vc6A 8CF9D	F>I c"
w"w(x) 6A >Iscw2=
vc� P$	P.9�3>P<G�@KPP[tWbtc�	P$
t) -8t6A�<GPALtIT P[tVatc
    +
v,7v6A CNxLW c#x!, +6x@Kxc !,v8CxHS R]vc
 ' +6	ZEPZHSZcs %UCN c
 />x=Hsc 2= c 8C HSxc 'xNY
vQZvc=H LWZP[	Zc
  #.
v7B 9D DO FQxcvv#x + *5 AL c $ -8
�cc 
t$t#.t(3t/: 7B	P<G�@KtGR�KVPc +6 4?�GR cx (3 <GxXcU\g	Uc
 -8F7B <Gdc' !,n@K�R] U` c}&1
v7B IT c 
��
�!�$�2=�7B�c! 8C HS c  �"
t#.t.9�0;P5@	P=H P[tct '�!,P(3t7B :EtIT c��Ɍьٌ������������	������!�%�)�-�1�5�9�������1�~�����9�z�Ǐ��5�n�Ð�9�����9�����$�=�������=���ϔ �a���˕�i�Җ�� �%�&�
SS�
�
�
�S&�
,�
.SCSGPUPVPZ�
[�
c"w+F,F0wBnCn_!t`"tc%t&t
FFF'n(n1n2n7}8}AwMxNx\z]z`}a}lwcwK#K.K2w5K?x@xJnKnNdOdSsTs_!t`"tc%t&tK w#K%w*K+K7K8K<|
A|
FKGKHKV|
[|
\|
a|
c'r(r-F.F1F8m
B^
HrIrU|
V|
Z|
_!t`"tc%t&tdd,{
0F1F8v9vAvBvFnGnbFc
KKvvw!|
"|
$F%F7m
D�E�HrIrR^
Y2`!ta"tc%t&tKKK,|-|@wDKIzJzNzOzTwiFjFcFF	|

|
nn#|
$|
(|
EnFnJsKsOxPxU}V}_!t`"tc%t&tF
|
2F3F@|
A|
LwZK[F]Fc<<wF!|
'n(n/F8m
B^
C(D(YF_!t`"tc%t&t+|
,|
2F3F9m
NwQFRFXF^F_FcwcFF|
|
AA&w.|
/|
2|
3|
7AAwEwIwMwQwUFVF_!t`"tc%r&r1�	 2�	+1�	,2�	6F7FS1�	T2�	c1�	2�	FF'1�	(2�	51�	62�	?1�	@2�	C1�	D2�	HFO1�	P2�	Q1�	R2�	_!r`"rc%t&tBFllw#F$F-|
.|
3F4F9F:F>v?vCsDsHdIdTvUv\|
]|
b|
c|
c
KKwFFwFF'n(n1�2�IFU!tV"tc%�&�&F'F/F0F3|
4|
<F=FKFZKc5F=K>KI�J�OPQP_!t`"tc%t&t|
|
|
w*F/F0F6m
7m
?n@nDsEsIsJsQ^
iwcwF	Fh2737?d@dDdEd_!t`"tc%�&��
�
P�
 P!P"�&�*�.�2�=P>P@�
A�
E�
F�
J�
K�
MPRPSPZ�
_�
e�c�&K.K/K_!t`"tc%t&t22{
{
/w6272HdIdL|
M|
N|
R<U|
V|
YFc}
}
'x(x3w_!t`"tc%t&tnn#F$F-|
.|
2|
3|
5F6F>x?xH}I}LxMxUsVs]|
^|
cFFFF'n(n,d-d0d1d=F>FBFCFU!tV"tc%�&��
�
�
�
 P#P(�,�1�3P4P9�
:�
;�
?�
@�
A�
M�Q�TPUPc$F%F(|
)|
-w1wBpCpSzTzY|
_!t`"tc%r&rFF1�	2�	1�	 2�	+1�	,2�	7F8Fc1�	2�	FFFF'1�	(2�	<F>FA1�	B2�	C1�	D2�	JFKFO1�	P2�	Q1�	R2�	S1�	T2�	_!r`"rc%t&t	|

|
7282<<>s?sBsCsMnNnWl
Xl
c2<3<9x:x=s>sFnGnMw_!t`"tc%t&tF|
|
|
FF"z#z1x2x6n7n?|
UFVFc
F|
|
 F!F%F3w7w>s?sCnDnHsIsM�N�QxRxV}W}_!t`"tc%�&�
UU�
�
$U%U(�
-�
.�
2�
7�
8�
FUGUJULUU�
V�
Y�
[Z\Z_ZkZlZcZZ#w'w-F.F1w6w:w_!t`"tc%r&r
FF+1�	,2�	S1�	T2�	c1�	2�	FF2F3F51�	62�	?1�	@2�	C1�	D2�	O1�	P2�	S1�	T2�	_!r`"rcs�{���������������������������×Ǘ˗ϗӗחۗߗ���ǘ����c�?�C�g�����c�?�?�c���������ǘ�g�C��ǘ?�?������ǘ����g�C������ǘ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'��������'�'�'�'�'�'�'�'�'���������'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�'�ݙ�	��5�K�a�w�����������������������Ϛ����'�=�S�i��������������1s���������1s4p��������.v1s4p�������+y.v1s4p������(|+y.v1s4p�����%(|+y.v1s4p����"�%(|+y.v1s4p���"�%(|+y.v1s4p7m��"�%(|+y.v1s4p7m:j�"�%(|+y.v1s4p7m:j<h"�%(|+y.v1s4p7m:j<h�%(|+y.v1s4p7m:j<h��(|+y.v1s4p7m:j<h���+y.v1s4p7m:j<h����.v1s4p7m:j<h�����1s4p7m:j<h������4p7m:j<h�������7m:j<h��������:j<h���������<h������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o����������������������������������������������������������������������������o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o��o�'�'�'�'�'�'�'�'�'�'�����������������������������������������������������������������������'�'�'�'�'�'�'�'�'�'�'������������������������������������羚�������������������������������������������������������������������������<h:j7m4p1s.v����������������������<h:j7m4p1s.v���������������������������������������������������������������������_�w���������������������_�w���������������_�w������������������_�w������������������_�w���������������_�w������������������������������������������������������_�w������������������_�w������������������_�w������������������_�w������������_�w��w��w���������������_�w��w��w���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                        VVVVUUUU����������������VVU�VVU�VVU�VVU�VVU�VVU���������V�VVU�VVU�VVU�VVU�VVU�VV��������VVU�WUU�WUU�WUU�WUU�WUU���������                                                            VVVVVVUU����������������VVU�VVU�VVU�VVU�VVU�VVU���������U�VVU�VVU�VVU�VVU�VVU�VV��������VVU�VVU�VVU�WUU�WUU�WUU���������U�WUU�WUU�WUU�WUU�WUU�WU��������WUU�WUU�WUU�WUU�WUU�WUU�����VVVVUUUU����������������VWU�VVU�VVU�VVU�VVU�VVU���������U�WUU�WUU�WUU�WUU�WUU�WU��������WUU�WUU�WUU�WUU�WUU�WUU���������U�WUU�WUU�WUU�WUU�WUU�WU��������WUU�WUU�WUU�WUU�WUU�WUU���������U�WUU�WUU�WUU�WUU�WUU�WU��������WUU�WUU�WUU�WUU�WUU�WUU�                                                                                                                                                                                                                                                 � ��
 ��; ��� ��� ����ՙ[ֵ����������������������������������j���j���Z�Z�Z�V�Z�U�VeUUVeUUUUUUUUUUUVeUUUUU�V���Z���Z��������������������������������������������������������������������������Z���V���U���Ui��UY�jUYUfUUUfUUUUeY�UUUU��ZU�jje�VZ����j�j������������������������������������������������
���*���*���*�����j���j���Z��Z��Z��VeUVeUUUUUUUUV%UUUU�V���Z���Z���������������������������������������������                                                                        ����
���
��������*����������������������������                                                                �    ��
 �** �
����*�*��������������������������������                                                                                                                        ����
���
��������*����������������������������                                                                                                                �    ��
 �** �
����*�*����������������������������������*��+���>��>���7�UPUU7�]w��� ���: ���� ��������z���_� U]�             
  ����  
                 ���������?����|��_u{�_w�5|� �                                        �    ��
 �** �
����*�*��������������������������������0   �   �*  ̀
��*          ��������?, ����������U�U�u�u���� < <                                            ����
���
��������*����������������������������0   �   �   �               ��������?, ����������U���u������ <;<  ;   �   �   �  ��  ��  ��  ��  ��  ��  ��  �⨀��������������*����������������������������      3   3   3  ��  ��  ��  ��  ��  �����������8����_�?�Ww�U�_�]_����<�<  �   �   �   �   �  �  �  �  � �  � *�� ������
���*�
������������������������������                                                            ���������ꫮ�ꪺ�z���z�_�_�UUUU�VU�WVjUU�ZUu�U]UeVU]UYUUUe�U���������ꫮ�ꪺ�z���z�_�_�UUUU�VU�WVjUU�ZUu�U]UeVU]UYUUUe�U�V��������������W�W�V�W�^�W���W���_�W�^�W�^�W�^�U�zUW�������                                                                                                                           �  �� �ꬪ��������������������ZU��UU�j�uuUW]UUU]�Z�Z�j�j�տ����^�^�W�^�W�^���^U��^U�zU��UnU}U_U��_�������_�������                                                                                                                        �   ��  ꬪ ����������������꯮�U���UU��]W�ju�U]uUUU�j�Z���j�W������^�^�W�W�W�W�U���U��U���U���U}U�W�U���V������V����                                                                                                                        ����VV�VUUeUWUeU��U���������U��zUU�_UUUUUUUUUUUUUUUWUU��U���������W��UU�zUU�_UU�_UU��WU�]UU�_UU�uU]u�WU]U]W]]UU_UUUUUUU                                                                                                                        ����V�VVUUVUUU_�U����U�z]U�zuU���U��U��Wկ������W���^���^�W�z�U�z�U�{�UU�UU��UU��U��W]�UU�WUU�UuU_]UUU�UUUUWWUUUU]U] �� ��? �� �w5 �u5 pU �U  U  �  V �Y �ie ��e  j  �  �  \  T    �? �� ��? �W �w5 �u5 pU �U  U  �  Z �Y �ie ��e  Z �o �� �   �< ���� ��? P_? pu? pu= PW5 PU @U  �  @U dU& d�Y �UV ��_ ��� _�_ _�  @   =  �? �� �� �� \� \] �U TU PU  �*  `U `i `�	 �i	 he	 f� �� T�= T@= � < �   �� �� �� \� \] �U TU PU  �*  `U `i P� �� e� �� T�  �  �   <  �?  �� �� �� \� \] �U TU PU  �*  @�  Pe Yi YV P�  ��  ��  P�  P  P�  ��  �� �� T� \� \] �U TU PU  �*  P�  Pe Yi YV ��  p� �� P� TT  <� ?�  �� �� �� �] |] \� pU @U  �  @U �U eV �U �� ��� ��� �_� P  |   �  �� ��? �� �w5 �u5 pU �U  U  � @U	 @i	 `�	 `i
 `Y) ��� �* |� | < ?   � �� ��? �� �w5 �u5 pU �U  U  � @U	 @i	 @f @� �VY ��V  �  T  P?  <   � �����X��X^��]]P�UPVU@YU @�*  UU Te	 Te	 \e	�_	_�W_�� @U   T=  @=   0�� �����e	�]m	|]�\�epUe@UY  �V PU XV XV XV X�0P�W=��U=@U _  _       �? ��� ��� Y]]i]]��U�U�P�j@UU  U� U� �?�����������S�  W              U @� @� [�w_�w||��U����  �?@ �?p U|@U��PU�pU��U  �   =            �  � ��? �_� �W� ��� �U��W�\_W5�� pU �U��� |�� ��? �?  �  p  �  � �� ��? �� �w5 �u5 _U wU5 �U \�3 �U��W� \�  �� � �_� ��� � ?�? ��   �       �?  ��  �� ��_ ������� _� �U _U�]� p5 p�? ��? _�� �W? \ �  �?  �������������U�U�U�U�U�U������V�V�V�V�V�V��������         `   T   _   pU    U
  `��  p��
 T��* W��: W��* U��
 T�� \UU  U�                  �*   ��  �� ���
 ���
 ���
 ���
  ��  ��                       � �?���~$ �0  30�<�������������|������UW�UU=�UU?�W�?��� ��   0� ��<��?������?���?���=_���_�U�|UU��UU��W�?��� �� �X~UZ���V���ZYUu�Z�_XU�UZ]~}��_�~U� �UWU�U)U}U)UUV��_�%���
~UU P  T  t  T  �  P  �  �
  x�  Z��j�
�`%
 �-  ��  
�� 
 �
  �*  �*  �*  �*  �
  �  �*  `�  �� �%  �
   
   
   
  �
  �
 ��  �     �� �j	 �Z) �V) �Z* ��* ��
 ��  �? � ��� �<���?�� �� � �����?<���?���� ?��  �<<�� <� � ?��  �<<�� <��� �����<<������� �����<<����� �����  �<<�� << �����  �<��� <� �?� �����?�?��?<��� ��� � ��?<����?�303  303  �00�� �?0 000 00������ `YU�XUUUVUUUV_W�������������X_�]X]UU����  �   �   �   �   �   �   �     
   �   U  U  U  U  _  U  �                                 0�w����O���0�w���|=��   �� �� _�?���> �> ��> ��> �� p� \�  \?  \  |  �?   �   � �� ��> |���]� �U� �W�  _�  |<  p>  p  p  p  �  �   <       �   X   V  �U  ��  �u  ��  �U   �   V   �                            �*  V��UUU)UUU��w}���ݝ��}���ݝ��ݕUUU���� �*  �*  �*  �*  �*  �*  �*   �:  ������e*�ٮ/��f�f}�f�j��Y�=��j���  � ����
 Z) �� ��� �  �  �  �  & �
 h � ����
 Z) �����  � (� �� �% �
         ����������>�>���<T P�W�_�>����T�<  P<T����>�>� P<T����>�>���������?, ����������U�U�u�u���� < <���������?����|��_u{�_w�5|� �    ((���������*�
�?�??���� <<�� < ?< ��� <?<�  <�<���< < �< ��< <<��< ?�??�� � ������������������������������                                                                                                                                                               ���ة��  ��� ��� � ��� � �ߍ& ��" t ����9 ��: �� � �9����: ��� <�X � u�L �H�Z�� �
0)8�
�� �� �� �
08�
�� �� �� �
0	8�
�� �� �� � �Λ  ��z�(h@H�h@                                                                                                                                                                                                                                                                                                                                                                  ����  �� ��L �� ����� �
 \��� ��� �  π ����� �ߍ& �  �� <�  � ��덉 �   ����Ή �0��  \� � �� �� ;���� �  g� n� <����  \� \� \�  ��L �� �� ���� ��'�� �� �Lj��� �Lj��� �Lj� �Lj���'�� �� �Lj��� (�Lj��� (�Lj� 5�Lj���#�� �� ��_�� B��V�� (��M N��H��#�� �� ��8�� ��/�� `��& 5��!�� �� ���� ���� `�� 5� <���  ^� �� �� +� �� �� ���L�� �� �� �� �� �� ���H�Z�� �� �ɀ�� �ˀ�� @� �� �� �� ��֮  ���   ��� � �� �� �� �� ����  \�������� ���� `� +� ��Ls���� 3�Ls���� l� �ɀN��� l� �ˀB��� l� @΀6��� ��Ls���� `� 3Ȁ ��L,��� u���}� u���~� u�z�h`��� �� �ɀ���� �� �ˀ���� �� @΀���� �ǀ���� 3Ȁ���� 3� `� +� ��Ls���� ��Ls���� 3�Ls�L��H��� ��� �� �� �; �f �< �g  (�h`H�< 8��g �; �f ��� ���  �h`H� ��  (ũ��� h`xHڭ� 
��O��9 �O�m� �:  H��hX`H�Z�� �� �� �� �g ���7 ����8 �f �9�� �� ���� 7�� �� -� �7�9 i�9 �: i �: �΋ �� � �ȭ� �� �Ό �� � Шz�h`H�� ����  j��? �? � � +� ��h`��? �� i�� �d08�d�� �� 8�d�� �� �� ͥ $�� �� ͥ �� �� ͥ �� �� ͥ ��  �耣H�? �= �� �� �� ���� �� m�L���� 7�L�� D�L������ ������������ �L������ ������ q��?���������� ����������LFƀ��� ��LV���LP���LF� ��� �� �� �� �@ �>  ��� �= i�= �,L8�h`H�Z�� 8�
��i��9 �i��: �� 8�
��9�7 ȱ9�8 �� 
��7�9 ȱ7�: �� 
��9�� ȱ9�� �> ���� ����� �= ��-� ���� i�� �� i �� �΍ �⭰ �� �Ύ �� ��z�h`H�� ��
������� ��X� �� �G�; ��3 ӭ� � � ���;  �ĭ� � +� �� �� ��E��  \� ;�h` �ĩ��  \��Щ�� ���E�� � �� �$ -ɭ; �� ���;  � �� +� �� �� \������ ��H�� ��
�����
�� ��L��� �� �0K�
G�; �G �ѭ� � �4 �� �ҭ� ���;  � �� �ĭ� � +� �� �� ��`��  \�h`��� �� �ҭ� ��� �� �� �� �� �� ��5��  \���� �� �0.�
*�; �* -� ���;  � �� +� �� ���5��  \�L�ȩ�� �� -� � �� �� �� ���%��  \�L��H������7 ����8 �; i��7� �h`�< i�<  <� � �� +� �� �� ���H�< �08��� �� �� h`H�< �208�2�� �� �� h`H�Z��� �� ��
�����
�� ��L|ʭ� �0��� ��
�� �� � �R�� ���� �� �� ��  �ĭ< 8��<  �� +� �� �� �� �� �� �魝 i��  \�< �
0͵ 0�����  m˭� � �6 �ĭ< i�<  �� +� �� �� �� �� �� E쭝 �0�8���  \������� � �� z�h`�� � ��� � �L+˭� �0��� ��
�� � �� �< ͵ 0} �ĭ< 8��<  �� +� �� �� �� �� �魝 i��  \��ĩp�< �� �� ������7 ����8 �; i��7� ���� z�hL�� �ĭ� �
�� �� ����  ��Lnʩ�� �< �p� �ĭ< i�<  �� +� �� E� �� �� �� �魝 �0�8���  \���H�Z��� �< i����7 ����8 ��� �� �
��; ��; i��7� ��Β �� � ���Α �� � ��z�h`�8�� � �č< �� �
�� �� ����  �ĩ �� �� ��H�Z��� �
�� �� ��
�����
�� ��Lͭ� � �L�̩ �� �; ���; �� �x �ͭ� ��V�� ���
� �� �� �� ��V ���; �< 8��< ͵ 0L �� �� �� �� �� �� �� E�< �0#�E��  \�L̭� ������� ���  ��z�h`��� �� �ޭ� ��ש�� �; ���; �� 0� ���; �< i�<  �� �� �� �� �� �� E�0��  \� �̀��@�� � ��� � �=� �� �< ͵ 00�; ��) ���; �< 8��<  �� �� �� �� �� �� �� \��í< �p6��� �; ��# ���; �< i�<  �� �� �� �� �� \��ʩ�� � -ɩ �� ��  �ĩ ��  ��L��H�Z�< i����7 ����8 �; 8���7� �z�h`��� �� ��H�Z��� �< i����7 ����8 ��� �; ��7� ��Β �� � ���Α �� � �π" N�8��< �	 �č<  �ĩ �� �� � �� z�h`H��� �� ��
������� �� ��L Ϝ� �� � �L1� �ϭ� ��L ϩ�� � �� �� ���
� �� �� �< ͵ 0ͭ; �3 ���; �< 8��<  �� �� �� �� �� �� �뭝 i��  \�Lq� �ĭ� ��;�< 8��< �05͵ 0: �� �� �� �� �� �� �� �� �ϭ� i��  \������� h`��� �� ���� �� ����� �; �1 ���; �< i�<  �� �� �� �� �� �� E� Щ5��  \����� ��9 �ĭ< i�<  �� �� �� �� E� �� �� �� Э� �0�8���  \���L �H�Z�� �0.��� �< i����7 ����8 �; i��7� ��Α �� � ��z�h`��� �� ��H�Z��� �< i����7 ����8 ��� �; i��7� ��Β �� � ���Α �� � �̀$��  ��8��< �	 �č<  �ĩ �� �� z�h`��� �< i����7 ����8 �; i��7� ��Β �� � �ܩ��� �ũ�� �� ��H�Z� ��� ��� �� � �K� �� �< ͵ 0z� �� �; �4 ���; �< 8��<  �� �� �� �� �� �� �魝 i��  \����:�< ͵ 02 �ĭ< 8��<  �� �� �� �� �� �� �� �魝 i��  \��ƭ< �pk��� �; �( ���; �< i�<  �� �� �� �� ��5��  \��ŭ< �p0 �ĭ< i�<  �� �� �� �� �� �魝 �0�8���  \��� -ɩ �� ��  �ĩ��  ��z�h`H�Z��� �< i����7 ����8 �; i��7� �ȱ7� �Β �� � ��Ӎ�  ��8��< �	 �č<  ��z�h`��� ��  �ɀ�H�Z��� �< i����7 ����8 �; i��7� �Β �� � ��ڊ8��< �	 �č<  ��z�h`��� ��  �ɀ�H�Z�< i����7 ����8 �; i��7� �� �� ���� �0��� �< i����7 ����8 �; i��7� ��Β �� � ��z�h`�8� �č<  �Ā�H�Z �ĭ< i����7 ����8 �; 8���7� ���� �I�< i����7 ����8 �7� ���� �)�< i����7 ����8 �7� �	�< 8��< � ��  +� ��z�h`���� �� � �����  �� �� +� �� �� \� �ĭ< 8��<  <� �� +� �� �� \� �  g� n� �ĭ< i�< ��  �� +� �� �� ꩀ��  \�< ɖ0� <� +� � ����� ����  \�Β �� � ��  ��� �
0	8�
�� �� �� � �L �� �� ���� L � wթ�� �d �0M�� �* �ԭ� � � ?Հ �ԭ� �e �Z ��#��  (��Z `�Z ��$��  (��Z �� �Z ��,�d �t�e ��� �ӭ� ���;�� � �4�d 8��; )�d i�; 0�e 8��< �e i�< 0��� L��`H�� � �8�� � �1�d 8��X &i�X 0�e 8�	�Y ��� �� i�� � �h`H�$�� ��� ��� �d �f �� ��e 8��e �g  (��� h`��� ��H��� ��� �d �f �e �g �#��  �h`H�� ��0�{ �0+�y �| �z �� �" ح� ��5 ׭y �{ �z �| h`��� ���� ��  �֭y �{ �z �| �� �� �ک�� �����H�� ��0�} �0+�y �~ �z �� �" ح� ��5 ׭y �} �z �~ h`��� ���� ��  �֭y �} �z �~ �� �� �ک�� �����H�� ��0� �0+�y �� �z �� �" ح� ��5 ׭y � �z �� h`��� ���� ��  �֭y � �z �� �� �� �ک�� �����H���  ة�� �� ��z 8��g �z  (�� h`��� ��H ة�� ���  hحy �%~�f �z �q-�x �9� �	�z i
�z �z �g �y �f ���  (��x �>�^�,�y �2�z � �x �+�x �&��	�z i�z �y �f �z �g � ��  (��x h`� �x ���y �f �� �z �g ���  (ŀޭx � � ��y �y �f �z �g ���  (��x ���x �����y �y �f �z �g � ��  (��x ��H��� ��� �z �g �y �f  �h`H�� � �?�y 8��X 4�y i�X 0)�z 8�	�Y �z i�Y 0��� �� i�� � �h`�� ���+�; �y #i�y 0�< 8��z i�z 0��� L��`�t �0\�r �u �s �� � � �� �٭� ��&��� � ���� ��  ڭ� �� �s �u �� ��� �u �s  q٭r �t �s �u `�,�t ��H�v �0]�r �w �s �� � � �� �٭� ��&��� � ���� ��  ڭ� �� �s �w �� ��� �w �s  q٭r �v �s �w h`�,�v ��H��� ��� �r �f �s �g ��� ���  (Ŝ� h`�� ���4�r 8��; )�r i�; 0�s 8��< �s i�< 0��� L��`H�� � �:�r 8��X /�r i�X 0$�s 8�	�Y �s i�Y 0��� �� i�� h`H��� ��� �r �f �s �g ���  ŭ� �
�s 8��s �g ��� ���  (��� h`H�� �E�i �0@�h �n �m �� �7 �ۭ� ����� � ��!�� �n �m  #ܭh �i �m �n h`��� ���� ��  �ۭh �i �m �n �� �� ��H�� �:�j �05�h �o �m �� �, �ۭ� ����� ��� �o �m  #ܭh �j h`��� ���� ��  �ۭh �j �m �o �� �� ��H�� �@�k �0;�h �p �m �� �2 �ۭ� ����� �!�� �p �m  #ܭh �k �m �p h`��� ���� ��  �ۭh �k �m �p �� �� ��H�� � �:�h 8��X /�h i�X 0$�m 8�	�Y �m i
�Y 0��� �� i�� h`H �ܩ�� ��� �� ��m 8��g �m  (��� h` �ܩ�� �,�h �� �� �ܭh �04�� ��1�� ��'� �� ��� ��� �h �f �m �g ���  (��� `�h �� � �(��� ��� �h �f �m �g ��� ���  (��� ���h ��H�h �f �m �g ��� ��� ���  �h`�� ���4�h 8��; )�h i�; 0�m 8��< �m i
�< 0��� L��`H�Z�� 8�
�����9 轷��: �� 8�
��9�7 ȱ9�8 �� 
��7�9 ȱ7�: �� 

��9�c�4ͤ �*ȱ9�� ȱ9�g ȱ9�� ��� �= i�f � ��  (ŀ�� ������ ��� �� 8�
�����9 轷��: �� 8�
��9�7 ȱ9�8 �� 
��7�9 ȱ7�: �� 

��9�c�L�� �P�� �K�� �F�� �A�� �<�� �7�� �2�� �-ͤ �(ȱ9�� ȱ9�g ȱ9�� �= �0�f  (ũ �� z�h`�� ��H �ޭ� ��L�ޭQ �0- ߩ�� �Q �R i����9 ����: �Q i��9� �	�0��� �8�R i����9 ����: �Q i��9� ��R i�R �R �g �Q �f  (�h`�R i����9 ����: �Q i��9� ��R i�R �ĭR i�R ���� ���4�Q 8��; )�Q i�; 0�R 8��< �R i�< 0��� L��`H��� ��� �Q �f �R �g �'��  �h` �߭S �0 �� %�� � � k��\�� � �]��,�S ���T � �� �� �?�T �F0@� �� �T �P8��T �g �	8��T �g �S �f �(�� ��� ���  (�`� ����T ɇ��� �T i�T �g �S �f �)�� ��� ���  (ŀƭ� ���9�S 8��; .�S i�; 0#�T 8��< �T i
�< 0��� ���� L��`H�� � �<�S 8��X 1i�X 0)�T 8��Y �T i�Y 0��� � ��� i�� h`H��� ��� �S �f �)�� �� ��T 8��g �T  (��� h`H�S �f �T �g ��� ��� �(��  �h`H�K �
���K �C �f �K �g ��� ���  ŭC i�f  ŭC ��X�-�C LR� ���� ��� ��� �� � �9� �� �C �f �K 8��K �g  (ũ�� �C i�f  (ŭK �<��� h`��� �C �f �K i�K �g ���  (ũ�� �C i�f  (ŭK ɇ0ǩ �� ��H�� ���,�C �A �K �I  �᭳ ���� � � �ĭ< 8��<  ��h` �ĭ< i�<  �Ā�H�A 8��; M�A i�; 0B�I 8��< ��< 8��< �j�I 8��< ��< 8��< �T�I 8��< ��< 8��< �>� �� h`�I 8��< ��*�I 8��< ��< i�< ��I 8��< �˭< i�< ��� � �� ��H�� ����� ��� �
��� ��� �U �f �V i�V �g ���  (ŭ� ����� �U i�f  (�h`H�U �A �V �I  �᭳ ��	�< i�< h`H�H ��,�H L��� ���L�� ,��� �� �P ��� �H �A �P �I  �᭳ ��L��H �f �P �g �� �������� ���1��  (ũ2�� ���� ���  (ũ�� �H i�f  (�h`�P ɠ� ,��� ���� ��� �P i�P �g �H �f �� ���������  (ũ�� ��� ���1��  (ũ2�� �H i�f  (ŭ� ���� �ĭH �A �P �I  �᭳ ���< i�< Ɍ ��L���� hL��H�H �f �P 8��g ��� �� ���������  ŭH i�f  �h`�� ����H�C �f �K �g ��� ��  �h`�G �f �O �g ��� ���  ŭf i�f  ũ�� �G �0
�� ���L%�-�G � �O � �� �O�� ���I�G �A �� �O �I  �᭳ ��0� �� �G �f �O �g ��� ���  (ũ�� �G i�f  (�`���� �� ��� �ĭO �0�8��O �g �G �f ��� ���  (ũ�� �G i�f  (ŭ� ���� � Ю�< 8��< �< �0 ��L$��� L��H�� ���Lb� ���� �� �N �� � �Ln�F �4���N ���� �y �0��y � ��y �f �N �g ���  (��y Lb� �� �� �0�F  �ξ �� �F �f �N �g ��� ���  (ũ�� �f i�f �0 (�� �� � � ��� �� �� �0ξ �� � ���� h`���� �F ���F �0��� �F �,N�� �0 ��F � �� �F �f �N �g ��� ���  (ũ�� �f i�f  (�� �� �К� �� ���� ��� �� �� ��� �� � Lb�H��� ��� �F �f �N �g  ŭf i�f  �h`H�� ���& �ĭF �A �N �I  �᭳ ���� � ��;  ��h`�; �0 �� ���F ���;  �Ā�H�� �0:�� ���3� �����  �ĩ��  �ĩ ��  \� �ĩ��  �� \� ����  �� ��h`H�Z�� � ��� � �L��� ��� �X �f �Y �g  ŭ� � �-�� �� � �Z�X i�X �Y i�Y �F� �.�� �� ��6�X i�X �Y i�Y �"�(�/�� �� ���X i�X �Y i�Y  ��� z�h`�%�0�� �� ���X i�X �Y i�Y �0�� �ͩ �� L��< 8��Y �; i�X ��H�Y i����7 ����8 �X i��7� �6���7 ����8 �7� �#�< i�Y 0�X �,�X �f �Y �g  (�h`� �� ��H�� ���� ��6�� �Z�/�/���� ��"�� �Z����E�� ��.�� ���� �Z�h`�� i�� �
L��� 8�
�� �� ��� � �٭� �P�Ҁ����� ���� �о�� �Zз���� �Ю�� �Z�L6��� � �����  \�; �,�D ���; �� ���r�< �����r�< �  �� +� �� ���� �	���� ����  \�� ���  �����  \�L �H�� � ��=�� �  �h`�	�f �
�g �X�� ��� ���  (ũ�f ��g ��� ��� �Y��  (ũ�f ��g � �� ���  ŭ� ���E�� � �?�� ��Ρ �� �� �� ��f ��g ��� ��� �,�� �� � � (�μ �f ��`��� L�ӭ� ��I�� ��$���< Ɍ06��� L�Ӏ,�< �}0%��� L�ӭ� ���� �#0�< ɇ0��� L��`���� ��Ȁb�< �q0��� L����'�� ������< ɀ0ɩ�� L�ӭ� �<0��(���� ������L�ꭟ �������L��< Ɍ0���� L�ө�� �< ����9 ����: �; i��9� ��Β �� � �$�ڍ� �� ������ �� � � �� ��`�� ����歞 ��	�� ���J��� �< ����9 ����: �; 8���9� ��Ή �� � ��ڍ�  �ﭞ ������ q� ��`�� ������ ��
�����	�� ���R��� �< i����9 ����: �; 8��W ���� �9� �Ș�W Β �� � ��Α �� � ��Í�  �� N�`��� �< 8�����9 ����: �; 8��W ��9� �'��� Ș�W �9� �Α �� � ��λ �� � �ʀ� r�`�< �20�� ����������|�	�����` �ĭ� � ��; ��< i�< �;  �ĩ�� L�ӭ� ����0�` �ĭ< i�< ���  ��L�ӭ< �20#�� �0���������������	�=��?�` �� �ĩ�� L�ӭ� ɀ�ɰ����ɫ�ɛ�	�[����` }���� ���	ɀ���` �ĭ< i
�<  �� �� }�證 ��P����  ���;  �� \� \��� ��� �; �3 ���;  �� ��� � \�λ �� � �ۭ� �08��� `� �� �� <� � �� �� ��� �����  \�λ �� � �ڀ�H�Z� �� �� ��� ���  �ĭ; �{�;  � �� +� �� ��� �����  \�Β �� � �ͩ�� �< i����7 ����8 �; i��7� Ш�; 8���7� Л���� �� �08��� �� z�h`� �� �� �� � �� �� ��� �����  \�Β �� � �ک�� �< i����7 ����8 �; i��7� е�; 8���7� ШL��Hɪ�ɠ�h` ���H�� ɠ�
ɨ�ɪ�h` ���H�� �@�
�	��)�h` ���H�� �� �	�� i�� �W 8��? 0� ��� � ��� m� �� �0�� � ��� m� �� ��� � ��� m� �� �
�� m� �� ��  <� �� +� �� �� �� i�� � �h`H�Z�9 �@�: � � � �9����: ���z�h`�Z�� � ����� ���� ��z�`H�Z g� n���)��&  ���f �M�g ��� ��� ��� � ��  (ũ���  (Ů   ����������� ��  (ũ���  +� �ĩߍ&  ^� ��z�h`Hڭ  �����h`Hڪ�J�




�� ��)� �& �h`H�Z ��
��M��� �M�i@�� �č� �@�� �� � � ������(���� i0�� �� i �� �� i(�� �� i �� �   ������ � �� ��  \���е�ߍ& z�h`��� ��H�Z� ���Q� ���.� � g�� � � �  ^� � n�� � � �  ��� � �	 � $�� � � � �� ���.�( � g� n��! �" � � � �  ��( �( �# � ��(z�h`� �� ȱ� ȱ�	 ȱ�
 ȱ� )
��/�� �/�� Ȍ � � �	 � �'� �1� ȱ1� � �� � �� ��Ȍ � ��`� ��! ȱ�" ȱ�# ȱ�$ ȱ�% )
��/��& �/��' Ȍ �( �) �# � �#� �  g� n�� � � � � � � � `� �� ȱ� ȱ� ȱ� ȱ� )
��/�� �/�� Ȍ � � � � �'� �3� ȱ3� � �� � �� ��Ȍ � ��`H�Z�
 )?	@�+ �
 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �/ �� �/ z�h`H�Z� )?	@�+ � 4��-+ �+ � ��� )@��J��+ �+ Ȍ ����� � � �+ �0 �� �0 z�h`H�Z�$ )?	@�+ �$ 4��-+ �+ �) �&��% )@��J��+ �+ Ȍ) �&����) �% �) �+ � � �/ �0 z�h`� �/ `� �0 `H�Z�* z�h`� � �  g� n�� � � � � � � � �/ �0 �ߍ& `

�����1 ȹ���2 ȹ���3 ȹ���4 � �1� �3� ȱ1� �3� � � �� �  $� �� ^� ���� `H�Z
���� ���  � ��*  �� ���� z�h` �� ��� ��� ��� ��� ��� ��� ��� ���  �� ��� ��� ��� ��� �� q�� ��� �� j�� q��  �� q�� T��    _�� j�� q�� j�� �� ��� �� j�� ��� ��� ���  
�� �
�� ��� ��� �� ��� ��� ���    ���  ��    ��  ��    �'�T'��'�T'��'��'��'�}'�T'�  '�T'�.'�T'�'� �'��'�T'� �'��'��'�  '��'�T'�   }'��'��'��'� �'�@'� �'��'�}'�@'�T'�  
'�T
'�.'�'� �'�T'��'�T'�   �'�  '�    �'�  '�    �� ��� ��� ��� ��� ��� ��� ��� ���  �� ��� ��� ��� ��� �� q�� ��� �� j�� q��  �� q�� T��    _�� j�� q�� j�� �� ��� �� j�� ��� ��� ���  
�� �
�� ��� ��� �� ��� ��� ���    ���  ��    ��  ��    �'�T'��'�T'��'��'��'�}'�T'�  '�T'�.'�T'�'� �'��'�T'� �'��'��'�  '��'�T'�   }'��'��'��'� �'�@'� �'��'�}'�@'�T'�  
'�T
'�.'�'� �'�T'��'�T'�   �'�  '�    �'�  '�    ��� ��� _�� ��� �� ��� ��� ��  �� �� �� w�� ��� ���    �� ���  �� ��� ��� ��� ��� ��� ��� �� �� w�� ��� _�� _�� j�� j�� ��� �� �� w�� ��� _�� _�� j	�� ��� $�� ��� d�� w�� �� d�� q�� ��� ��  �� ��   @����� ���    O�� G�� O�� O�� _�� O�� O�� ;�� O�� _��    O��    w��    ��� ��� ��� ��� w�� j�� _�� Y�� ��� ��� ��� ��� �� q�� d�� _��    ��� ��� ��� ��� �� q�� d�� _�� ��� ��� ��� ��� w�� j�� _�� Y��   @��}�����@��    w� 2�    w�� _�� O�� ;�� /�� '�� ��    O�� w��    _�� d�� d�� j�� j�� q�� q�� w��    �� ��� ��� ��� ��� ���    O�� ?��    ��� ��� ��� ��� ��� O��    w�� ;�� _�� ,�� #�� �� �� �� w�� _�� O��    �� �� ��� ��� ��� ��� d�� ��� w�� ��� ��� ��� �� �� �   	 �		� �

		�
	 ��
		 ����������������@�  ��  /����/��������������  !�����!�����{����{���  �C��K�  ��  S�  ��  ��C�P�{��������  R�[�g�n���������   @�?���O���_�����ߵ/��϶�o����_���߸���/���ǹߧ�#�C���úͻ�����M�����5�}�Ž���2!""C�K�[�k�{�����Ӿ2b�a�a�a�a�a�abb$b@b�b�bchc@yJyxczy�c8d�d�d�B~��2n��"!#W0�C� 	 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____H��� ���  (�h`� ��L ��  ��L�� ��L �                                                                                                                 S� ���