                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �����������������               �               �               �          �    �          �    �      �  �    �      � ��    �      � ��    �      ��?��    �      ����    �      �S���    �      �W���    �      ����  � �      ����� �� �      ��+�� q�      �s)���T\�      sq=���T\�      �}���0W�      �����LW�      s�����U�    ��]����W�    ?��W�_W�   ��5���~UOW5�   0u5��^OU\5�   Lq�]��^;��5�   \}]��^E;}\?�  ��_W� �^E�Wq��  �_��U�^Q;Uq��  �T5�TU�^Q;Uq��  �T5�TU�^�;U���  �T55UU�_��T�}�  �T54UUU��T��  �T�4U����T���  �TM��WU�������  �TOM�_������  �T�5u|��ϺSW�  ����p����OW�  �_���_��OW�  �Tӫ��U��;�_�  �TS�z�_U���_\�  ��S�_�UU����_�  �_SU]�UU���_|�  �TSU]�UU��;U��  � MU]�UU��;U\�   �OU��UU��;U\�   LMU]�U��NU\�   �OU]�U��NU\�   S=U]�U��NU\�  �_7U��U���NU\�  �_7U�����OU\�  ��5US����SW� ���5�T����SW� �����T�w�o_SW� ���������_SW� ������w�o_SW� ����7�����TW� ����=�w�o�TW�����7�����TW������=�����T�U������6����� �U���~��;�������W���~��? �ױ����^���������q�?��z����U����ձ� pS�����W�ݪ��q� \S�������]����fWs�����:p]��UǙ�s�ÿ�W?pW�W�f�\�ÿ�WpWlWǙ�W�ÿ�}pW�W�f�W�����pgWǙ�^�c�����Wg�� �s�{�pgW5��? ����p�\�g   ����pg\�   ����? \�\g6   ���  \�f\U�9   ���  \ř\Ul6   ���  \�f\U�9   ���  \řpUl6   ���  \�fpU��   ���   \řpUq�   ���   W�fpU��   ���   WřpUq�   ��?   Wqfp���   ��?   �����   ��?  �ofϵ[  ��?  �m�� ���9  ��  �m\� ����;  ��  s+WU����7  ��  �W]�TUř;  �� �T�Uw�T�f�  �� ���Uw��W���  �� ��U]�TUqv�  ��  �U�UU��ŝ�  ��   �W����m�  ��   wי���� �?   w�fӵ�gf �?   {������ �?   w{lf��gf �  ���� LU�� �  �UUl� LUUlf �  �U�� LUU�� �  �Ug� LUUlf �  pU�� LU���9 �  �_�� �_W\g6 �  p]�� L]���9 �  �W�_� �WU�W7 �  pU�y� LU���� �  �W��� �_W��� �  \�ŵ� L]��� �  ����� �WU��� �  \U�]� LUU�_��  WU��? LUUq�w�  WU��9 LUU����  WUqf6 LUU�f~�  WU��9 LUUř��  WUqf6 0UU�ff� �UU��9 0UUř�� �UUqf6 0UU�ff� �UU��9 0UUř�� �UUlf6 0UU�ff6� pUU��9 0UU��9� pUUlf6 0UUgf6� pUU��9 0UU���� pUUlf6 0UUg��� \U��9 0UU���� \Ug�6 0UUg��� ��W? 0UU���� Sq��� 0��Ul���T|۽�0S�U�����{��gf0S�U����0�����:�T������0{�gf�:�T������?����:�T���v�WU�gf��:�T|�����  �����:�T\qf�����gf���:��W���v�_UU�����SUg���_�_u�����TUř�����U_ժ��:0UUqf����w�^ժ��0  �٪���w�^ժ�����o�������^����WUU����o�w�^���  W�ի�������� �UW}U��  ���    ��U{ժ  �       ��{��  �       �U{�:   �       �U{�   �       �U��    �       ��     �               �               �               �               �               �               ������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���                (  (                  �               �                  0���              0l�*              0k��              �j��             ��j��             ��j�����           ��j��UUU         �K�j��UUU         �K�j����V5         ���j����X5         ���j����X5          ��j-��]�V5          ��j���}]U5          ��j���uU5          ��j��u��5           �j���]U5       �����j��u��7       <  �j��UUU5      �3  �j�����?      �� �j�����      ��_U�j��         \wUUU�j��         \w����j-��         �� ��j���         ������j��         ������j��         ������j�� ��?     ������j��  �      �����j�� WU�      �����j�� ��?          �j��  _5         ��j�� ���         ��j��           ��j-�� WUU       �K�j��� ���       �K�j��  �U       ���j��  �U       ���j��  �U        ��j��  �U        ��j��  �W5        ��j��?  �W5        ��j��?  �W�    000  �j��� �W�    ���  �j  0  _�    ���  �j  0  _U   ���  ����� 0  _U   ���     ��?  _U  ���ު�   �U5  |U ����     �U5  |U5 ������������U5  |U5 �\wuu��]UUU�U5  |U� �������^UUU�U5  �U� �������^UUU��?  �U�  ������_UUUժ:  �U�   ����_UUUժ:  �W�   �?pU�������:  �W�     |U���ݝ�:  �W�     _UW��ݝ��  �W�     WUW�����    �W�     _���������? �U�     |��j @���? �U�     ����������? p�W     �{]� C��? p\     �{]� C��? p�\     ���������? p|      ������:   p��   ��������:� p]5     W���U���U= �]5     \Uo�{U�k�W� �u�     pU��zU�^U�w�   �*�Ֆ�zU��VzU w�   0������U��Z�U�w�   ���o������Z�W�u�   ���[�*���j�^�]�   �?�V�*U���Uz|]�     �U��JU��V�_W5     l���JU���V���U5    �[���JU���Z��uU    �V���JU���jU�]U    �U���RU���jU�_U    kU���RU����U�^U   �ZUꫪRU����VUz�    �V����RU���ZU��    �U����TU���ZU�7    kU����TU���jU�>   �ZU����TU����UU:   �����������������  ������UUUUU������  \UU��WU�W�UU��UUU  \UU�W�WW�U_UUUU  \UUUu5\W��puUUUU  \UUU�5\W��p�UUUU ��UUu�WW�U_uUU����_UUUUW�UUUUU�����UUUUW�UUUU���7������������������7������������������������������������sW_���������������U_\U���������������WU\U��������������?\Up� �������������p� �? ������������� �?     �����������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ������������+���+����������������������*������������+���+����������������������*������������+���+����������������������*������������+���+
���������������������*������������+� �+� ��������������������*������������+
�?̪"��������������������*������������+����������������������*������������ ����
 ������������������*�����������
�l��3 ��������������������*������������!k��ê�?������������������*�����������r"[�T���������������������*�������������Y�Tآ�
?������������������*����������
��Z�T��  ������������������*�����������'�iE�밪�������������������*�����������'�jU��  �������������������*�����������?�iU�?說������������������*���������*k?�jU�?� ������������������*����������Z��iUj=���������������������*����������ZU�jUj5:0 ������������������*����������VUWgUj�:��������������������*����������VUWkU�j�?�? �����������������*����������UUW'P�j�0�������������������*����������UU_�����<�������������������*��������*kU���[����������������������*��������*kU��_]W����*�����ꫪ���������*��������*�Zժ^�W�:5��+�����ꨪ���������*���������j���z]׊���+�����:�����������*���������Z���ꭷ�[���������>�����������*���������V��Ϋ_��o�������������������*���������Ve�����W�
����������������/���������Ve��ê:<��T��*����-�����������/���������Ue���?��P�� ���^�����������/���������Ue��?�����������������������/���������UY �����T�* ��������������/��������ʧX (����U ����z5�����������/��������ʫV (�����UA���^M�����������/��������ʫV ������W����WM������������/��������ʫU �����_T���US������������/���������nU�������Tq��W�T������������/��������*z��������S��U5U������������.��������*x��?�����\wwUUMU������������.���������諪>����:|w_UUSU������������.������������>�������UU�QU������������.������������� � ���}UU�QU������������.���������:����� ȫ _UէQU�����������-�������������;� �/�UU��QU�����������^-���������:���?�� ��_UU��Q�����������_-������������� � ���U���Q�����������^-���������_}� 8 ���W���Q������������^-�������: �WW�0   pU߫��Q������������^,������� ���U   TU����Q������������,�������0?�p]U	  � WU����Q����������z�,��������7�0LU�    W���������������z�/�������<C5�0T  �կ���������������z��+�������� 0@,  ��������������몮�z��*�������    ��   �     ��������^�:�� ������� S             ����������^�:�������� S�            �����������^�:��?������� S�?         �������������^�:�?������� SU�>          ��꿪�����������?������� SU�/       ������������������?������� SU���        ��������������
��?������� SU���       ��������磌�ժ����?������"�TU���     ���������ꪫ�ժ����?������$�TU��       ���������k�W������?������$�TQ�       ���������W��.����?������$�TQ�        ���������W�������?������$�TQ�        ������ꫫW�������;������$�TQ5          ������ꪫ�������:������$�TQ"*       ������Z���������:������$�TQ ��*       "�����V��
�꿪��.������$�TPŪ�*       �����W����뿪��+������$�TPŪ�"        ������W�+��￾��-������$�TPŪ�       �����z�W�����￻�{5������$�TP�
�    �
 ����z�����������������$�TPŪ*      ��ȫ��z�����ﯺ��������$�TPŪ*     �*����z������﫺n��ꪪ��$�TPŪ
    �������z�����类^��ꪪ��$�TPŪ"      ��*����z��������^�>�ꪪ��$�TT��*      ���⪫�:�.����^�*�ꪪ��d�TT���    ( ��"�Z���¯�￺�*�ꪪ��$�TT�*
   > ���U�����￺���*������$�TT��* � �  ���U���￺���*������d�TT�� �� � ���U?������ﻺ��Ϋ*������$�TT��
 �> � ��������ﻺ�����.������$�TT�� �: �/ ��� �������z�5���?������d�TT�� �� � ���  /������z����?�./���� ST�* ��������� ��������z� ���?莏����US�*
������ �� ��������^� ���?�.����� S�* �����  ���������������?������US��"������> ����������찪��:Ȯ���� SŪ����:��
< ����������謪��0�������USŪ
���?��*��������꯾�뫪��>Ȏ类�US��"��#2���+�*�����꫺�������� ��类� S�� ���>�� ���������5������?�����*TS�����30��*Ȫ�������ﺺ�������/�����*U[�����;�����*��������j� ����� ����* [������� * �����������Z� �����*�>����*T[�
��8����*����꯫�W������� �>���?U[�����: �*�¿���ꫪ�W�����/�?����* [�����?�� ������ꪪ�W쬪����/�? ��?"T[�����?���
�����ꪪ��꿎�?? ������*U����������������������꯺��*�¿�?"���* ��?���*������諭����"�������ø* *��������������磌�:�?몮�3�*��»�:`�
����>(����������������� ��3�����
�
ÿ���
 �*�������ڪ갪�着����*      P��    �� ��������� ﰪ         ������
�ʏ������������������찪��������*������V�������������������>쬪��������*����������*��������������쫪��������*��������?������������������ �����������*������UU���*�������������� �����������*�����:U������������������������������*�����:������������������� ������������*������������������������ ������������*������eU������������������������������*�����WUeV�������������k��갪�����������*�����UUef�������������[��ꬪ�����������*����ꥪYf�������������W��ꫪ�����������*����z	@�e������������W����������������*����^RU�Y�������������W����������������*����^UU�Y������꿮����W����������������*����WUUVU������ꫮ�ꫪ����������������*����WUUUU������ꪮ��������������������*���������������ꪮ��������������������*���������������ꪮ��������������������*���������������ꪮ[�������������������*���������������ꪮW�������������������*���������������ꪮW���ê���������������*���������������ꪭW�������������������*����������������j�W������������
�
�
��*����������������V�W� ������������������*����������������U�W  ������������������*����������������U�  ������������������*����������������U� 𪪪��������
�
�
��*���������������zU� �������������������*������������j��zU���������������������*������������Z��z�𪪪����������������*������������U��z ��������������
�
�
��*�����������zU����ë�������������������*�����������zU�������������������������*�����������zU�������������������������*�����������zU�� �����������������������*�����������zU�: � ���������������������*�����������zU� ,��*�*���* 
���*��� *�*�����������zU� ���**����������������(�*�����������zU? ��(�**��������**�����(�*�����������zU ����**��"������**�����(�*�����������z  ����*�������
�( *��� *�*�����������z   ��(�**���������**�����*�*�����������:  �����**���������**����(*�*�����������:  ��*��**���������**����(*�*�����������: ���� �*�*�������(**�
�((�*�����������: ��������������������������*�����������:���������������������������*�����������:���������������������������*���������������������������������������*                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����  �������8��:�꣎�>���
�����>��:�㠪�㪪���������   j��iUUSUU�SU���������������������������������������䪪��    �     �
�    h	h    J$X    B�Z	    FPb)   �E��   �EP�  ��`�  �`�  �X� (�F V�* d`� JY�UU �*R�UV���UUVU��     �        ��
       ���
      (h%      h�Z�    �
�UU
    �
�UU)    �@aUU&     XUU&   � UVU�V �*@UU�R	  PI�UU)P)�
T�UU
@�� a hU� �
P	�ZU�j������UUUU���;  0;  ��  33 33 �� ���*���*��������� �� ������ �������������������������������ϫ������ϫ������������������������      ��
U *U�
*(nU�*jf(nU�*jf(nU�*jf�*nU jf�
nU(jf�*nU(jf�*nU(jf�*nU�*jf nU�
jf(nU�*jf(nU�*jf(nU�*jf(nU�*jf�*nU          �*  �  "�  "�  "��"�
�"�
"�
"��"�Z"��"�Z"��"�Z"��"�Z"��"�Z"��"�Z"��"�Z"��"�Z"��"�Z"��"�Z"��"��0l1l1���������������<3�03332>?û��?����۟��V[k�EVViQ�XA��F@fEQQUQPEUUDUUUUUUUU      ?  ��  ��  ��  ��  ��  �; ��; �p� ���� �U����� ��� ����� W5  �? �W5 �W� 0_U0�U��W:�W�g��W��� ��5 ��� ������     �   �  �  �  �  �  ��  �C W��U� �~� �� ��� \�  ��  \� W��U�pU�Տ:��0p�00������� [� \� W�ð�������     �  ,  ,  ,  �< ��|UU\Zi|UU���j�5�e�5���5�]�=���; Ǵ����U� pWup�_p5Wp\�� p\|\p\����\\�:�:�?�?     �  �:  08  00  <� ��>�ʏ>�*�:��j=pWU7\�_�\5\�\5���?|��5|���� �?� 7|�����|��_�5p /��5p�5p=�5p�7p?�7pp5p5�������      ?  ��  ��  ��  ��  ��  �; ��; �p� ���� �U����� ��� ����� W5 ��� �U��U�U-�U����p�� p5 |6 _�� ��� �   ;              �   �  �  �  �  �  ��  �C W��U� �~� �� ��� \�  ���sU�pU0xU��U�× �o �\ 0�= �~� ���   �   �   �   �      ?  ��  ��  ��  ��  ��  �; ��; ������U�0�������0 ��� �  �?  W5  �?  W5  W�  _U �� \�  W� �Y� p�� l�� �Ճ�� ?�  �:  �?     �   �  �  �  �  �  ��  ����U��?����  �  ��  \�  ��  \�  W� �U� �V>  �5  _�  �e _ _9��W��0�� �?  �                    � ��? 0�� �W� �������0���_U0������ s]� �]� 0�� ��?  �          � �� �W� �������0���_U0������ s]� �]� ��  �             �  � �������� �  �� ����UUp����Vp�V������  �?          �  0  �  �  0  �� ����UUp����Vp�V������  �?      �?  0< �?7 ���^��W���_��_ \��_����^� �� �?7 0< �?        < �?7 ���^��W���_��_ \��_����^� �� �?7   <     ��  �� �� �� �� ��  �9  �?  �  �?  ��  30��� ?         ��  �� �� �� �� ��  �9  �?  �  �  �  �  �  �  �?       � ��?|�7;W�7�U���W���^�� {���^��W���V�7;k�7��; ��?  �      � ��? |�7 W�7�U���W��ް��߰׫^���W���V�7 k�7 ��; ��?  �    0   �� ?�� ��0���Ϫ��:�ί:\��5���:�������V:0 ��� �?   0   �� ��� ����pj�����:�.�:�5x:���:�������: ��� �
3           �3  �� ��:��� �� ��� �:��  ��  �   0          �3 ?�3���0���"�*/  � *  �  �;  �?  8,  ��*�̿�� �� ����<�<�0�0�?��>/�/�/�?��>�  �<?<<<<�<�  ��������,8,8,8,8,8,8,8,8  ����    ����      ����  ��        00?0?0    ���?�:�����3  �3��<�<;��;��;��;��<�<3�?�3  ������:����?����0�������  �3�?�?<<�?<<�?�?�?���3����  ��������0������� �( �� �p�p�����+�2��������*����:��:� �  ��������?�������3  �?��;<<�;< �;��; ?�;?�;�?�?  �3  �����������?����  ����� �33�3�0�����k����5���������:�������                                                                �             � ?            0��?           �*��?         �����:        �����         ?�����         ?�����       ������       0�����        0�����        �*�
�          �*����������
 �*�ʪ�"       00������������ �à�, ���� ���� ��*���*���ꫪ�ʢ����?�������2�" ��0��0� ��" ������������" 򪪪��������������:����������������*���������  ����������>   ������������  �ê:�ꬪ��Ϊ ������￿���? <Ϫ��:�� �>� <�����;<��� <�������?;���� ��������?;��� �?����;<���   00��  >  <3�3���?3���  ������������           <  � ������:������  �  �  �: ��� ��� ��� ��� ���  �:  �   ���Sݫ�����    ��W׬��    �> ��@5>�@5�  �@5>�@5�  �@5>�@5�  �@5>�@5�  �@5>�@5�  �@5>�@5� ��>         ���?��������?       � 00998900� �� ��  � 1���  ���-J�J�(J�8J�BJ�MJ�SJJ�pLj� ɐ ��� JJJJ�5J�;Lj�` � ��� JJJ�!J�'Lj� ��JJ�J�Lj� ��� J�J�Lj� )�J�Lj� ?�J�Lj�J���� �е�f 	��f  ��Lj� ��Lj�HJJ��� 	�� L�J��� 	�� h`HJ��� 	�� L �J��� 	�� h`�e J�(�e )��e �z �� � � ��8�� ���� L0�� �� `��| �e )��e `H�� �� �e J�@�e )�	�e �� � �/ ���� ��� JJJJ��� ��  ��8�� ���� L��� �� h`H ���� )�	��  ��h`H ���� )�	�� ��|  ��h`H�� )�	��  ���́ � ��΁ �e 	@�e h`H�� )�	��  ���g JJJJ�� ����L��� �(�L��� ��L'� ��� �e 	@�e h`H�� �� �Z �[ �\ �] �^ �_ �� J�J�J� J�*L�� Ւ�Z � �*L�� 7��Z � �L�� ���Z � �L�� ��Z � �L��h`�� J�J�	J�L�� P��Z � � P��Z � � �ꭝ �o )
�o ����o �� )�o �� L��� �n 8�� ��T��P�Z �� i
�[ �� JJJ��Z �\ 8�[ ��[ �[ i
�] �� JJJJ��Z �\ �^ �� �[ i�] i�_ `��n �� i�+�S�Z �� i
�[ �� JJJ��Z �\ 8�[ ��[ �[ i
�] L���� JJJJ��Z �\ �^ �� �[ i�] i�_ `��n 8�� ��Y�[ �� i�Z �� JJJ��[ �] �� �Z i�\ L ��� JJJJ�'8�� ��Z �� i�\ �� i�^ �[ �] �_ L �`��n �� i �x�V�[ �� i�Z �� JJJ��[ �] �� �Z i�\ Lf��� JJJJ�$8�� ��Z �� i�\ �� i�^ �[ �] �_ `��o �n � ���!��#��%��'��)��.��'Lϔ ДLϔ וLϔ �Lϔ T�Lϔ ��Lϔ ��LϔLĔ���  ��Lϔ���  ��Lϔ`�� �� �� �� �� )�� �� ��  ���� �� �� �� �� )�� �� �� �� `�� �� �� �� �� JJJJ)�� �� ��  ��� �� �� �� �� 



�� �� )�� �� �� �� `�� �� �� �� �� JJ)�� �� ��  R��� �� �� �� �� 

�� �� )�� �� �� �� `8�Z ��.�Z � ����LՕ�� �(�� ���� N��o LՕ�o LՕ``8�Z �!����Z �[ i�q��[ L���Z L�� �o `�[ �`�8�Z ��9�Z L.�8�Z ��Z �[ i�[ L.�� �������� N��o LQ�� �o `�[ �P��Z i�,�9�Z L~��Z i�Z �[ i�[ L~�� �������� N��o L��� �o `�Z �$���(���� ����L�8�Z ��Z �[ i�[ L�8�Z ��Z 8�[ ��[ L햜o ` ?�� ����Lc��� J��l �
�W �Lc��e 


�L�� � �K�� 



�B�� �
�,�� i�,�t�� �� JJ�8�� ��� Ll��� i�� Ll� <�Ll�L�� %�L���� � �N�� 


�F�� �
�8�� i�,�#�� �� JJJ�8�� ��� L���� i�� L���� )��� L�� P�L��`�� � �B�� 

�;�� �
�.�� i�,�ύ� �� JJJJ�8�� ��� L
��� i�� L
� d�L
� %��� �� ����� �� I�� L���� 



�E�� � �>�Z �� �[  F�� 
��LN�� �� �խ� �X �� �Y  F� � �ޭn � � ���� 


�E�� � �>�Z �� �[  F�� 
��L��� �� �խ� �X �� �Y  F� � �ޭn � � ���� 

�E�� � �>�Z �� �[  F�� 
��L瘩 �� �խ� �X �� �Y  F� � �ޭn � � ��`�� �� 	�� ��� �� �� ��� �F�� �b�� �� �� �� �� `�� 



�L�� �� ���� �n  �� F�� �Z �� �[  ��L���� �� I�� J� ��� )�� �� 	�� �� �� 


�K�� �� ���� J�n  �� F�� �Z �� �[  ��L癜� �� I�� JJ��� )ߍ� �� 	�� �� �� 

�M�� �� �� �� JJ�n  �� F�� �Z �� �[  ��L;��� �� I�� JJJ��� )��� �� 	 �� �� `�� 	�� �� �� )��� `�� 	 �� �� �� )��� `�� 	@�� �� �� )��� ` ?�� ����L���� J��m ������L���l �F�O ��L���� � ��� ���� L���� �p�i�� �� � �$�� ��L���� JJJJ��� 	��  <�L��L���� ��B��� �p�!i�� �� � �/�� ��LF���� �� LF��� 



��� 	��  P�LF�L���� � �I��� �p�!i�� �� � �3�� ��L����� �� L���� 


��� )��� �� 	 ��  d�L�� %�`�� �� �� 	�� �� 	��� ��� �� �� �� �� �� �� �� `�� J�J��� J�	J� 4�L3��� JJJ�J��� JJJ�	J� ��L3��� 


�J��� 


�	J� ޜL3��� 
�
��� 
�	
� 3�L3�`�{  ���o ��  ��X �� �Y �� �� )��� �f )��f ` ���o ��  ��X �� �Y �� �� )��� �f 	�f `�{  ���o ��  ��X �� �Y �� �� )��� �f )��f ` ���o ��  ��X �� �Y �� �� )��� �f 	�f `�{  ���o ��  ��X �� �Y �� �� )�� �f )��f ` ���o ��  ��X �� �Y �� �� )ߍ� �f 	�f `�{  ���o ��  ��X �� �Y �� �� )��� �f )��f ` ���o ��  ��X �� �Y �� �� )�� �f 	�f `�x 
m  m� m� m� m� **� ��@�#�`�'ɀ�+ɠ�/���3���7���;L��� �o L ���o L ���o L ���o L ���o L ���o L ���o L ���o L �`�o � ���(��1��:��C��L��U��^L'��,�X �,�Y L���,�X ��Y L���,�X � �Y L��� �X � �Y L���,�X ��Y L���,�X �2�Y L���,�X ��Y L���,�X �<�Y L��`�m� �� �� i �� �� i �� �`���s ��Z ���[ ��  ў��  ў��  ў�  ў`�)�JJJJ��  螊)��  �`xH�Z�� �a��$��b��%��c��&��d��'�����X ����Y ��n �[ ����V ����W 8�>�W �Z �X-s �V�X ȲX-s �V�X ��n ���Z �Z z�hX`
��j��v �j��w � �v�$�*�a��b��c��d�8�7��  螭f 


� [� ��Ȁ�`H�y �  ����y �0�h`H�  ����h`��e �e `H�Z�X �@�Y � � � �X����Y ���z�h`                          �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  �?��ʫʫʫ���?�*V�V�V�V�V���*      �?�?        ����  �    �  +>  �  ?����\= ��� �W���W����� �\= ����  ?�  �  +�  �?  �  +>  �  ?� ��� \=� ��� W�� W�� ��� \=� ���  ?�  �  +�  �?��?Wp�W���  �7��<�?< ,8  �2  �2  << <�?<7���  �W��Wp���?        �?�p�Wp�Wp�p-x������p=|p�p�Wp�W�?�                              �  ����� ������� ���  ��                      ?  �  �   �� �� � ������������� �  |  �   ?     �  �  �5   � ��W\U]��]5WUu��u�\UU��U��UU� �U=  �                 �?  \� ��Up�_��]5pw�p�u����p�]��]� WW= ��              �? 0��?����?������������:��������� ����� ��� ��?              �?� 0���?�����������������:�ê:���?  �  �  �   ��  �U �U= pU� p�pTpU=pU5pUU��UU��U����<�� �� �0    ��  �U �_5 ���  �W��?�=���7������������ ��� �_= W� ��           ,  ��  �  <      �����  �    <  0  ��   /              #  �   0�  <�    �
��� �
   <�  0�  �    #     �? �������������� ;�  ��  ��  ;� �������������� �?  �? ���������:��:�����  ���3���3��  �����:���:������ �?      � �3���� � �S�?�T�T3�T3�T�S�������3� �          � �3���� � ���?��?��?3��?3��?���������3� �     00�� �  � �0���0���0�;�§�[�p��\��5��?�7,9�,90 ,9  � ����p�|=��w��s5\��_�{p���s���s�����W=�]u3��03���� � ����:,�8,�:80���>�3�������>�30��,�:8,�8��:�� �  ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                   ��        �      ���      ?j�2      3ڟ2    ����:    � 3�2    ����:      3ڟ2      3j�2     0̨�    ����    �������  ������� 0������ W��gf�U ������  0W��gf�U ������٪  ��������������� �}�����  �������  �]WUUUU=����UUU�\�]U������7����������U���������U}�UUi]���U}�   \���U}�   ]���U}�UUU]���U�uUUU�����������]U������7���UUU�\�]WUUUU=��������  �}�����   ���������   ������ ������٪ 0W��gf�U ������  W��gf�U 0������ �������  �������   ����     0̨�      3j�2      3ڟ2    ����:    � 3�2    ����:      3ڟ2      ?j�2      ���       �       ��    �       "  *  �  �  ���*��
���*�!B)` h	h�!X��(X*Z��
h�� HY*���*(T`�*j�
 ��*���(��* 
�*���
 ��  ��
 �� �  �  �    "  " � �� �(�b
�*�**j**bJ)bR(bR�X��j��j���Z)�V&�Z$�Y)��)��*�(
���� (  �  �  
   * ��" `�� ���(��
(�Z*�*�*h
d�& �
�H�*H�i* j�
�d����@�* � �������} ���} ��p Lc��} ���} ��p Lc�� �p �� J� ���� JJ� ��� JJJ� ���� JJJJ� ���� 



� q��� 


� 䯭� 

� X��� 
� Ͱ` �� C��n � �L�� �n �p � �*�� �� �� ��  g��o � �,�Z �� �[ �� �� I�� �� �n ��  �� F� ��L� �� �ڜo �n `�� �Z �� �[  C��n � �M�� �n �p � �*�� �� �� ��  g��o � �-�Z �� �[ �� �� I�� �� J�n ��  �� F� ��L�� �� �ڜo �n `�� �Z �� �[  C��n � �N�� �n �p � �*�� �� �� ��  g��o � �.�Z �� �[ �� �� I�� �� JJ�n ��  �� F� ��L�� �� ,ۜo �n `�� �Z �� �[  C��n � �O�� �n �p � �*�� �� �� ��  g��o � �/�Z �� �[ �� �� I�� �� JJJ�n ��  �� F� ��Lp� �� xۜo �n `�� �Z �� �[  C��n � �P�� �n �p � �*�� �� �� ��  g��o � �0�Z �� �[ �� �� I�� �� JJJJ�n ��  �� F� ��L� �� �ۜo �n `�� �Z �� �[  C��n � �Q�� �n �p � �*�� �� �� ��  g��o � �1�Z �� �[ �� �� I �� �� JJJJJ�n ��  �� F� ��LW� �� ܜo �n `�� �Z �� �[  C��n � �R�� �n �p � �*�� �� �� ��  g��o � �2�Z �� �[ �� �� I@�� �� JJJJJJ�n ��  �� F� ��L̰ �� Yܜo �n `�� �Z �� �[  C��n � �S�� �n �p � �*�� �� �� ��  g��o � �3�Z �� �[ �� �� I��� �� JJJJJJJ�n ��  �� F� ��LB� �� �ܜn �o `��n �e JJJ�J�Z i�o �� �o �9�� i�o �Z �o �(�[ i�o �� �o ��� i �o �[ �o ��n  ��`�e JJJ�!�� ��8�� ��� �e 	�e �� Lı 
�`�g 	�g �{  �ͩ�� ��� �"�� �� ���  �� �̭{ ��!�{ �� J�J�	L� ��L� �L� u�L� � d� ���g J�- (� 9� Q��k  �ѭ� ͱ ��� ͱ � 
� [� ��L�`�� �b �� �c L̭� �Z �� �[  ��� 6� �խ� �Z �� �[  ��� 6� ��`�
�a �<�` `�� � �I�� � �B�� � �;�� � �4 ���� � ��� i�@�!�� �� �� � ��� i�@�
�� �� L�`�� )�	��  ���� �"�� �D�� �� L� � �\�� � �U�� � �N�� � �G ��� � �8�� ���� �� � �+8�� ���� Lt��� )�	�� ��� �"�� �� ��  V�`�� � �P�� � �I�� � �B�� � �;�� �
� V��� � ��� i��!�� �� �� � ��� i��
�� �� L̳`�� )�	��  ����� ��� �"�� �� L̳�� J�J�	L� �L� ɴL� Q�L�`�� � �Y�� � �(8�� ���	�� �� LD��� ��  $� +� ˷ � $��� � �#8�� ���� ��  2� 9� �� �Ln��� �� �� � �S�� � �"i�,��� �  N� U� U� l�L���� �� �� � �#8�� ���� ��  @� G� '� >�Lȴ�� �� `�� � �>�� � ��� i���� L𴍠  $� ˷�� � �8�� ����  2� ��L��� �� � �;�� � �8�����  +� �L2��� �� � �8�� ����  9� �LP��� `�� � �b�� � �/8�� ��n �� i�n �	�� �� L���� �  $� +� ˷ ⷭ� � �%�� i�p�	�� �� L���� ��  2� 9� �� ��� � �b�� � �%�� i�p�	�� �� L�� ��  @� G� '� >��� � �/�� i�n �� ��n �	�� �� L#��� ��  N� U� U� l�` �� \�` �� \�` 6� s�` �� s�` �� s�` � s�` i� \�` �� \�` h�� �� ��`��a ��` ` �� �� ��`��a ��` `�� � �48�� ��� �� �� i	�� i�� �� i�� i�� 8�� ��� �� �� � �4�� i	�� i�� �� i�� i�� 8�� ��� �� �� i
�� �� `�� � �#��� �� i	�� �� ����� 8�� ��� �� � �#��� �� i'�� �� ���&�� 8�� ��� `�� � �2�� i�� i�� �� i<�� �� �� i
�� �� �� �� i�� �� � �4�� i�� i�� �� i<�� �� 8�� ��� �� �� i�� i�� ` �� h� � �ޭn � � ��` �� h� � �ޭn � � ��` � � � �ޭn � � ��` k� � � �ޭn � � ��` �� � � �ޭn � � ��` � � � �ޭn � � ��` L� h� � �ޭn � � ��` �� h� � �ޭn � � ��`�� � ��� �X �� �Y  �� � �ޭn � � ���� �X �� �Y  �� � �ޭn � � ��` �� [� z�f 	 �f ��Z �(�[ � ]���Z �2�[ � ]���Z �<�[ � ]���Z �F�[ � ]��n  ���n �n �
�� �� [ө�Z �
�[ � ]���Z ��[ � ]���Z �(�[ � ]���Z �2�[ � ]���Z �<�[ � ]���Z �F�[ � ]���Z �P�[ � ]���Z �Z�[ � ]���Z �d�[ � ]���Z �n�[ � ]���Z �x�[ � ]���Z ���[ � ]���Z ���[ � ]�L� z� �� [�d � �� ��  
�
���I�L�� �� ��` �ө(�[ ��Z �  ]��<�[ ��Z � ]��<�[ ��Z ��  ў��  ў��  ў�  ў�F�[ ��Z � ]��F�[ ��Z ��  ў��  ў��  ў�  ў�Z�[ ��Z � ]��n�[ ��Z � ]�����h 	�h �Z�[ ��Z  �L庭h )��h �n�[ ��Z  �L� [�`�	 ���a ��`  ��`�� �� �� �� ��� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �l �� �� �� `�n )� ���&��;��KL̻8�Z ��V��R�Z �\ �^  ͻL̻�Z i�+�9�Z �\ �^  ͻL̻8�[ ��"�[ �] �_ L̻�[ i�x��[ �] �_ L̻�Z �[ `�� � �M����"L!��[ i�x�3�[ �] i�] �_ i�_ Lͻ�[ ���[ �] ��] �_ ��_ L!��Z �[ `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ���ة��  ��� ��q � � �r � �ύ& ��"  P� t ����X ��Y �� � �X����Y ��� ƟX�P�U �# L �H�Z�x �y �z �{ �} �~ �� (z�h@H�Z�' )�	 ��U �# �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                                                                         � z� ,� {� �� 
� ,� ũ �J  Y�g J�3J�< ǭh J�� v� 9� ^� (��f 
� z� ,� �L� 
� Q�L\� C� [� ��L � �h JJ�� z� ,� �L©�Z ���[ ��\ ���] �i �i I�i � �
�[ �[ �D�c��a �[ ɐ���8�[ �` L�©�` � �� yխ[ �r�V�Z �^ �[ �_ �] �] �C�!�[ �\ �Z ��a �] ɏ�8���] �` L� ��L0é�` � �� yխ^ �Z �_ �[  ��L���Z �Z �	�]��a ��` � �� yխZ �^ �[ �_ �\ �\ �Z �] �[ ��a ��` � �� y��\ i�n  �í^ �Z �_ �[  ��L0é��N  ��i  ���i �i �x��i `�Z H�[ H�D�[ �n �Z ��a ��` � �� y�h�[ h�Z ` �� [ө(�a ���` ��Z � �[ � �� �ө�J  Y�  
�� z�`�� �� �� �� �� ��� `�� �l �j �i ��k �m �c ��b �e ��f �g �h ��� �� ��� ���s �P�� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �{ �} ���� ���� �� �� �� �� �� �� �� �� �� �� `�� `�o  �� [ӭo ��& G� [ӭ{ ����{  �� [ӭ{ ����{ �o L�`�<�[ ��Z � ]��<�[ ��Z �  ў�Z�[ ��Z � ]�` }� 5�`�� � �{�l ��t� ����-��G����!L�ŭm � �d��X��T��H��T��HL�ŭm � �>��J��.��J��6��*L�ŭm � �(��,����$����L��`��� L(Ʃ�� L(Ʃ�� L(Ʃ�� L(Ʃ�� L(Ʃ,�� ��� L�ŭ� � �= �ƭn � �	 ���� LyƩ��T ��H  )�� �� ��������?��JLy�`� Lyƭ� 	�� Lyƭ� JJJ�J�Lyƭ� 	�� Lyƭ� )�	�� Lyƭ� ������ Lyƭ� ������  ��Lyƭ� �X �� �Y  F� � ��`��  �� F�� �Z �� �[  ��`�x ��8�x �e 	 �e �l �i �i ̀ �'�l �� �� �m �m �� O�LNǜi LHǭe )ߍe  �� ��`�g 	�g � ������������L�� u�L�� ��L�� űL��`�i ��  �� �� �� �� � 1� 
ԭg J�" (� 9� Q��k  �ѭ� ͱ �
 [� ��L��`��b ��c L̩�� �� ��� �� ��� �� ��� �� `�,�� �� �� �� �8�� �� �� �� `��a �p�` ��Z ��[ � ��`�i ������LU� V�LU� �LU� ;�LU�` f�8�� ���E�� �� 8�� � �O���7�� �� 8�� � �;���)�� �� 8�� � �'����� �� L�� ��L�Ȝ� L�Ȝ� L�Ȝ� L��`�i �i ����L�� �ǩ�� �� �� �� �T�� �� �� �� Lɩ�� �N�� L�` fɭ� ����� L:��i ��� �
�� ��� ��� �� �� �� �� L:�` fɭ� i�x��� �� �� �� �� Leɜi  �� ��Le�`�i ����k��dL�ɭ� � ��� � �%�� � �3L�� � N� � �� �� � +� P�L�� N� � �� � +� P�L�� � �� +� P�L�� �� P�L��`L� �� �� � �� �� � � �ޭn � �� ��L�� � N� � ��L�ɩ�a �(�` ` ��i ���L.ʩ �� �� �� �� �� � �ޭn � � ��` ��i ���L_ʩ �� �� �� �� �� � �ޭn � � ��` 6�i ���L�ʩ �� �� �� � �� � �ޭn � � ��` ��i ���L�ʩ �� �� �� k� �� � �ޭn � � ��` �� �� �� �� �� �� � �ޭn � � ��` � �� �� �� � �� � �ޭn � � ��` i� �� �� �� L� �� � �ޭn � � ��` �� �� �� �� �� �� � �ޭn � � ��` �� �� �Ӝx �{ �} �� �� �� �� �� �� �� �� �� �� �� �� �� ��Z �b �X�[ �c  s� [� �� 
� Qέg J�" (� 9� Q��k  �ѭ� ͱ �+ [� ��L�� C� s� Q��k  �� [� �ӭg JJ��L�`�� �� )��� �� 	�� �b i�� �c i�� �� �� )��� �� 	�� �b i�� �c i�� �� �� )��� �� 	�� �b i�� �c i�� ��  ��L̭� )�	�� �n �o �x  �ӭo ��H�� ��
�� �_�	L��΁ L���� i�� L�̭x �(�	�x �o �n �n J� ��  � [� ��L��`�� ��L:� �� k� ^ͭ� J�� �� �� ^ͭ� JJ�� �� ��� JJJ��� �� 	�� L�� z� �� [�� � ���P�� �h 	�h ` ɸ  � Q��k  �� [� ��`�~ ���~ �g )��g �b �Z �c �[ �  6� F� ���b i
�Z �c i�[ �g 

�� ��L�ͩ
 ���a �
�`  ��`�� J�Lέ ��������L�ͩ��� L5Ωȍ� L5ΩP�� L5έ ��������L-Ωd�� L5Ωd�� L5Ω(�� L5�`
��.��t �.��u `��a �(�` `�� J�B�{ ��_�{ �� ��L{��b �b ��b �EL���b �b ��b �5L�έ� )��� �x L�έx �(��� 	�� �b ����� L�Μ� L�� sͭe JJJ�,�b �X �c �Y ��a �(�`  � �ޭn � �	 ���g J�a �� �� .� g� �� �� � Lѭg J�C�� � �<�� � �5�� � �.�� � �'�� � � �� � ��� � ��� � � Vϭg 	@�g `�b i
�� i�� i�� i�� i�� i�� i�� �c �� �� �� �� �� �� �� �b �� �c i�� ` �� � �ޭn � � ���n `�� � �18��)�� �Z �� 8���� �[ �  }� �� �ϭn � �L�Ϝ� `�� � �18��)�� �Z �� 8���� �[ �  }� �� �ϭn � �L-М� `�� � �18��)�� �Z �� 8���� �[ �  }� � �ϭn � �LfМ� `�� � �,�� 8��!�� �[ �� �Z �  }� k� �ϭn � �L�М� `�� � �3i�,�)�� �Z �� 8���� �[ �  }� �� �ϭn � �L�М� `�� � �3i�,�)�� �Z �� 8���� �[ �  }� � �ϭn � �Lќ� `�� � �3i�,�)�� �Z 8�� ���� �[ �  }� L� �ϭn � �LKќ� `�� � �)8��!�� �Z �� �[ � }� �� �ϭn � �L|ќ� ` 7� �� ��`�e 


�8�k ���k L�ѩ�k  F�k �Z ���[ � ����������L�ѩ  ��L�ѩ ��L�ѩ ��L�� ���Z i�Z �,��`��a ��` ` :�� �V�qV�n �i �n � N�L��i i(�n � �V�n �L9� `� N�L�`� :
��7��V �7��W `�V i�V �W i �W `� �V�i �8�i �Z � �\ L�ҍn 8�i �n �\ � �Z ��V�[ �] ��V�a ��V�` �e 


� ��V �� ��`
��{��t �{��u `�[ ����v ����w 8�>�w �Z imv �v �w i �w 8�a �\ �o �Z �n � � �\ mt �t �u i �u �t-s �v�Z �Z �,���o ��n �Z �v i0�v �w i �w �t mo �t �u i �u ��` Ц`Z��u �t �@�Y �X � ��t�X����Y �u ���z`��u �t � �� �t����u ���`��u �t �p �o � �� �t�o ɀ�#�p �p ���0�	�p �o L������u ���L������u ���`��u �t � ����t����u ���` �� S� ��` I� �� Sխe JJJ�*� �� ��#�������������e )��e  ��`�e J�a�� �_�Z�z �| �S ���� )��Luԭ� 	�� �� i�_�	�� �z L�ԭ� �_�!�_�� �� �n )��
�� 	)��� �z L��`�e 

���� J�J�	L��� L��΁ L�ԭ� J�J�!J�4J�6LRծ� �_�JJ�-L��JJJ�*�LRծ� �_�J�2L�JJ�0� LRթLRթLRթLRխz �� ���� )��� �LRթLRխz �� ���� )��� �LR�`
�����t 轢��u ��a � �` �� �Z �� �[ `�[ ����v ����w �Z mv �v �w i �w � � �t-s �v��a ���v i0�v �w i �w �t ma �t �u i �u ��` ��`�[ ����v ����w 8�>�w �Z mv �v �w i �w � � �t-s v�v��a ���v i0�v �w i �w �t ma �t �u i �u ��` ��`��\ ��]  M� 5� �`�� � �B�� �Z �� �[  ٭n � ��� �n �� �o  )߭Z �� �[ �� L�֜� ��n  ��L�֭� � �G�� �Z �� �[  ٭n � �"�� JJ�n �� JJ�o  )߭Z �� �[ �� L�֜� ��n  ��L��`�� � ���� �Z �� �[ �٭n � �&�� JJJJ�n �� JJJJ�o  )߭Z �� �[ �� L�֜� ��n  ��L�֭� � �?�� �Z �� �[  ٭n � ��� �n �� �o  )߭Z �� �[ �� L{ל� ��n  ���� � �G�� �Z �� �[  ٭n � �"�� JJ�n �� JJ�o  )߭Z �� �[ �� L�ל� ��n  ��L��`�� � ���� �Z �� �[ �٭n � �&�� JJJJ�n �� JJJJ�o  )߭Z �� �[ �� L�ל� ��n  ��L�׭� � �B�� �Z �� �[  ٭n � ��� �n �� �o  )߭Z �� �[ �� Lc؜� ��n  ��Lcح� � �G�� �Z �� �[  ٭n � �"�� JJ�n �� JJ�o  )߭Z �� �[ �� L�؜� ��n  ��L��`�� � ���� �Z �� �[ �٭n � �&�� JJJJ�n �� JJJJ�o  )߭Z �� �[ �� L�؜� ��n  ��L�حg JJJJ�k jڭn � �` �ڭn � �V �ڭn � �L Hۭn � �B �ۭn � �8 �ۭn � �. +ܭn � �$ uܭn � � �ܭn � � �ܭn � � ��Lu�`� ����L�� �� �ޭn � ��� L������L�� � �ޭn � ��� L������Lu� 6� �ޭn � ��� L�� P� �ޭn � Е�� L�٩��T ��H  )�Lu٩�\ ��] �b �X �c �Y ��a �(�` `��\ ��] ��X ��Y ��a �p�` `��\ ��] �� �X �� �Y  ��`��\ ��] �� �X �� �Y  ��`�� J� �� F� �ޭn � �	 �� ��n `�� �X �� �Y `�� 	�� �� 	�� �� )��� �� `�� JJ� �� F� �ޭn � �	 �� ��n `�� �X �� �Y `�� 	�� �� 	�� �� )��� �� `�� JJJ� � F� �ޭn � �	 ,� ��n `�� �X �� �Y `�� 	�� �� 	�� �� )��� �� `�� JJJJ� k� F� �ޭn � �	 x� ��n `�� �X �� �Y `�� 	�� �� 	�� �� )��� �� `�� 



� �� F� �ޭn � �	 �� ��n `�� �X �� �Y `�� 	�� �� 	�� �� )�� �� `�� 


� � F� �ޭn � �	 � ��n `�� �X �� �Y `�� 	 �� �� 	 �� �� )ߍ� �� `�� 

� L� F� �ޭn � �	 Y� ��n `�� �X �� �Y `�� 	@�� �� 	@�� �� )��� �� `�� 
� �� F� �ޭn � �	 �� ��n `�� �X �� �Y `�� 	��� �� 	��� �� )�� �� `�g 



�*�� �X �� �Y  F� �ޭn � ����N  �� J��� `�� J�V�� 



��� � �
 Oݭn � �4�� 


��� � �
 rݭn � ��� 

��� � � �ݭn � �LNݩ��N  ��`�� �X �� �Y  F� �ޭn � �	�� J��� `�� �X �� �Y  F� �ޭn � �	�� J��� `�� �X �� �Y  F� �ޭn � �	�� J��� `�� J�<�� JJ��� � �
 2ޭn � ��� JJJ��� � � Uޭn � �L�ݩ��N  ��`�� JJJJ��� � �
 xޭn � �ݭ� 



�ܭ� � �� �ޭn � ��L�ݭ� �X �� �Y  F� �ޭn � �	�� J��� `�� �X �� �Y  F� �ޭn � �	�� J��� `�� �X �� �Y  F� �ޭn � �	�� J��� `�� �X �� �Y  F� �ޭn � �	�� J��� `�Z m\ �o �X �o �:�X ma �o �Z �o �(�[ m] �o �Y �o ��Y m` �o �[ �o ��n `��n L	߭� �Z �� �[ ��\ � �] ` a߭Z � � 9�`
�����t 轲��u `�� J��  7�L]ߩ 7�L]� ��`�o )�o �n )� ���'��d��nL�8�Z ��s��o�Z �o � �n �L�g JJJJ�� ��!��L���Z i�+�>�Z �o � �= �L��Z i��$�Z L�8�[ ���[ L��[ i�x��[ L��Z �[ L�`�o ����L8��[ i�x��[ L8�8�[ ���[ L8��Z �[ `�g JJJJ�� ����LW�Z �� G� ��` � �� � x� � +��f )��4�{ ��7�{ �f J�J�J�J�L�� `�L�� ��L�� 
�L�� _�L��{ �2� ˛`�� JJJJ� ��L��� �
��g )�g �� 	�� �� �� L��`� �� ��g 



�T�e 


�!8�� ��9��  k�n � ���  ���g J�íg I �g �� �Z �� �[  F�  � ��L��g )�g LO�l �FБ�<�� �,�� �g 	�g L��� �X �� �Y  F� � ��`�� �� ���� �n  �� F�� �Z �� �[  ��L��� �� I�� J�L�� ��� )��� `�� J�o�� JJ��� i�,�R�� L��8�� ��D�� L��� JJJ��� m� ɀ�+�� L�8�� �� ��� L� ��n � � ��L/� ��L:�� )��� L:�`�g 



���� 	�� �� ́ ��� )��� 8�� �� �n L~�� 	�� 8�� � �n L~�� ͂ ��� )��� 8�� �� �o L��� 	�� 8�� � �o L��Nn No �n � ��o �� �� �� �� �� L:�� �X �� �Y  �� � ��`�� �Z �� �[ �  7� �� ��`�g 


�� ��L� ��`�� J� k�� JJ� ��� JJJ� ��� JJJJ� C�� 



� ��� 


� ��� 

� )�� 
� v�`� �� ���� �n  �� F� �� y�L�㜢 �� I�� J�L��� )��� `�� �Z �� �[ `� �� ���� J�n  �� F� �� y�L�㜥 �� I�� JJ�L��� )��� `�� �Z �� �[ `� �� ���� JJ�n  �� F� 6� y�L5䜨 �� I�� JJJ�L5�� )��� `�� �Z �� �[ `� �� ���� JJJ�n  �� F� �� y�L�䜫 �� I�� JJJJ�L��� )��� `�� �Z �� �[ `� �� ���� JJJJ�n  �� F� �� y�L�䜮 �� I�� 



�L��� )�� `�� �Z �� �[ `� �� ���� JJJJJ�n  �� F� � y�L圱 �� I �� 


�L�� )ߍ� `�� �Z �� �[ `� �� ���� JJJJJJ�n  �� F� i� y�Lh圴 �� I@�� 

�Lh�� )��� `�� �Z �� �[ `� �� ���� JJJJJJJ�n  �� F� �� y�L�圷 �� I��� 
�L��� )�� `�� �Z �� �[ `���T ��H  )�`�g JJJJ�/�(�[ ��Z � ]� [� �� �� z�  
�� �� �� �J  Y�`�g 	�g �� �� �� �� i�� �� �� i�� �� �� i�� �� �} `���T ��H  )��n �} ���} �n  �� �� � Y筠 � �"�� � ��� � ��� � ��g 	)��g  ��`�� �Z � �4�� �[  F� �� �խn ��8�� ���� 8�� ���� L�朠 `�� �Z � �6�� �[  F� �� �խn ���� i�,��� 8�� ���� L眣 `�� �Z � �6�� �[  F� �� �խn ��8�� ���� �� iɐ��� LX眦 `�� �Z � �8�� �[  F� �� �խn �� �� i�,��� �� iɐ��� L�眩 `Hڪ���




�p ��)p �& �h` ��
�����t 轓��u  �� [өύ& `�n J�� ��L�� ��`�� �� ���� �� ��
�� �� �� �`�� �� �� �� �� �� ` (� R� ~�`�� �� �� �� �� )�� �� ��  ��� �� �� �� `�� �� �� �� �� JJ)�� �� ��  ��� �� �� �� `�� �� �� �� �� JJJJ)�� �� ��  ��� �� �� �� `�� � �l�� J��� i�,�Y�� L��8�� ��K�� L��� JJ��� m� m� ɀ�0�� L�8�� �� �!�� ��� L�  �n � � ��L� 6�L�� `�� �X �� �Y  �� � ��`�� �Z �� �[ �  7� �� ��`�� � �*�� ́ ��� 8�� � �n L���� 8�� � �n L��`�� ͂ ��� )�� 8�� � �o L��� 	�� 8�� � �o L��Nn No �n � ��o �� �� �� �� �� L�o � ��7��3L��n J��o 
�����t 轾��u LE�o 
�����t ����u LE�n J��o 
�����t ����u LE�o 
�����t ����u LE�`��a ��` ` X� ��`�� H�� �	���� ��a ��` ���[ ��Z �  �� ���Z i�Z �� ����� ��h�� `
�����t ����u `�Z������ ���� ��z�`�Z����� ���� ��z�`�� � �l�� )�n �� �� )�� �� �Z �� �[ ��  9ଡ଼ JJJ�J�LH�\ �� �Z �] �� �[  9ଡ଼ JJJJ��^ �� �Z �_ �� �[  9�LH�L�뭋 � �z�� )� �n 

� �� �� )�� �� 

� �� �Z �� �[ ��  9ଡ଼ JJJ�J�L��\ �� �Z �] �� �[  9ଡ଼ JJJJ��^ �� �Z �_ �� �[  9�L��`�� � ���� )ύ� �n 



� �� �� )ύ� �� 



� �� �Z �� �[ ��  9ଡ଼ JJJ�J�L��\ �� �Z �] �� �[  9ଡ଼ JJJJ���^ �� �Z �_ �� �[  9�L�� � � � � � � � � � � �( �) �* `� � � �  !� %� � � � � � � � �* �G �P � ���H �T `� ���%�+ � !�$ � �% �  W��+ �+ �& � �� ���%�8 � %�1 � �2 �  ���8 �8 �3 � g� ���X� ���� � !� � �	 �  �� ���� � %� � � �  ��� � �
 � }�� � � � ��T ��� )� ��`� �� ȱ�	 ȱ�
 ȱ� ȱ� )
����� 轡�� � )0� ȱ����H Ȍ � � �
 � �Lf�  Q�� �� � �� ��Ȍ � ���! �"�$ ȱ"�% ȱ"�& ȱ"�' ȱ"�( )
�����) 轡��* �( )0�- ȱ"����H ���T Ȍ! �+ �, �& � �� � � �N )����� �.  g�`�. �/�1 ȱ/�2 ȱ/�3 ȱ/�4 ȱ/�5 )
�����6 轡��7 �5 )0�: ȱ/����H ���T Ȍ. �8 �9 �3 � Ц� � � �N )��@Е��� �!  �퀈� �� ȱ� ȱ� ȱ� ȱ� )
����� 轡�� � )0�  ȱ����H Ȍ � � � � Ъ�  o�� �� � �� ��Ȍ � ���J 
��u��L �u��M �L� ȱL� `�J 
��y��L �y��M �L� ȱL� `H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; � �8�� �� )0� Ȍ ����� � � �; � z�h`H�Z� )?	@�; � I��-; �; � ��� )@��J��; �; �  �8��  �� )0�  Ȍ ����� � � �; � z�h`H�Z�' )?	@�; �' I��-; �; �, �)��( )@��J��; �; �- �8��- ��( )0�- Ȍ, �)����, �( �, �; � z�h`H�Z�4 )?	@�; �4 I��-; �; �9 �6��5 )@��J��; �; �: �8��: ��5 )0�: Ȍ9 �6����9 �5 �9 �; � z�h`� `� `H�Z�H ���%�I ���H �P �I )?
�����R 轻��S �Q  f�z�h`�P �* �G `�Q �R�C ȱR�= ȱR�> ȱR�D )
�����@ 轡��A �D )0�E ȌQ �? �B �C � \�T `H�Z�P ���LU�= �F �C I�F )��F �B �@��D )@��J��F �F �E �8��E ��D )0�E ȌB �@����B �D �B �C )�; �I )����
�@����; �; �F �( �; �G ��* �G �? �? �> � f�z�h`H�Z�  Q�  o� � �� �  }� �� �� �� )��� z�h`H�Z� � �
� � ��O �N )?�O �Q�� �K�O 
�����" ����/ 轕��# ����0 �! �. � � � �N )�����  g�N ���  �� )�z�h` �<�!B ��!@ �<�!B ��!@ �<�!� ��!� �P�!� �<�!B ��!@ �<�!B ��!@ �<�!B ��!@ �P�!C �<�!B ��!@ <�!B ��!        �!� ��!� ��!� �!� qP�!� (�!A _(�!A q�!@ ��!@ �(�!A ��!@ ��!@ ��!@ ��!@ �P�!C     � ���!� ��!� �P�!� �(�!� �(�!� �<�!� ��!� �<�!� ��!� �<�!� ��!� �(�!� �(�!�     � ���!� ��!� �P�!� �(�!� �(�!� �P�!� �(�!� �(�!� ��!�.
�!� �(�!� �P�!�     � �� � �� � �4� � �4� � �4� � �� � �� � �4� � �4� � �4� � �� � �� � �4� � �4� � �4� �     � �� � �� � �� � �� � �� � �� � �h� � �� � �� � �� � �� � �� � �� � �� � �� � �h� �     �.4� �.� �� �.� �� �� �.� �.4� �.� �� �.� �� �� �.� �.4� �.� �� � �� �� � �� �.� �     �.4� � �4� � �4� � �4� � �4� � �� �� � �h� �     � ��� /���     �     � /d���     � w!� w~!� w}!� w|!� w{!� wz!� wy!� wx!� ww!� wv!� wu!� wt!� ws!� wr!� wq!�     �	
	 �
	�
	
�
�
�	

	�
�
	�
	 �
�
	 �
	 �
	
	 �}���������q�  ��%�  s���  9���  ��������w���������������������0�Z�����������%�,�_      H   H      _   ?  !    _   (  ! 8      �"   o   �_2    �o� �Od    E�����E�����E�


(
.@

G
RZ
cd
�
` ` ` ` `  ` $` (` ,` 0` 6p<` @` D` H` X` \` `` d` l` p` t` �` ` 	


` 	pd
(
*` 	.2` 	:d
@
CpGHd
RX` 	Z
cd
f` 	jpnd
{d
 ��� �@��� ��� �@����� � � � @ ` P�� ��� ��� ��� �0� �@�P�`�p�������������ЇP�ЈP�ЉP�ЇP�������������ТP�УP�ФP�ХP����Њ��Ћ�P���Ц��(�P�Ч��������x�����P����Ќ�� GAME OVER $PAUSE$LEVEL  $HEIGHT :$READY  $HI SCORE$SCORE   $CONTINUE$END     $MAINaSCAN$VERNIER$POWaLEVEL$MAINaENGINE$ALLaGREEN$dddOK$GOODaLUCK$THEaEARTHaDEFERDER$BROKEaDOWN$THEaENEMYaAND$DEFENDaEARTH$STAFF$PLANNERa$aaLOUISEa$PROGRAMMERa$MUSICa$LIaWEIaXIAO$XUaHUIaHU$PICTUREa$YONGaBAN$LIaZHANG$TESTa$YAaLINGaJI$2�>�D�L�U�]�f�o�x������������������������!�(�4�>�G�P�Y�_�����  0@P`p��������  0@P`p��������  0@P`p������������������������������������������ 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          Z� �x�