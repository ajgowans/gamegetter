�?�&���q� ?��-
��+����,���l�  X� À� �?` � � � ���Ǜ3�ި������������)�
���|����`��Х����������	8�
�� ��`� �����������`�-��������	� ��� 
����`��)�摥�)�Ƒ��)�搥�)�Ɛ`��JJJ�P��B�3�E�2���� �2��P�� .����EeP���2�B�3��)�J��,����� ���2 .�������2�2�B�3�� ��2���� .����` ?����#����8�T������ �����������`�#� � ���2�`�3�!��� ��`�P �`�#���� �ey���f�@�g}��h`� �ei�f�@�gi�h` ��)�� � `� � `���h�6�-�B}H��B�
�8�
�B�A�A}M��A�
�8�
�A�@栩�� �����`)���M�1��JJ��R��1�l��0����P��)�� ���� A�`�-�M��PLD��-�H��PLD��-�P |�`     MMMMMMMMMMMMMPPPPPPPPPPPPP��������������������������         ��4擥�0. Yĥ�JJ�����晥	8噅	�����	� �����-��` @��P��1
��)����*���� ����P� ���������2������ .��P��`��P� ��2���� .��P��`/���O� ���  � ��[����}������.����;}����~��fT����UT���nAy���Pz���V�f���Y����j����������~��ޛ����m�f��y|���=�}��o/��������W� ���  ���                           ��   �  �g�>  �  ��� ��٫��W����k���k��U�z��f������� �j��  ���  ���?  ���   ��                                                          �/    ��  ��  ��Z  �E.  ��9  ��F9  ��V.  �~i  ���   ��   �/                                      �n�PʆQ�R� 
**���H�R=�� 
h(*=�
�
��P��`�����?� ��� 
�Ă��� � 
��)��R���n�n ߄� � 
���Ă��� 
����e����懥�i0����Ɓг`��@ �¥�9������� ��������� ��� ����@� @���2���3�`�"`擥�� ϐ`� ���)� �`�� �`�� ��`�� j�`�� &�`�� 9�`��� ��`�C�3�҅2���� � �Z��2�ȽZ��2� .�ƙ��C�3�܅2���� � �j��2�Ƚj��2� .�ƙ��E�3�N�2���� � �z��2����� .�ƙ��` � [l�5�6�ְ� � ���p6�6���� ��l  ?�  �9� p�0l ��G �90�p� ���Z��p p�p�5 ��իu�p L�p�6 ��Z��p Lp� 7 �6�~��5� � p� � �6l���5� � p�: ���:�U�o�:��� \�F�3�ʅ2�N��0�O��1���� �0�2���� .å0i�0��1ƙ��`P��  ��: �ۼ����?�00� \�  �0�?���[S��������O�����8��?�@3lWuۯ@���ٟ�4� �:O ��0Mm��k�E ���ٯ�v0T��� ��rDym��i�A���i�6v��6�  p���Zy���i��?���i�vvM���w9  ����j靭�������zڮvvC���  ����k幱����k�{��NnS��o  ������z��v�:�����������  ������z���y�?�{^���������?  ���O��{3�w�޷{�T��������  �����{3����{�S������z�� �I�3�
�2�Ԉ�0�Ո�1���� �0�2���� .å0i�0��1ƙ��`ֈ���_��{3���=|�C�����n�z��C���~O�w��ON��=����������W��L�_w���?N�W3����Z��z����Wz?L�W����M��������������W��O��G����M�C�V����������_��N�_9�[:T������?�����_�j5�e~�=�[N��W��U��;������_�:���~?�[^������W�;�W������?�e���?������������w��������5y����~��������������?�y��j���W�����> �����O�y������������~�� ��K�3�L�2�
��� � �I��2����� .�ƙ��`�z�����y��_�Ӕ�����~^�;�y�;��_�����S�������7�����_�����S:u�����7���:L�~������S:u������7���:ӗ��_����S�]�o���?<��:כ��������O�^�����><��6כ��g�����O�o��V��>{��6׫�������O��꫟�^�{��6ׯ��g�k���O�����y�{��6l�o����]u�S���ڜ�y�M�3�+�2�m��0�n��1���� �0�2���� .å0i�0��1ƙ��`o��y��6����_���nS��z�֌�y��M���p�j����޷ە���^5�y��Nn޶����_֞���������y�pNn����z�{����?���_��N~zvpNn���N�ۯw�N���]�>�:~zvpNn�m�Nyn����W��W��:~zvpNz�m�?]�P��U��[� �9z^vpNy�m �\�U��U����9y]upNy�m�����_W�����k�99u�9mm0������뿮:�6�99u�99�kL>�������������]�99����������� |��M]�O�3�p�2�
��� � �ʌ�2����� .�ƙ��`�< C���?��o1 ���P��k�C���     �T������    ���9�Z���Z    ���9ܫ���?   �п�:l�_�\��   �����<�  ��6   �?   �   �=        ��    �        �?  �O�3�l�2���� � ����2����� .�ƙ��O�3���2���� � ����2����� .�ƙ��`;�7������������1��p�zp�z��~�����;���?��s>|�w~}�{�~�������NGݧ_GݗOGۜ�[;\�[;p�[;������������l�;���?>|�s>|�w~}�{�~�����ϥ��0��)����$�K�3�V�2���� � �t��2����� .�ƙ��Ɵ`�Ye�[��[��  �  v�  vq�M�PS��]\5ut���s�N������?7p����W �� �� � ?� � ю }� À� �?`��I���E���A��)�;��JJJJJ)�0��c����k����[����T���������1���s��� b��ƚ��`���s���������V��� b�ƛ��ƚ��`�^��������V��� b�ƛ�`$&          Jr^6�Jn\4���q���m��ei�f�	�gi�h�	��������a���b���c���d �¥�/ƚߥ��2������)����ay摅b��cyd �¥� �é ���`��ͩ@�a��b�\�c�c�d �¥��`L<DlTs�S{k"::<":MMG �����#���  ����	� ��� 
����� ���� 
����\�����I�� ����`��)�����P�8�PJJI����Ś��JJř�ܦ��I�P��8���JJ��������� ق`  8Ph��hP8  8Ph��hP8 ,,,,,DDDDD\\\\\�� ��� #�`�� ��`�� ��`���!�!���� �#�#� �
 y� >�ƙ��#����`�#����;��� �� �� �� 
�L7��� 8�;���  W�`���/������!����ay摅b��cyd �¥� �`��թ��������a���b���c���d �¥�Pƚߥ���@�a��b�\�c�c�d �¥�1�@�a��b�R�c�[�d �¥��R�a�e�b�R�c�[�d �¥� 0� W�`          Hp8((0,0�@Ow�����?�$0<FRRR#/;EQcc[����Q�3�P�2� ��2���� .�ƙ��`��)���.�$�d��� ����JJJJ)��w����6�� b����� b�������`$&$���F >���)�
��:����������Q�3�P�2� ������ڒ�2��ƛ����� .å�i��ƙ��`��������� ��  �`  �    � *���*��jT�jBdBE�VEj��j��* �*�������ʓ����)��� @����� ��2���� .�����`��������� ��2����� .�����`������ �S��2����� .�����`������ �ӓ�2����� .�����`������� ����2����� .�����` 0`� (Px          @ @ @ � � � � � �? �� �� {� 4 4 p �        
  
  
 �? �? �� �/���p� p� �5          (  (  (  �  � ��0������A�A �  <  P  P  P  �  �  �  � � ���2��:�^;   \ � � p 4 4 {� �� �� �? � � � � � @ @ @   �5 p� p� ����/�� �? �?  
  
  
        <  � �A�A����0��� �  �  (  (  (        �  \  �^;��:��2 � � � �  �  �  P  P  P  ?   ��   \�  ��V ��V \�  ��    ?    �   �+  p�?  ��Z��Zp�?  �+   �    �   �  ���  p��jp��j���   �   �   �   �2   �� �A���A�� ��  �2   �    �    �  ��5 ��� ���  ��5   �   �    �   �>  ��� T��AT��A ���   �>   �   �   0�   �^P��P��  �^  0�   �    ?   ��  �z@��4@��4  �z  ��   ? �����	���� ˖`������)��������� �� 
� � ����`������������햕�T�����`4�����y����y����� 
�` �             ��(�a���b��c�c�d����ei�f��gi�h �¥�����`������	������`�������`���`�����
���`���`���	����`���`���������������������������������������������������������������������������������������������������������������5����6��������� &� �� O� �� À� �?`��� ��`� ���)�
�������#�!���
����i���i���iz����� @��2���3�� � X�` HX<TQTTRFBBBBB���D�!�@��� �#�#� �- y���i�a��i/�b��i�c��i7�d �¥� ؘƙ��#����`��i�ci�d �¥�`��i�ai�b��i�ci�d �¥�A��i �ai�b��i�ci�d �¥�"��i�ai�b��i�ci�d �¥� 0� W�`��J���F��ai�b�	�ci�d� ������}���e}���f��}���g}���h �¥� �é ���`晥����`   .00 ���Q擦����R�� a�`)�>���ƐƐ���(� y�`��(桩���`���摥��.��`�����摥��f��`����ƑƑ���/��`��ƑƑ�����`���ƐƐ���^� y�`�C�ǩ ������`��  �����7��i���i�)������ @������� ���12�2����� .�ƚ��Ɵ` 	  � � �? �擥��` �����H�����I�� ����`)����� �JJJ8��P��� 9������4�$JJJ�P�P�P��	�� 9����$�JJJ�P���� 9�`�� ��`��� ��`                ����}O����}X�� ق`�,�,�,��**�*������)?� ��`�� y�`��i����i:�������� b���i$�� b�`��i����i0��� ���������� b�Ɓ�`$&                                 ���          ��^�         ����        �����?        ?����        �����       ������      ������    ��������  �?l�����O9�?  O�lQ���_A9<�  O�lA�k�Z�<�  ��l���j�|�  ��|���j���  �:ܗ��j��p;  ��\��������  G�9��O����  �9y�?����  �9y�8����  �99�����[�  _�9���k�  ��p9��Զ9�>   ?�9��Զ��    �;-����      �>-�����    K;m�?��  K��K���  [��
��{�  [�<k���  l� �� [�  �� �9 [:  �� �? [�  K���?��  [�0��:��  [90�<:{�  l�0�<:�  ��0�<:[:  ����?[�  K� Ǐ��  K� ���  [9 L� {�  [� L� �  l� 09 [�  �� 09 [:  �� 0: [  L� � �;  L�   �9  \9    {9  \�    9  p�    [  ��    [  ��    �   �    �    �    ;    �        �                          ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������7����8��� @� �� !� =� À� �?`� ������
��?�(�� ��`����.���0�()�$� �������i����iK��������� b�ƛ�` o�`������"� �������i������������� b�ƛ�` F�`     )*$&���)��3��
����� �������������}&������#��� b�ƛ���ƚড�3��/���� ����i$������}&������ ��� b�ƛݩ��ƙ�`"*&%?      ���: ����0�1 �����|�����݅�� ��ݎ����)��桥��	�� �����|���`
L���LLUUUU���!�!���� �#�#� �
 y� ��ƙ��#����`��i	�ci1�d��i�ai�b �¥�A��i�ci�d��i�ai�b �¥�"��i;�ci�d��i�ai�b �¥� 0� W�`��~���z��ei�f�	�gi�h��i	�ci1�d��i�ai�b �¥�>��i�ci�d��i�ai�b �¥���i;�ci�d��i�ai�b �¥� �é ���` ��� ���H�����I�� ����`��� ����3�����P��}����8�� ق�����P��}����i� ق`����` $%&12>3333   �� ��� ��`�� ��`�� ��`擥�� $�`� ���)��擥�)���}��������}������}������ @��2���3������
�� ���)�� ��` 4  ���V��i;���i� @�� ��� ����� 
������ � 
�n��)�R� ߄� � 
�2���� .å�i���0��ƟƟ` �ک  ���> ��ޭ� �C�[� ��� �	�       (  
                                   �         �        <p      ��      �y�      �^�      ��_� �    ��\^�9    0:]�]    �8�n�     �k�      L5�9     �S?��    ��0��   �?5[��   �� Mn��    cOMn>9    �vMnC   �?��n��  pͬ6[�^  �N�6���    O�?��>    l�0כ    �Mn�   ��CM����  L? MnY?4  0�Mn�@  ��vMnd   ��NnC�    O�zg�6   �3��U��?  \ç�e�{  �U:�V�  �N�?���    o�0[�?   ��>5���   ��M���   �@Mnj�  L�@Mn�O  0Yuk=�   ��yu[C�   ����ZS�   �N�:���    ��O��:   �[��֪>   �k=�j��   ��C:���   P5�Z    [@9[�6    �M^�7    �<M^�    l�M޴    ��Nޭ    ��zW�    ܦ�V�    0k��     ��      ���>     ����     �o�[�     �����     ���      ��.      �k�      �\�       �O�       pM�      ��      <??      33       �        �                                   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ٮ �� � � À� �?`���������ei�f�	�gi�h������ �ai�b��ci�d �¥�>��� i�ai�b�i�ci�d �¥�ƚ��T�a�k�b�@�c�_�d �¥� �é ���`��JJ)���2�ڨ�3�:��1�9�}ܨ�0��1�� �0�2���� .å0i�0��1���`LO ` ��?  SO�� ��PV�05�U]�TV�5L�U[6C�W֖�S���f�W�����W��f�[���[�}tf��x�:���8�:��}4�?\����:�Z�A�����W꾾�霾�:�ʫ�������ҫ� 뾾�  ﾽ� �����������K���pk�<ܯ�;<��?;� ?�3� �P�թ��P��� �٩�2����� .��P��`� �y��2����� .��P��` P P �?   � �  0TU ee5 \�m� [�� ���� ���� ���:  ��  �    �    <    <    0    ��   <   @0 �PU1 p��� p��Ul��Z���j��������  �?  �   p   �    �    �     �  � <   �  CU� �QVV�U�V���j���������?��  ;�  �   �   �   �        �  ��  0  U GYY Wy[5����5����6����: ��  ��  ;    7               @��� ��2 .����` @�� ��2���� .�Ɲ��`�����"0� ��� �Lg�� i��� ������0��� ��� *�`I���杽 ��i8坅 *�`�@��� ���T���&�� b��$�� b��l����� b���� b��\���&�� b��$�� b��d����� b���� b�`���;��)����1�)�*�JJJJ)� ��������������������� b�ƙ�`��'��������������������� b�晥���� ��`������ ���^���$��������� b�ƛ�`���������������� ������������ b�ƛ�暥����`�^.<T$T22$&��)���0F�����)������/���� ?���� e�� �)�P�e��� @� ���晥����`�  �   �  ������������������������������������������������������  �            �  ������������������������������!�!���� �#�#� �
 y� խƙ��#����`������ �ai�b��ci�d �¥�X��� i�ai�b�i�ci�d �¥�5ƚ��T�a�k�b�@�c�_�d �¥��Z�a�e�b�X�c�_�d �¥� 0� W�`���@�$j� )�� 8���8����JJJJ)�P ق`�`�*)����)JJJ�P���T��8� ق���P�T��P� ق`����I�� ����``�� ��� �� R�`�� ��`�� ��`擥�� ��`��)� �� �� �`���,��)�&�M�3���2���� � �$��2�Ƚ$��2� .�ƙ��Ɵ`����        ��[��E�B�C�B�.��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ����	 ^� � � À� �?`���9����3�������օ�`ɀ� �`��� ������N���X�� b��d�� b�`�0���� ��`�P���� ��`�h�� �� ��` ~�`��ɠ�3)�/��JJJJ8�
)��అ��N��� ����������ڰ�� b��ƚ��`���అ��N��� ��������ڰ�� b�ƙ�`&$\Jn\����������N�������� b�ƙ�`DPht擥�� 3�`��� ��L2���)JJ���� ��� �� �� ��`�� ��� l�`�� ��`�� ��`��)�$��JJJ���������i��ԅ���P قƚ�`�����������҅�ԅ @��� ��2 .������ ��2���� .����ƚ�`��)�-��JJJ8���豅��������� ��P�$���H�� ق�ƚ��` 
!#         <<l<l<<l<ll<l<<l<ll<lT<lTTlTTTTTTTTT888888$88$$8$$$$8$8$8$8$$ ����� � O�`ɀ� ��`����I�� ����`��ʽ�3�ﲅ2�粅��벅��<�}���1�;�}���0��1� �0�2�ę�� .å0e��0��1ƚ���Х���� ��`
��!CFHK ��n  ��)�� E���
��m��0�n��1����ѵ҅�ԅ @�� �0�2���� .å0i�0��1ƙ��`�ѵ��$�� 
��Ѥ���yp��ҵ�yu���� � z�` ó`   � �  �������w����`�����Y����`�%��� �օ�`����� ����`����Ʉ�۩��`�������Y����`�w����`�����%�� ��`����� �����`����Ʉ����`�Ѧ��� }3���� }8�� @��ѵ��� =�` P�`      �� ��2���� .����`�� ��2 .����`���!�!���� �#�#� �
 y� ��ƙ��#����`�������a����b����c����d �¥�H������ }��a}��b�� }��c}��d �¥�ƚ��\�a�h�b�J�c�L�d �¥� 0� W�`D8Dlt�S{?? >QQ   
     ��q���m��ei�f�	�gi�h���������a����b����c����d �¥�/������ }��a}��b�� }��c}��d �¥�ƚ�` �é ���`L<DlTs�S{k"::<":MMG���,��)�&�I�3��2���� � �յ�2�Ƚյ�2� .�ƙ��Ɵ`)h��              �)h��Y�YiUY �� @ �  �2 � L>  k � 0� � � ��� `
 �Tl<`
<�T9l��3p�3Z9[Yp2p�e�kV]|>pv��U�w�p�U:�֕�u�sf��z%�u�s���^&�u�Ù���&�}���� �&{���� ��&{���k��&{���op�&{���op�&<{�|ٯ�?  \��0�\ֿ5  �?0� ��[2��ճ6 �W�< �3o2����6 |y��� �3o2_��=�� �n Sj�?o2Wڜ=����o Sj_�o��k�=�����  S����orի��Z�?��  �گ��orի��ڵ���  �ڮ��onU��mvm:��  ����j������kΟ� ����庚WV��魛�_o�������U�ij���_n������y_�V����n�3�����^W�k���R>p��?�����_U�����V���Ci���WU.�eڭk:���Wj�~�W���շ�:���j������Vڷ������ ��[������ ���� ��W�����__� ���6� �ח����ZU���6��P������ߪUU0\�\��Z�w����ޫf�?p�� �keWe���ֿ� �� ���^Y�kf���� �P��]Y��f���U0U�j}VY�����VL����WYi���j1L��> �UY> ���5��? �V�? ���֓�;  �V�?  ���:  �[�>  ���<�?  8[�,  ��<� �  �_�  T0Dj �_� ��0Uj  ~�  �T�0Uj  �  �T�<�k      �ԯ=��3      �?��WT5      \P��}�7      ��}ߧi�2      ��i����      ���?q�J�  �?    ��?   <U�  �jU� 0��j̰�(�Z̰�j1��<�5L�?  ��0� ���T0 0� ��� 0� �j�� �?�� ��� � ��  � ��   � L�   � L  � 0  � 0i  � �d  � ��1     S�     L    0d    �C�     <    �S�     �U?     �   �    �W�  �W�Z=  _��[ �����p鯾�7\����7��<��5��  �_6�; �W�� ��j��U�� ����� ���� � � �� �   �6 �   �6 �  ��6 ;  �� ;  p� :  pn :  \o   ��   ��6   p�    ��   �>    _�   �?     �            ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��� �?�q�A��=� ����0$��
 ����0�����
�����6����7 b���
��� �ɰ`� ����0,�� ��n����o�@��`����3���2 �� �� $� J���� ��`e�e�e�e�������΄$�z�Ѕ�N�Ԇ�;�X�����#�N�y�ǈ�`����-�l�"�������΄$�z�ԆX�����#�N�y�ǈ�`����-�l�"����������������������������������� �S)��@�S)��@�S)��`�S)��`�@��ɰ��`�ɘ�  �`������`l6 �� � )�������������� � �`�`i�`�@i�@  �`�� � )JJJ������ �S)�0�S)��S)��@�@ɠ���   �`�@�@���� ��`8�	������@�� `�� ` �� � )JJJ��^���� �R)��@y`��@�R)?i ��`y`��`  ��� )����; ��`!�������������������� ��� �  �                    �  � ��� ���������������������� � )JJJ��X���� �S)�+�S)��`ɏ���� `�@�@�Z�
��� ��   �`�S)��@�@ɟ�쩘� ��S)�� Z��� ɀ�ө� ��"�� �R)?��R)@��@y���@�
�@8����@�Ri )?��R� ��`��`8����``�`y���``     � ������������������������������ � )JJJ��9���� )�$ ;��� � ɀ��� ��� ��; ��  �`� �0����� �� `#�� �R)?��R)@��@y���@�
�@8����@�Ri )?��R� ��`��`8����``�`y���`��``    �  �  � �� �� ���� ������������������ ���� �� �� �  �  �    �� � )JJJ��"���� �S)� a��� �@���   �`�@�8�ɘ���; ��`ɐ�
�� ��� `	$�� � )JJJ��x���� �S)� a��� �@���   �`�@�8�Ɉ���; ��`ɀ�
�� ��� `
%�� � )JJJ��΅��� �S)� a��� �@���   �`�@�8��x���; ��`�p�
�� ��� `&�� )��`�(�
�� ��� `� � �1���:� �; ��`�Q��� `�� )�"�`� ���:� �; ��`�x�"�� � � `� � �1�����Q��� `�� � )��`  �`�� �R)��R) ��@y���@�
�@8����@�Ri)��R���0��`8����``�`y���`��``  � ������������������������ �  �� � )JJJ�������#�@�W�� ��;������: �������`'$&"*)��`ɀ��P�� �� �;�"�: ��`��`ɒ��h��8�� �;��: ��`�� � )JJJ������� )��`�@����ɨ��� � )��@L���@  �`(�� � )JJJ������� )� �`)�� )JJJ��!����`�$�8� � � �� � �;��: ��`�� � ���@�`��� `�� `�@��� �;��: ��`*�� � )JJJ��L���� ��� � � I� `+�� � )JJJ��w���� �(�� � � I� `,�� � )JJJ��ň��� )0��`�H��� `���`�X��`�𩩝 `�`�0���; ��`-�� � )JJJ������ )0��`�8��� `���`�@��P�𩩝 `�`�(���; ��`.�� � )JJJ��^���� )0��`�(��� ����`�@���� `�`� ����; ��`/�� � )JJJ������� )��`���(��� `�8����� ��; ��`0�� � )JJJ��䉝�� )��`�(��8��� `�X����� `�`�0���; ��`1�� � )JJJ��+���� )��`�8��H��� `�`����� `�`� ���; ��`2�� � )JJJ��"���� )0� �@�Z���� �� `� )��`  �`� �� )��`  �`� H������ h)�� JJJJJ)��$��:� �; ���� H)?�PI?�h�@��@y,��@�P�`8�,��`L�ɀ��`8�,��`�P�@8�,��@L�����@8�,��@�P�`y,��`L��`y,��`�P�@y,��@  �`3*"&     �  �  � � � ��� ��������������������������������������������� � )JJJ������� )��`�x�
�� ��� `� �I?H�@y⋝@h��`y⋝`  ��� �����#��/���; ��`�@о�� `4   �  � � � ������������������������������������������������������ � )JJJ������� )��`�x�
�� ��� `� �I?H�@8�⋝@h��`y⋝`  ��� �����#��/���; ��`�@о�� `5`�� � )�� JJJJJ)iC��`���/������ 0 �� �L匽p���� L��&�� � ���`���P�^���� ��`�0�^����p����P�3�`�2� ��2����� .æ��3�P�2�`�0
�����0����1�3�^�� �0�2����� .å0e��0��1����`���&����$�d�����T�d�t����������� � @AJ�)D�Y�ZdAJj�)�E��Y��ZdAAj��E�P�Z@Aj )   @@ P TATVeIA�fD@�U@YVAe�EDYUEdYUdVV���@�f T @U        PQ  PX�  @aM @��5	  A�  iX  �a  D��%  $A  �i �� @J�  )T�  @I  T Y    �    T     T @�VPZZ�ZUdVYU��ZETUYUUUAD�UUY ETY Q@DT   D   @ 	 PPAPU@@P Dd � D�QY`dj@�YUeDUP@U@&  �    ADBADDP E D R AT@!e�PD!RE�Q!e�AA EThPPT@DA�UDDiJFTV�Y��Vj���T��Ye�ZY��TYiA �fV TZE @    T T @T P TP��ZAAfTQUUUQTUTUdTEPiTAU�U�P��@)j T  P @UTPEPTUPT PQ @EUTUTPQ@U P  P @�Z�
�dPD$QIeIDQdIEEdEEaEEaQQa$UTdU��@�Z P  @@Q@AETA@PAA   A @@@@ AA@@ AV PT $`T T @U AEP A@AD@ @  P    EPP  @P��  TQDPaUU�TY��Y���iP�Z  �  T    @   PU@  $ P @ �TDDiTDI�ZQ�vUD�U����e�A����VBUi�iDATj�iAQ՛�eHQ���VID���YD�WgiDQ�Z)DYZYPdUU%@�X� PP  PE   T  P Y@�QTF T QPAYDP@DiDeDdDdeDDT�d  ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������q��%��$�%)� ��` D�`���'�'� ���
��ߨ�.�ਅ/ ܨ�'�&�'��`��8�&��� ��`�����%)���{��` j��&���%�2� �$�+Ħ������ �&� ���� �&L��� �������`� ���� ��䦐�`��`l. y�ũ��5���ɪ��M���ګ�v����P������S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S���R�8��P�I��P�P�R��S�8�	�Q�
I��Q�Q��S�Q���R�(`�P���S�(`�ReS�(`�'���-��������( �©��������( �¦'� ��'����� �� ��`� � `�'������Z���� �( �¦'� ��'����� �� ��`� � `�'�����������( �¦'� ������ �� ��`� � `�'���-���O������( �©���������( �¦'� ��'����� �� ��`� � `�'���+���	�������( ����i ����'� ������ �� ��`� � `�����p�����( �¥i����'� � `����� �����( �¥i����'� � `�'���)�����������( �¦'� ���`� � `� ������{����������( �������'� � `X���XLL�������'���
��������� ���������( �¦'��`�0���'� ��� �� � `�'�����������( �¦'� �������� ��`� � `�'������ �L���a�� /� �¦'� �������� ��`� � ` ��hH00Hh������ =[y������y[=� �������(����� �������'� � `*Br���'�����6� ������(�� �¥i���( �¦'� �� � `��`�0���Н�п jjj:::���RRR"""�'���.� �G�������(�� �¥i(� �¦'� �� � `�����(�� ��` $8L`t����� ���|������( ��������'� � ` 8P��� ����������( ��������'� � `p���'����������(�� �¦'� ������ �� ��`� � `�'�����������(�� �¦'� ������ �� ��`� � `�'����������(�� �¦'� ������ �� ��`� � `�'��8�JJ���������(�6� �¥�/��'� � ����� � `���� `�#��� `�� `8Xx������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ O�� �� ��������-�{����-
�����J����K����L����M����N����O���J� �L���N����`�-������



�� �� �@�P�۰iJJ�`����0�+��p�����`
     �   ���	
	
������X0xp0P0HpP0Hp0PpH0pHp0x0p0x�p0P0xPH0p0Px��xHP0PHPp0PPp�PpH0pPp0x������(*5ACGfk %),2;>FIS`o�%?CIOXZdgj��&+.8>[\]_`c�$'(?AFM������skiX���z���������(�U����R�����`�� � ���� � `�@� @`��  ```�` �� @`��� `� @@����@��  ���    �  @`� ��@�  `���  `�� @`���  @`��� ���� ��@`� `�� @`��� ���� `�@��    	
      !!!!!"""###% 
	
    


"    &!'    '!&
		  

" "

&

&		         $		"		



&	
   

    	


     !!!!"""#####$$$$%���@� @��� `� �� @���@�� @��`` `� `� � @��@��` @� `� `� @��@`�`��@� ��`�  ���@�@`�@� �`�� @`�� @`�� @��@��@`���@`���   				

   !!"""###$$$&@`� `�� `��`�� `��� � `�� `�@`�  �� �@�� � @�� `�� `�� �� �� @� @���  `�� `  �@� @��  `�@  �� �� � `� �� @�@
    
#		
  

	
	
"		   
       				


    !"""###$$$$%@`�� @��� ��� @��`�`��@�� `� `�� ��  � @ `�  ����  ��@`� ` `� `�@����` `�� � � `� `�  �ࠠ `��   ` �� `���!




$	!	
%#   	

!
'


     		

  !!"#####$$%`���  @�� @�� `� ` @��@� �` ` ����  @�  `� ��@�@`���@�`@  `�� ���� ` ` @�� ���@�  `���@��%


   
$  %	$&&"   	#

	! ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������%�j)� ��L���	�i�
� ��j � �ʩ �� �?�`��l`�@ UU}}�Ã��~��s�]ux��|�x x��x��x � x�����x �����x ���� x�x�x x�x��� 0 x�����x � ��������P�̀�1�ހ�0 A�晥����` LLLLLLLLLNNNNNNNNPRTVXZ\^�)��(� �@�A�B�C�D�E�F�G�k�<���I��H��=�m�`�P�3���2�i


��������K���� ��� ��� ����=5��� �2ȑ2�Lg���
��;��2��;��2�朥���� .�来�����ƚб�i`���g�)�9�����1���8��
i��0�D�1�8���
i��0�A�1��	��P A�����������������	�� ��`�� ` &0=Rjz!-5I]t
      
   
  � ��������P�R�1�
i�0 A�晥����`�)��ɩ�� �� �`� ɂ`���
�!� �D�3��A�3���2�� ��2���� .����`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������I '��� 9�� � ��L� ��� �� �?�`�����z��� ��`� ��)����PL^��)���JJJ)�P b�`�P����������������X�3����2���1���0�� �0�2���� .å0i�0��1���ƛ�`���p� � �@ ����"(��(�P"�T����� ��  R�  B�  B�  H&  H&  H!  H!   	   	        �  �  �  B� �P P V��R�
��
�T
�R� ��  R�  ��  ��  �!  �"  H"  H"  `
   	   	  �  �  �  �  �  B� �P � �Z �Z � �Z �V d
�T�D�D�@�H�@ � �(��(����������� �         ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
������������Ð���Đ������@������������� ���� w��������� ����懥�i����ƃ������iX�����Ɓ����оƂ����ж`��JJJJe�����)



e�����`� ����Q��P���������P��i.�����Q��`ǐW��� ?  F M   FM M M F  F    F M M    FM?    M$+29@GNU\cj F  	%,3:AHOV]dkF  1
&-4;BIPW^el  F  '.5<CJQX_fm M  !(/6=DKRY`gn ?F")07>ELSZaho M  F ? M  F ? M �MF  F ? F  F M F M#* FF  �s  MFF? F ?   FM tx|�������� M FMF M{uy}�����������M F8ivz~��        ���� prw  ���� �����  ���q                 ��     ����������          ����������         T[bb� ������                        **************************************************************sty*****************uvz*****************wx{******************************************)5************* *46*GR]e********"+7@HS^f********#,8AIT_g********$-9BJU`h*********%.:CKVa**********	&/;DLWb**********
'0<EMXc**********(1=FNYd**OZkl******2>****P[mn***** *3?* ***Q\op*****!****!***ijqr*********************���������������������?�O�������������������������O�?�������������?�C?�O�Oj����ƤƤƤƤƤ��ZOj?��P������������������������� UTZ�j������?�CƔƤƓƓƓ�i�T�U� ��������  UU �������������������?���TV�U� ������������������������  UU ������������������1�1i1iFjUU  ��������  UU��ƓƓƓƓƓƓƓƓ�V��ƓƓƓ�T  ������������������������  UU�ƤƤ�d�d�d�d�d�d��V��� ������S��������� ?U0�œ�OOOO���d����<�C�ZOjO�?U? ����������������ꪮ�g  UU�����������������œƤƤ�UU  �������� �UŤƓƓƓƓƓƓƓƓƓƓƓƓƐ�UEi1T���������D�UA�O?D� �U�j������������������������??j@UU  �������� SU��ƓƓƓƓƓƓƓƓƓƓƓƓƤ�i�������������g�[I[F�A�P���� OU?������������������ĤĤ�iiFjUU  ��������� US����j����jS���PS���VT� ��P����������������j�f�UV�[�  UU�ƤƤ�d�d�d�d�d�d��V��� ������S������������V ��@�?����V�jũƤ�����j�U0 ������������������������ ���?�O�S��������������Ɠ�S�O?U� ���������  TU��Ɠ�O�O�O�O�O�SƓ���U�����U� ���������������o��������� U�i���������������������?i@��PU ��������  UU��ƔƓ������O�O�@�Uƪ�@OjOU �����������������������  UU ?�?�?�?��������O�O�O�S����?�O�?��������  UU�V��ƓƓƓƓƓƓƓƓƓƓƓƓƤUU  ������������������������  UU��ƓƓƓƓƓƓƓƓƓƓƓƓƓƤUU  ����������?�Y���ƓƓ������ƓƓ��Y�?�����������O8�?�?8�O��T�SLOL?L�L�O�O�O�O�O�O�O�O�O�O���T���������  UU��ƓƓƓƓƓƓƓƓƓƓƓƓƓƤUU  ����������?��?�?�?�?�?� �U�j�?OOO��������OOj<U� ���������  UU d�T1���������T1� U� �����������������������TP��j�������������������?j@��PU ��������  UU��ƓƓƓƓƓƓƓƓ�V��ƓƓƓ�T  ������������Uj�jZP ��������������������O�O�O�S����������������� �U�œ�OOOO���d����<�C�jO�O�?U? �����������n��A��E�����������������T PP�����������������������������﮾Z�V�EfUAV E@                        @A�U�������������[UED                                 @@UT����n�[�Z�[��V��V��U�D� � T QD @@ @D  D   A @ T@�T������������������������k��������f���e���d�UdQ P@�P��������������������������������jfU  UP�U�������������������������������������UU PU�������������������������V  U���������������������������U ���������������������������U� @�
����������������������������UU  �*����������������������������U� P�*������������U� U* ��������������U��� �*���������箧��z�e�U����������@�
T����������������Q���Q��_���������������������������P�I�'P�
�'��������������T���@����������������������������������A��k@���o������������������������������������ �����WUUUUUU�W�_�U�U�W�_UUUUUU������տ�_�W�V�U�U����U�U�U�}����U�U�U�U�U�U�U����U�U�U���������oUWUVUU�U�U������U�U�U�U�U�UU�U�U�U�UUVU[U���U�U�U�U�U�U�U�����������U�����oUWUVUU�U�UUU�U��������UUUUU�U�UUUUUU���������U�U�U�U�U�����U�U�U�U�UUU�U�U�U�U�U�U�U��UUUUWU_UU�U�W��������o��7x7s7x7s�o������������� ������� ����������������������������������������� ��������� ������������������ ����� ������� ��������������������� ����� ����� ������� � �������  ��  ��  ��  ����W�W������   � ?W�������������쵬��W�w���������������^�z { � � �w�w޻o{o�oOO�o]u�n_�u�׿_��������^�z����װ^p^p^p^�לל���m�m���U����������� � �p�                        � ��G�N�_y�yݾ�y�y���y�y���y�y��y�{���u���Z�o�������������_�_�_^�y��o�@ 5��\^�r���u�m�m�m�o������� { { � �@ ���(��P�T���� � R B B H H H H         � � �               � _���_������盓G�G曑G�G曑G�Gv�і�[��w�w�_�ߑ��ו7�5U5�5�7�7��@�@^ y�5��P� ^]�ysy_yUy��������������� 3 � �"�("�� � � � & & ! ! 	 	              � 3>0�ž�zo�^��o�^_�U�[� 6 � � ?         � ����:�:p�_�U�_�^��������8�8�8���� 2            7 7 7 7 � �                 �pް��  � W �{{1{���k�����>}O}L~�SzSz����w�w��� � � � � � � � � � � k � � � l , , l � � � l , l � � � l , l � � � � � � � � � � � �    � ����ps�]������ � � � � � � 7 7 ;7��u�������� � � : ���0�L:������[�k�|�|�1�ڬŬŻ��������?� � � � ; � �������:�?�:�9�8�8�9� ; : 9 8 9  ; : 9 8 9                        � 0 O���S�������n�n�����U����z W���� � �            �� � wv^^�^U^�v�vuv5���U�W�^������  �                     � �PUP_�z��v�v��������F�����Ɲ����F�F��F�F���F�Fכ�V\�\U\�ܪ�V����m�W����p]p]s}UU��������^�N �  ��S�LLLL00i�i�i����>�   � 0 L ���0�         ��??0@�կ���~m^mn�mmm�m9mw�7m9my�m�m~_][�ߥ{�{�_������o�o�_�W��W�^����AP@ �W��u�W������2�2�2�2�2�2��� = ; ;  � �  �0�ᰅ�nijj����o�l�������l���6�6���   � ?�@�T��ګ��۷������������u�]����u�]��������{�[�V���_��:��mmm����6�6�6�6�2�2�2�2�2�2�6�6��� <               ��?�@����;�;�;�;�;�;�;�;�;^;W;�:������������� � � ? 0e0i��p��?      �� � � � � �    � ��303Kϒ  �?�@ŐƑ1�1�1���������K:?.�.�1ffji���.>���9���pp�    1 � Z��       Yi�W�          ? �g�5��\V      ����pfp�pj�Z���   ��r���n����6���� � l k���� ?    �s��������       ���p�\6�6�5������    9 � �W�     ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`� Q���@JJe2�2��3�2���3��`��������������������������� Q��JJe2�2��3`�H)��n��2hJJJJ)��~�y���3` 0`��� P���@p��@@@@@@AAAAABBBBB 	� �R��`8�	�	I��Ș��R�P�@8��I��ȘH�Ri�Rh�Q�R�Q���P������	�PJ�Q�����:`(*"$&" �¥�*�;�� ��� �;���� �
�P
�Q����RJ�S�;� s�`���`ɘ��i�@��;���@eP8�;8�;� ������  @���2���3�`�"`���@eP8�� ��`eS8��@�� �����:�  @���2���3�`�"`� ���� �	��� ���` ̥��� � �(� `� ��f�a��b�e��h�c�
�d�g���`�� ��2ȑ2 .����`�#����R�P�Q� ��2��Q� .��R��`�2i0�2��3`�0��1`�PH



���Ph��� ��ԑ0����� g��P��`� ��Ց0����� g��P��`�P



���P� �ԑ0����� g��P��`�=0��<�� �=�
�� ��`�	�=�<�	�� ��` 	ɦ� )@� 3ɦ� )�� ��`�o�Z� � �n�[� 	� 
���[��� � 
��Z��)��R �ɥo�Z� �nȽ 
� 	����Z�� ��`�o�Z� �n�[�[� �2= 
 	�2���[�� .��Z��`���������`�k�{���	� @��2�
�3���A�� ����@�V�=<�� �i�j��k`��`�������	�	�	�)JJJ�����ą� ��n����o 	� �� $ĥ��>� ��` �M�3���2� � � �2���
�� .��P������-�� ��`� ���+ŅP�0Ņ0�M�1 A������` ������`����V�eE�E�`� � � ��� ��`     ��@�
�	�
�@�?L�����`��b��I� �`�`��06��2�@�ayƅb�`�cyNƅd�`���A��!� Ǧ`���� ���`�`� �� �� �ʥk����  �� �`                              �"�v��r��ai�b�	�ci�d� �\���@�g� �eytǅf� �	�gi�h��g�h8���g�g �¥�)��| �é �������"� � �`�3���2 ��`�� ��`� � �R���@�g� �eytǅf� �	�gi�h�
�g}��h�h �¥�!����!� � �`�3���2 �©�| w�`�� ��`�`���� ��L���6�� iA��� � ` 5�`� ����ǅ:� �;�`� �������`&"*��9��ei�f�	�gi�h �¥� �`���A�� �� � ���� �� 5�` 6ȩ�{ �`�`��������2���3���� ��2���� .�Ɲ��`�`���A��)��9�`�B��>�.�>`�C��)�!�	�`�D��)��)�`�H�	��H`�eD�D ��`� �Q�Z� 	�P�$P���Q�QP���Q�Q&P&P���Z�Q� 	`� @�n�Z�Z� �[�o�[eZ�[���� � 
�P� �Q�$P0	p��Q�Q&P&P��Q� 
��[��`0��
�� �4��5�o�Z� � �n�[�4� 	���[���Z��`� �Z�o�Zen�Z����Z ���Z��nJ�V�X� �W�o�R�W�en�ʹ 	H� 	� 	h� 	���X��Wen�W�V�X�R��`� �V�W�o�J�R��Wen�W����V�W�n�X� 	H� 	� 	h� 	���X��W8�n�W�Ven�V�R��`�o�S�nʆQ�n�P�Q�R� 
**���H�R=ʙ 
h(*=�
�
��P�ۥQen�Q�Q�S��`�����?�� Q��JJe2�2��3�)�	�R� �X �ɥV�R� �0�2��R��`�0�0����1`�2��3`�2�2����3`�0i0�0��1`�08�0�0��1`�28�0�2��3`��O� �������:)�� ��V�V����W���1���0� �V� �0���� g��W������������ ��` �˩��2�@�3� � �cˑ2����� .�� ��<�P�@�1���0 |å=�P�@�1���0 |é ���[˅0�@�1�@�P |������
�P���0�@�1 |åH�P���0�@�1 |�`��������    <<  ��<����>���<3�  0  �@Ũ�E��Aũ�=��BŪ�5��{�=�=�
�8�
�=�<��������i���
�8�
��橥��
��`�������`�������`� �����`��& �� �� u� '�q� ��  � S� Y� �� �ө �` Ḁ� ������ � ��@��`  � J��`� ���������`��� ��`������`�I�  ��  �`�k�T�>�/��3�
8��2��3��W� ��2������ �2��
�� .��W����̅W��̥
�2��3� �W�2�� .����`�)��ͅV��3�1�
i�0��1�
8��2��3��W� �V�͑2�0�����V .� g��W��` 0HUU }} �� �� �~ �� s� ]u TU�����5t�PU��0<0��0<0��U@U@_��0�`0@���0�\3@W� ���� �	��� ���`�)���ͅ���ͅ����	}�ͅ�}�ͅ��ͅS C��Ƣ��` ��������*&"��&� ��>� ��  Υ	8���
��΅8�΅9l8 `8�uΎι����-�\ϥ)�	�}�� �{`�}���|`�i���S ~ͥ�*���@�� � �����S�  @���2���3�`�!`�8����S CΥi
� C�`�i���S CΥ8���
�S CΥi
��	�S C�` �Υ8���*�S CΥi���S C�`���i���S ~ͥ�,���@�� �S�������  @���2���3�`�!`����Se� ��`���i���S �������8�� �Υi� ��`���8����S �Υi���S ��`�#����R�P�Q� ��2��Q� ��R��`�!�-� �#�#� ��`�3���2����P �L�� ���#�#� �ץ"�-� �#�#� ��`�3���2����P }�L�� ���#�#� ��`�#�S)�� �S) �� �S)�� �S)�� �S)��@�@�S)��@�@� ���ɰ�	�@�ɠ�� � �"`� @��#�2���3�`��P� )


�� �2=3�ґ2�ȱ2=3�ґ2� .��P��`�#�@ɟ��������B� ��� �"`�����gӰ��ymӝ��@yjӝ@L���@�@�@�@ɟ����@�@�� � @��#�2���3�`� )�V���R���� *�`�� Q�`�V
�V� �V�2=���ґ2�ȱ2=���ґ2 ��R��`�V��ӅV� �V��P�2=���ӑ2���P�� ��R��`�#�S)�� �S) �� �S)�� �S)�� �S)��@�@�S)��@�@� ��ɰ���@ɠ�� � �!`� @��#�2���3�`��P� )


�� �2=3�ґ2�ȱ2=3�ґ2� .��P��`< � � < � ��� ���� �?�?  � � � �� � ������?�  ?��!�#� �#�#� ��S��� ��Lr� x��#�#� ��"�#� �#�#� ��S��� ��L�� ���#�#� ��`�V
�V� �V�2=���ґ2�ȱ2=���ґ2 .��R��`� ���? � �� �#�@��������B� ��� �!`�����gӰ��ymӝ��@8�jӝ@L#��@�@�@�@��� �@�@�� � @��#�2���3�`� )�V���R���� ��`�� p�` (  �V��ӅV� �V��P�2=���ӑ2���P�� .��R��` 	�?��0�3���  �  �    ���6���3� ���	ԅP�
i��0�J�1 A������-�P�P�J�1���0 |�`�J�1���0�� ��0���� g����`    �<?�<?<<�  �������  � < <�  �?  � < <� < <�   ?�?�<<<<�< <  �?  � < <�  �0 �<<�  � < < < < < <  �<<�?<<�  �<<�? <<�  ?;;;;;;;;;?   < ?�?�<�<?<  �?<�?<�  �<0   0�  �<<<<�  �?  �  �?  �?  �?     �0 �<<�3  <<<�?<<<  �������     0�   <�� 0        �?  <??�<<<<<  <<?<�<?<<  �<<<<<�  �00<?�   �<<<�?<��  �0<�<  �?? � �� ?�  �?��� � � �   <<<<<<�  <<<<��  <<<<�<??<  0<��0<0  <>0����   � ?��� ? �?                ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��2��s�� .��t��`�u����ʽC؅v�G؅w�w�K؅3�X؅2�e؅s�r؅t  ��w�v��` ISJJJRLLLPMMM��������00  � �� � �� ���y�7�� �`�`���A����6�� iA��� � L�� 5��`�`� �ө�|`�q�k�r)�� � L��� � �r���y� ��!�"�x�r�M��B�Uمs�]مt�t�eم3��م2�
���م0��م1 ��t�s���x�r�r�p�� �q��  �`)���x����u ��r`  01@P`		  MLLOOJJJMMMPPPIIIILLLLOOOORRRR�������������]ڝ����]۝������]ܝ����]ݝ�����]�]ޝޝ������]ߝ��� P @�i�Z���edUU�D*eQii eY DYiEPi�D*dUU�Ye���@�j P   P�  jZ PZ TU TU  @j�%@e�ih��i �iiQ�VY�jZ@* �Y Z�j Z  ��  U� �� TQ @Q PYUZQ*�%T)fZ@j�jQi�e@�A� YA� ��f@ Z�fVPjAiFYA�Vi�����hPfPU�ePeA T dQ h�U �Ve  ��  P� iA� �F�PiA�QZPi�iTe�ZTe�&P&fU)UEU
EP�	 TZUQ U� e�
 ��  Z             P  @�  �Z  � @�U �V d YU  i @Z@@P U�i@d�@�    TUUU���jj��eU�QeVRT�TU @       EEUQE��U��U��j
  �        U   �  �  ie  e� U�	 QP) U�  @�  � @TPP VUP�dP���&�T)T)A	X 	hT	�D
hE
hE	TP*dP%�@$dUP�`A�F TA)XU)�T*hD)`P*`P%�@$�%�@)`P%hP�)h@)XUVP
�@��FT�V�j@@@ ZQ  �U  � �E @VF  �V  �Z   �   @        
  ���jY��Ue�QUYQTEE@A @    QQ�EU�VZ���f�VP�V     Z U e T�T� D� @Ei @) U	 QY D�  T  �  Z                          �  �F  �  V  �  `  X P X @    )� e�P����`P� �Y�ZU�E @        PQD�eT�iUYTVYdY�je��Z�j*h�U	�� ��  ��  UU�P@� @DT    EP UT Z�QAZ�Q��������*��j��   �   �            *   �  T*  @�   V @	  @% Q � TYDZPY 	Z `i`iX �X �Z E* P
@U)@)�PZ
@�@�@�T@�P � �
 �
jYA�V $�E %�djUe�V��j� Z��V��Z��j��Z� jU� ZP �P�P i)@�
P��� ZP�P�
P�@�@F
X@�X@U
X@Q* �Z ��` ��`����Rhj�U  �F � ��J�����V�� ��V �� e�V i� %�@%j )`��DU�PQ  T V T h  h  `  �U   f  h  �Z   �               j� ��*�����Z��Ui�UVe�DEU� EU AE     @ Y AjUU�j�U ��   � ��� ����������U��eQ�FUQ�UQVE@ Q      P   P T�UT�Yi���Z �@U@UP
Q � �  �  @�  D)  T	 D� E�  V*  �  *           ��p� �0�2�����0i�0��1 .��p��`�)��ɤ���)������)��	Ɍ��	�)��	���	`��U�I�Q�q�M���I�q�E�)�� ?� ��)�� � �� �� ����� � �) � ��)������� ��`�q� ���H����� ���H� �x�r��q��|`����-�#�&�(��7�$�F�%�U�&`���` 	R�%H�)N�(G�7�      �  @� @     @  R %H )N (G 7� �& �m ���� �$�%�&��� �>��H�)�� �� �� \⥔�� �� ���� �񩉍& `���&   ��-�� �񩩍& `� �����������-�5⅐�:⅑����D� �L��T���00�� ��Щ �ҩ%�ԩ��ө%�թ �ׅօم����� ������?⅞�`BLT<(@d�����yX6(6WyH&&Gixi  0@P`p� ��q����?�I���!�"��� ���\������	 @��2�
�3�� � � � ������ �� � �� ���  � `� �� ����`� ��������� � � � � ��`��� �2�@�3�/� �2�� .����`��5 ��5�5� ��� �5� �4��4������z�{�|`��0 ����)���� ��3��2���� ��2 .����� \����`���y��2��� � �^�� � ��`�3�


����� ���2� .�����`�`�`   U    &  *   �)�2���� +�������@� ��������)�����)��`)*** """   � � �
����� ��`��`������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������0�p����b����������z�����&�B�F�:������������������������J�f�j�^��������������������>�>�>�>�>�>�>�>�>�>�>��6�Z�~��< <�<�[��[��[��k}鬾:���<?�<��<�<<<     � 8_�<ܦVp�i�j�5�ZY5�YU6�eU�\UY5|V�5\�����_�0 ��   �  �? ����j���f:lf�9�UU�k�Z髩e�kiU�jU�kj�鬪�:���:p���g� �?      �   �  �= �e� p�f���lVf���=lee�Y��f����  �>  �  �  �
X)h&�)�
<�<70�7���P��P��VU��ZU7L��5L��1�4��?\W�5���:�_�:�: � ���:�Z���k�[@�P:[�>k�;����?�?<���óAάA:\}5����\}5�A:�A����?<� < ���A�A:\}5����\}5�A:�A�� < � �����A�����A��A���;�A���U �  <  < ���<�<�<�<�(�(���} �  < �<?��� � ��?��� � �</��3�0<���� ?��(��<�\�5p���?����? � ��Z � ��0�?��;�������{��w��7��7<�� 7� ��0�?��;�����;�������;p���       � ��8<,<�<<����� �?���<��<7p�O��<<���[���������������S��CU����<<<�3����Ǔ�Ɠ�Ɠ�Ɠ�Ɯ�6��:�<�@�+��0�0�0�p�p�p������<C� ��?<�� ���� 7���F��F����U3���� �?<�� ?��Ɠ�Ɠ�Ɠ�Ɠ�Ɠ�Ɠ�Ɠ�Ɠ��� ;0  �  ��������� � � � � �  0 <�C�LGk0��|����ڧG�=Cz4��0���?<�?<0����Cz4�=�G����|����Gk0�<�          ��W�a�����W �      ���V��5���� � �W�^E�\$6����<�3�������������i��i��?��:p�����0��(7��Ǔ�Ɠ�Ɠ�Ɠ�Ɠ�Ɠ�Ɯ�6����0������������������ �  <  <  �  � �������� �  �  <  <     �� ���?��?��������?��?� � �      �����}�}����� �      � ���:l}9��?������?l}9��:� �     � ���:��?������?��:� �    ��*ZU�����U�vA�v �v �vA��U����ZU���*��������A3�A;pp<�4�40��� <         �����VU��������� <       ?<����S��W��W��י�צ�����;,�8,�8 < 3\w|wp~����|U= ������/? �  �  � ��?�u��|U= ������/? �  t  � � � t  } ��?���kU�lA9�A �   @ @ @    } <}<���kU�lA9�A �  < ��L�1S�ū���A;�A?��ꗾ֓���A? �     < ��0}p���3��30�p~�� <     � �A?W<�������<��������U��U?(�( � �U?WU����7<�7<����7<����WU��U?(�(����>,P:�O��O��O���������, 8��>������>,T8���������3�����,T8��>������>, 8������������������, 8��>��eY�����zL9L9L9�ppp�ppp����������������������������& ���z�{�|� � � �* �}�~�� �����[�© �Åąȅũ�& �������� [� ������������i<����`�����`�����>�]�:��8�� ���i0�ƥ�i �Ǧ������Ƒʈ��ƅ�i0�ƥǅ�i ���������  ����a�.�]�*�D ������ȑʈ��� �ʥ�i0�ʥ�i �������� ���_��a�Ș ,���a�����`��`�����`���K�]�G��8�� ���i�ʥ�i �˥�i0�ƥ�i �Ǧ������Ƒʈ��ƅ�i0�ƥǅ�i ��������� ����a�0�]�,�D ���ȱʈ����'��� �ʥ�i0�ʥ�i ����ߩ�¥��a�����`��`



}I�ƽJ�i �ǊJ��� ��M�eʅʥ�i �ˠ�Ƒʈ�`� � �ʩ@�˥ɑ���������`H)����hJJJJ��
e�i@}��` 0`��� P���@p��      

�� �A� � �����`� �/ �O�O� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                  㩠�  � �� � � �� ���� ����& � �-��  ���� ���?�	�& `� �@�A�B�C�D�E�F�G�k���<���I�m�l��H��=`� �&  �� ��?��>�����!�"�I�m��l����ɍ& ` �����������z� ������`��
��5􅰹6�`�z`ƺ������Ƶ`������ �� ����ȱ��������U���ȱ�����������z� � � ������ȥ���ƶ����L2�����ȱ�����L2���ȱ���L2�HJJJ����hL2�}ȱ�� � �� h)� � �� ��� � ���� ��� � �� �L�n��0e͐ͅ�Υ���� ��`eͅͰ�Υ�0�͍ �΍ `�{08

����{��� � �����)� � ����� � ��� � �}�}�v���e)x�aJJ�����	���R��N��0.��8����΁� ������� � ��� � L��m����������թ ���}�� � � �|0

����|���( ���) �~���* �~�	�~�� �* `l�o�xo?9d*o/z Y � �� B B /B ?B OB _B oB B �B �B O����������m�5�K�]�W���U�U�"<  < < !�  � � !�"�!�"�"<"�#X  "<  < < !�  � � !�"�!�"�B<@ ! 	    � � � � � @ � @  T �0 @ 	@ @ @ !T �T � !@ T} � !�`   ��� 	� � ���� < �<  � 	� � ���� �T  � � � ����  }  � �� ��  �� � ��<  � � ��� �� ���  �� ��  � �� ��@ � � � ����  � � � �� ���p   ��� ��  � < <�  < � ��  � ����X�� � ��  � < <�  < � ��  � ������� �T  � } }<  } @ @�  @ T@T}�}T � ��  � 	 	 �� � � �� ��� �`   ��T T �T �@ @ �@ �  FT T �T ���} �  �  < < �} <�����0 � � <� <} } <} <T T �T �} } }  � � �� �  � @ @ �� �����0   ����� � �<�� �� � � � �<< �< X � � �<�� �� � � �<<�� <�  ��  X  �0   ��� �� � � � ���� �� � @ @ @h@ @h h � �@T  @0   ����X X ( ( X X � � X X ( (�  HX X � <  �  <� � � � � � � � � @ @ T T  
 
 < 
� 
�   ����  @ h �@h�h�   @ h �@h�!h  h   @h�@h�h� � � � 	@ @h�<�"  !!!@!h�@h�h� !!!@!h�@h�!h  !h!!@h�@h�h�A "�!�!�!@h�<"�B   s�s�<�<�}T 	   0	@ @T}T 
< < 	@ @T}T 	� �@�@� � @T� 	� �@�@� � � ���) T@T}T@ � .T0� <�<�}T  @ @T}I� ;�;�.}.�.�`� Q�Q� �!!T!�� c�c�!�!}!!}� T �0 !�!T �.T} � 0 !�!}!!}� T �0 !�!T � �  \� �  !}  � � 0 �}�} } �T�T�0 �T�T� .T}�}�0 �}�} � �����T0 ����T � �  �.T.  } h.T.0   ]�]�1�
< 2< 1�}1T !@ @!T!}A@ 1�
< 2< 1�}1T 1@ @)T1}�� ����a@`�1�@aTa}a@1T@T}a�a�1����1�T}a�A@!T1�@T�a}A*<aTa1@T}Ta�aTa1@��a@� �@�!@��Ta�A}!T1@T!}a�@ !�  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xة �& �� ���  �   � O� f̥)��� �� �-�>��������-��: d� �� �ťk����)@��津���� �� ��L<� ��  ��lЪ�m��Le����&  ����  �� � ������ ��ɍ&   �L��H�H�H� � ��  
� �?�?��;��7�� � f̥)��'� ���� ��L����)� f� x� �ͩ��?���h�h�h(@�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � �