  �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                  �?���?          ���      ���;�;��  �������������   �   �   ���?���������«���[i僾[U微ז׺^7�ܵ�7�ܺ�7�ܾ��i���Vi���VU��W�Հ[U��U����π��ހ����������JU���RU��   ����������� 0� 0�< <���>��U=�U����������������p��-�x��-�x���p���i_��UUU����W��VU���ZU��«��������� ���
���j�UB���U��   �   �����������   ����0����:������������������֪���ު�������2<�<��2댎�ʂ��r*è�©<j���ڀ����y�m���U[�r��Z������pU��\U5��_U��   ������� �<�<���?��[:隦k�i��UU�kf��k�f�kV��V���Ye:�Ye�V�:oV��k�f�kf��UU�ji�隦k��[:���?<�<� �      �  �<�<�:;�k���j�Z�>�f�:kj��[V��kYe�kYe�[V��kj��f�:�Z�>��j�k�쬺;<�<  �  �                    0�<�<��;����ii�V�s�ͬP:�P:s���V��ii�����;<�<0�                �������  �  �  �  �  �  �  �  �  �  �  �  �  �  �?  �?  �?  �?  �?  �?  �  �  �                                  ���?   �����   �����   �����
  �����
  ������  \UUU��  \UUU��  �����  �����>  �����  �����                                 ���������������������������������       ��������������������������      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��������������������������������       �������*�������*�������+�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +���      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      �������������������������       ��������������������������������      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�������+�������*�������*�       �����������������������������������������������������������������        ������������������������                                                                                                ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��                                                                                                      ������������������������        ��������������������������������      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�    �� ��* ��
 �z �v hv hV �� �]5 \��?�uU��wU�\�?\��|�� �5 |�5 ��? \}= ��? �~5 ��� ��� �
 ��� �j* �� ��5 ��5 �Y5 �V? �w� p��?�ו���U�p��?|��\�? _W� �U� �U� ��?  W  W  W  �  �?      �?  �� �V��0���Z��Z� �� ����]�����Z�:��v5�W������� �����_=p�W=��W�*�>���:  �?     �?  �� �V��0���Z��Z� �� ����]�:��5�Z�?����W���� ���|��|�Zp�Z)���*���?��       �� ��* ��* ��* p�* p�) p�) �_* \u���5WU]�WU�����5��W5 �W= \� \_= ��? |}5 ��? \� _������ ��  ��
 ��
 p�
 \�
 \g
 \e
 ��
 W���_V�7_U�?�w�ww= ��5 W�� WU� WU� �� p�  ��  ��  �?  ��      �*  �� ����6��r��r��J� �� ����.8����_�:��5p��5p��?��� �*���W=p�W=��WX)�?��_5  �?     �*  �� ����6��r��r��J� �� ����,8����^����>�5���5 ��?�|��|�Zpժ*��h%\��?��        �� �� p� �:> ��; �~: ���?�����nU����?�����6 ��6 ��6 ��6 ��: ��? �� �: ��� �����   �� �� p� �:> ��; �~: ���?�����nU����?�����6 ��6 ��6 ��6 ��: ��? �� ��> �: ��: �Z� �_�  0  0  �  �:  �� ̫���k��k?��������뫪��������?���;���?���:������������>��:�>�꼾�����  0  �  �:  �� ̫���k��k?��������뫪��������?���;���?���:������������:����:��:��?�: ���  0  �� ��? 0�= ��> ��? ������گ���_�����z����� ��� ��> �� ��: ��> ��? �� �� �� ��? �� ��  0   0  �� ��? 0�= ��> ��? ������گ���_o����z����� ��� ��> �� ��: ��> ��? �� �� ��>�:���? 0  0  �  \5  �� ������3���3�ʣ�������������o���_��[���Z��j������������������.���?���  0  �  \5  �� ������3���3�ʣ�����G��������o���_��[���Z��j�����?��������?���>������> ��� ��  ��<�����p�� ��� �� �� �������>�Vo5�R�?�Zn5��?��o5���? �+ �� ��  �: ����Ϊ���?     ��  ��<�����p�� ��� �� �� �������>�Vo5�R�?�Zn5��?��5��?��+ ����� ����>��� �  l9 <k�<�[�7p����j�W�|��=��������������������纮�纮����밿�>���p�=p�p�>���?���  �  l9 <k�<�k�7p����j�W�|��=����������������ۛ���ۺ��뺮����;����|�p��:��?�; ��?     � ��: ���<���7 ��������  �� �������?\��7���7\��;���;\��?�������  g��j�����?� � ��: ���<���7 ��������  �� �������?\��7���7\��;���;\��?������ ���  ��  �� ������� �  �: <��<���30�������z|�n=���������槮�槮�����箺������;����|�p��:��?�; ��? �  �: <��<���30�������{|�o=�������ڛ�ڛ��ڛ��ڛ���뮺������簫�>���p�=p�p�>���?���   �?  05  O= �P ��P=0�Wp}�:���:���.+��k^�:o�W5L���|���Z�����;��� � �� ܑ �� ��> ��?      �?  = �P ��P=0�Wp}�:���:���.+��k^�:o�W5L���|���Z�����;���? �� �� ߛ����������?  �7  �7�?�ܫ�7ܪ�7pZ�p���Ye����l\e�lne�ln��ln��ln��l����������6��6p�6�����=��;����*   �7  �7�?�ܫ�7ܪ�7pZ�p���Ye�����l\e�lne�ln��ln��ln��|������.���6p�p�=p����5|*�6���� ����  \  |�  � �_� |�p�_�^}������֪�������\շ���1��=�ϥ���?����� ��? �F7 ��: ��� ���     �  |�  � �_� |�p�_�^}������֪�������\շ���1��=�ϥ>���?������ ��? ��� ����:��?�  �3�?�3W���u]3�}}3��W�UU�����|j�=\��5\��?\��?\^�7\��5|��?�֫�����k\�k���K��6 �?  �3�?�3W���u]3�}}3��W�UU � ���|��=\�5\��5\��?\��7\��5���=�j�?�����k>���5��?��������+      �  ��  [z [� �� �:  �� ���p��z��_����z����皪ܪ����� �� મ�������:�:�:�:�?�? �  ��  [z [� �� �>  �� ���p��z��_����z����皪ܪ����� �:  �:  ��  ��  k�  ��  �� �� �  �:  ��  ��  |=  � ������?������뛫�����������������v:��o:�=l:�=l:�=l:��l:����  �� �  �:  ��  ��  |=  � ������?���뛻�����������������W����z:��o:�9�:�9l:�9l:�9��������   �  �� ��� ��� ���  �>  �� ������o����������������f�7������ �:  ��  k�  ��  ��  �� ��� ��      �  �� ��� ��� ���  �>  �� ������o����������������f�7������ �� ����.���:���:�ڳ:���? �  �:  ��  ;�  �:  � ������?�i���Y��۪���J����������V��l�v:l�o:l9l:l9l:l9l:��l:����  �� �  �:  ��  ;�  �:  � ������?����U��۪���
����������V����v9��o9�9l9�9l9�9l9�9o�������       � ����֫�֫�~���� ����~���֫������~��ֿ�V� ��� ��� ��� �������k��j����3�{������ � ����֫�֫�~���� ����~���֫������~��ֿ�V� ��� ��� ��� ��� ��� �k��k����#�{�>�ڪ��� �   �  �> �����?�k�?�n�?���?�Z�竪�����﫦������������������l��>������?��:����������  �   �  �> ���?����k���n�����?�Z�竪�����竦�������������������p��>������=��:������� ��? � ���?p��p������ ������?���?�����;��+���; ��; ��? �� �� �� �����
���Ⱥ�.���:�:����     � ���?p��p������ ������?���?�����;��+���; �� ��? �� �����>�������~����/��������    � �; �o�ޞKޞϯ����������o�����z�������v������������ϼ�~9���p�?�:�>�:��?o7 ��?    � �; �o�[ޞ[ޞ�����������o�����z�������v������������ϼ�������p��:�>�:�>�>�?��*      ��  W]��W|UU�Uj�_j�]� �u� ��������:��W������:����Z��� ��� ����=���h�������? ��  W]��W|UU�Uj�_j�]� �u� ��������:��W������:��������� ��? ��6 ��6 ����ZU������  �  �  �? ������:���:���:���:�������������������?���:�����6���7����:�7�>��>�:���?�  �  �  �? ������6���6���6��ڶ�����������������6���?���:�����6���7�������:�>�?���?�� T�? �? �u� ����UU=��U����� �u� j]��Z��������_�W�����������W�� ׯ� ��? �� ������U���� ��     �? �u� ����UU=��U����� �u� j]��Z��������_�W�����������W�? W� ��@����|�)�s*�?��� �  p50|���Z?�}�=l�;l���l���������_�o^׶����_W6��}>���w}�w}:�v}:�v}
�������:�?�: �� �  p50|���Z?�}�=l믿l���l���l�����_��_׶k�>[^W6��}6���?��u��u��u:��u:����o���:���?��
                                  V      QE                � R   � � @                  �`      � P P  (                                                                       �    � Z �  �*XU   ��V   �jUE�   �jU�   ��UUU�  ���   �jUU  ��e�V	  (���U�   �*��                                                                   ���   �jU�  � P�  �UP�
  �VQ��*  ��B��
  H�F�*  
��V�  
X穪  heU<�+  �eU�
   ����                                                                      �     �   ���3   < <��   ���;  / ���  �����3  ���ʮ>  ��� �;    ���;     ��     ��                                                                   �      @0     0<�  �/��=  _�<|��  ������  wU�U�  ��WU��  {�j�  ������  �D   � �                                                                   �@            @             	     @  �  �       @                     @   �   @                                                                     ��   ?  _U  ���WU  {U�UU=  ���Wf5  {W�}U?  {W���5  {_UjU:  �i��6  \�UUU�  \�����  \�UUU�  p�UUU�  p���  ��eff�  ������                                          ?�?��   �W���  ��Z��:  �[�= ;  {_�? ?  {����5  {_UjU:  �i��6  \�UUU�  \�����  \�UUU�  p�UUU�  p���  ��eff�  ������     ��   ?  _U  ���WU  {U�UU=  ���Wf5  {W�}U?  {W���5  {_UjU:  �i��6  \�UUU�  \�����  \�UUU�  p�UUU�  p���  ��eff�  ������                                          ?�?��   �W���  ��Z��:  �[�= ;  {_�? ?  {����5  {_UjU:  �i��6  \�UUU�  \�����  \�UUU�  p�UUU�  p���  ��eff�  ������                                   ���  �����:  �WUUU5  �w����  �W7  �  ��wUU�  ������  �����  ��z�m5  �׫�z5  �W��5  �wUUU7  �W�_�5  �:�;  ��?�?  �W��7  �UUUU5  ����6  _U}�]5  ��{��?         0���AUD�?0�                                                  @  @   @A         �YB              @j     A   P  
 �    �
 
  �*��  @ (  $  @  $   @
  �      P*    �$@                                            *      �@      � P   T( @  @�J         �         T@      $ P @  ��      (   (
 �    � �      ��*    @	   T T      	     U
  �    � �   ��*       (    �  �   $   P @  @U ��       H  @ @          @                                  �   *   �   B     �@  �  T   �
          �  � @  �  � P   *      @�ZA             @ @   @ @ @    T       D                                                                    ������ �갪�� ������ _�z��W� g�U�U� \UUU�VU lUUUiUU ��UUVUU ��UeUUU ��ZUUU� WVUUUU� �������                                                                 �     ��     ���  � �U� � �U�� �; UUի�W; UUU��U� �ZU�zU� YYY�_U� ��jVUU� ��UUUU� ������?                                   �vu    �vu    �vu    �vu    ��    �6p    ��    ��u    ��u    ��u    ��u    ��    �vu    �vu    �vu    �vu    �vu    ��    �6p    ��                                     ��     �_��    pUU�    p���    ����   �U�^5   ���U5   ���:   ���Y=  ��~�?  �:�~�  |%���  \9���  \��U�  l�oW�  ��UU�  �^���  �^���  ����U  ���WU  ���UU  ���i�5  ���?  �m���  ������  ������  �ꪞ��  ������  ������  ������   �����     ��?                                                                     ��     �UU
   *hUU%  ��ZQ%  jU@%  V�@U%  V� T	  UQU%  FU U�  FUU�  UP�  VEUA�  XQUU&  ZUUU*  TUUU	  VPYQA)  AjU�  FQj�V�  Uj��  �j�V�  V���U�  XU�j$  XU�ZU%  h��ZU%  �
�jU%    ���
    �*�     �*      �*     ���     ���*   P����                                 ��������UUUUUUUUUUUUUUUU��UU�UfU���UWUU��{�U]U���~�UyU���{�UyU� �~�UyU� �_�UyU� �^�UyU �_�U��� �^�UyU� �_�U���@�_�UyU�@W]�UyU@W_�Uy��@W]�Uy��@�_�Uy��@���U������   ��UUU ��UUU����UUUU��zU�UU��ZuU5����VuU�?��p�w 0S�~U1S#��^U1Sc�]_�:Sc��W�? ��TU 0����TUU1�� �TUU1��b�TU�:�kb�T��?����T� 0�k��T�U1��"�?U1�kb��5���   ��UU� �UUUUU���UUUVU���UUU\U]�WUU�U]�n���W�����^��T �^�TLU�uW�TLU<�W�T���U�� ���U��� UU�LUUUW��LU�_W�鬪�~����� ����  ����LU \�W��LU��������UUUUUUU�UUUUUUU�UU�U�UU�UUU�UW���UuU^���sUmUz�� �UmUz��U�UmUz��U�UmUz���UmUz�?��nUz� rUmUz�U�nUz�U�UmUz����UmUzu���_mUz�� �mUzu�U�mUz��U��U�?�@� �U �@ר�U��+@���U��@W_�Uy��@W]��y��@�]�W{��@W]��}��@�]�W{p@W]�U}�p@W_}Uup@WW��_��@WWUUU�@�WUUU��@�WUUU��@�WUUU��@�[UUU50@�_UUU�:@�W��_��@�WMUmU�@�UMUmU��:��b�n�  諢�U��૪�U��� p�^�����ժW��UUկ�_�����mx=p/>��m�s-���m��/�z�m��/�^�m��/^WUo���.^UUl���,�_�l���,���l���,�
l���,  n���,�
�o���,���n���,^�_�W�W�ꬪUU����  UU^�����U�_ પ�W�������WUU�WU�������Uw���-9Uw��x�/9U����/9�����/9UUյ�/9UUU��>/9�_��8�+9����8�/9 �*�8+9   �8�/9�
��8�+9����8W+9U��8W/9�� pU � �zU�*����U�?ת�mUz�տ�mzu�����zu�_}~u�yp��zu�y}U{u�yp]U}��y����ypUUU����UUU��9�UUU��9�zUUU��9\UjU��9�^��U���_%V���_U%V��^U%VU�@�uM�mU�@�UM�mU�@puM�mU�@pUMjmU�@��MUm��@��NUm��@\�N�m^]@\�O��_�@|UM��W�@{UMj]UU@{UMU]UU@sUMU]UU@��NU]��@�� \��@����z @��[U�  @UUkU}UU   kU     kU     ��  o8��+^UUl���/^UUl8���_UUl��կ^U|���� �s������o�UU���_xUU�WUUuxUUUUU�m�UUUU���UUUUՠ��U��Uը�������?�� �����    ���?      UUUUUUUU                        UUU��W/�UUU��W+�UUU�?W/� PU��W+y�
 �?�+}���:��/�U����U/yUUU�_U-��_UUUU-] �WUUU/y�
WUUU��*WU�Z�z�*�������*�� ����   �:      �UUUUUUUU                        �_U��W]?zU��UU_wUUUU]UwUUUUUU�������������?UuUUUUU5�UUUUU5UUUUUUU=UUUUUUU�UUUUUUU�UUUUUUU�������Z�������[�      [�      [�UUUUUU[�      [�      [�      ��o8��+^YUl���/_�Ul���U�U\X��_U5|���W������U��?�UU��UU7�U��W��u���_U��e _��WU��}UU�W��*ܪ* W����0�Vg��� ��U ��  �W� �  ��?UUUUUUU                        UP��U/�@w��W+���U�3W�u��Wy�~E�?h(u��T�X�u�Q�}!u_U�E�_ �UU�WUU,_U�A�_�{o�UuU��ZU�ګBUU��ð�*� �����  + ?     < UUUUUUUU                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                  �?���?          ���      ���;�;��  �������������   �   �   ���?���������«���[i僾[U微ז׺^7�ܵ�7�ܺ�7�ܾ��i���Vi���VU��W�Հ[U��U����π��ހ����������JU���RU��   ����������� 0� 0�< <���>��U=�U����������������p��-�x��-�x���p���i_��UUU����W��VU���ZU��«��������� ���
���j�UB���U��   �   �����������   ����0����:������������������֪���ު�������2<�<��2댎�ʂ��r*è�©<j���ڀ����y�m���U[�r��Z������pU��\U5��_U��   ������� �<�<���?��[:隦k�i��UU�kf��k�f�kV��V���Ye:�Ye�V�:oV��k�f�kf��UU�ji�隦k��[:���?<�<� �      �  �<�<�:;�k���j�Z�>�f�:kj��[V��kYe�kYe�[V��kj��f�:�Z�>��j�k�쬺;<�<  �  �                    0�<�<��;����ii�V�s�ͬP:�P:s���V��ii�����;<�<0�                �������  �  �  �  �  �  �  �  �  �  �  �  �  �  �?  �?  �?  �?  �?  �?  �  �  �                                  ���?   �����   �����   �����
  �����
  ������  \UUU��  \UUU��  �����  �����>  �����  �����                                 ���������������������������������       ��������������������������      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��������������������������������       �������*�������*�������+�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +���      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      �������������������������       ��������������������������������      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�������+�������*�������*�       �����������������������������������������������������������������        ������������������������                                                                                                ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��                                                                                                      ������������������������        ��������������������������������      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�      +�    �� ��* ��
 �z �v hv hV �� �]5 \��?�uU��wU�\�?\��|�� �5 |�5 ��? \}= ��? �~5 ��� ��� �
 ��� �j* �� ��5 ��5 �Y5 �V? �w� p��?�ו���U�p��?|��\�? _W� �U� �U� ��?  W  W  W  �  �?      �?  �� �V��0���Z��Z� �� ����]�����Z�:��v5�W������� �����_=p�W=��W�*�>���:  �?     �?  �� �V��0���Z��Z� �� ����]�:��5�Z�?����W���� ���|��|�Zp�Z)���*���?��       �� ��* ��* ��* p�* p�) p�) �_* \u���5WU]�WU�����5��W5 �W= \� \_= ��? |}5 ��? \� _������ ��  ��
 ��
 p�
 \�
 \g
 \e
 ��
 W���_V�7_U�?�w�ww= ��5 W�� WU� WU� �� p�  ��  ��  �?  ��      �*  �� ����6��r��r��J� �� ����.8����_�:��5p��5p��?��� �*���W=p�W=��WX)�?��_5  �?     �*  �� ����6��r��r��J� �� ����,8����^����>�5���5 ��?�|��|�Zpժ*��h%\��?��        �� �� p� �:> ��; �~: ���?�����nU����?�����6 ��6 ��6 ��6 ��: ��? �� �: ��� �����   �� �� p� �:> ��; �~: ���?�����nU����?�����6 ��6 ��6 ��6 ��: ��? �� ��> �: ��: �Z� �_�  0  0  �  �:  �� ̫���k��k?��������뫪��������?���;���?���:������������>��:�>�꼾�����  0  �  �:  �� ̫���k��k?��������뫪��������?���;���?���:������������:����:��:��?�: ���  0  �� ��? 0�= ��> ��? ������گ���_�����z����� ��� ��> �� ��: ��> ��? �� �� �� ��? �� ��  0   0  �� ��? 0�= ��> ��? ������گ���_o����z����� ��� ��> �� ��: ��> ��? �� �� ��>�:���? 0  0  �  \5  �� ������3���3�ʣ�������������o���_��[���Z��j������������������.���?���  0  �  \5  �� ������3���3�ʣ�����G��������o���_��[���Z��j�����?��������?���>������> ��� ��  ��<�����p�� ��� �� �� �������>�Vo5�R�?�Zn5��?��o5���? �+ �� ��  �: ����Ϊ���?     ��  ��<�����p�� ��� �� �� �������>�Vo5�R�?�Zn5��?��5��?��+ ����� ����>��� �  l9 <k�<�[�7p����j�W�|��=��������������������纮�纮����밿�>���p�=p�p�>���?���  �  l9 <k�<�k�7p����j�W�|��=����������������ۛ���ۺ��뺮����;����|�p��:��?�; ��?     � ��: ���<���7 ��������  �� �������?\��7���7\��;���;\��?�������  g��j�����?� � ��: ���<���7 ��������  �� �������?\��7���7\��;���;\��?������ ���  ��  �� ������� �  �: <��<���30�������z|�n=���������槮�槮�����箺������;����|�p��:��?�; ��? �  �: <��<���30�������{|�o=�������ڛ�ڛ��ڛ��ڛ���뮺������簫�>���p�=p�p�>���?���     �  �� ��: ��� ��� ��� ��� ��� �� �;� ������s�p����� �V9 ��9 �_? �+5 ��4 ����ͪ��� �  �� ��: ��� ��� ��� ��� ��� �� �;� �����5�s�5p����� �V9 ��9 �^; �^; �_?  _  _? ��� ��� � ����_=���l�l�~l_}l�����4�/�N_}������z��z�/���p�vp�~��� ��� �� �:��?� ��?� ����_=���l�l�~l_}l�����4�-N_}������z��z�����+p�vp�~��� ��� ����9��:���*   � � �z �> �z� ��� ��� ��� 0�� �������\��6\k�?�v �� l� l� � � �� ��  ��  �� ��      � � �z �> �z� ��� ��� ��� 0�� �������p��6pk�?��v �� l� l� �� \� ����:��s: ��� ?0�3�}�=���9�]�9���9�]�9�=�9�����^U�[^U�[��������������Z?�����z �^ WW �^�׬>���?��� � ?0�3�}�=���9�]�9���9�]�9�=�9�����WU�^U�[���[��������?��Z�����z �^ WW��^��\���: ��?     �  �  �? <�� ,� ��� ��� ��: �� �� ���������?�����[�?�o� ��  ��  �:  �? ��� ���3�� �  �  �? <�� ,� ��� ��� ��: �� �� ������?�����k�?�� ��� ���  �:  �:  �?  l  l  l  �?  <� � �<�7�۬�l�������� ��������?l���ln����������������:���:���?��������?��  <� � �<�7�۬�l������� ���������:����n����ꬮ�����?�:�:���:���?��9���9  �� �?  ��  ��  ��< ��8 ��: ��: ��: ��: ��:��:���?���
�w�
 �� �� �� ��  ��  ��  �9  �9  �9  ��      �?  ��  ��  ��< ��8 ��: ��: ��: ��: ��:��:�V�?������
�w� _� �� ��  ��  ��  �����?���< �; ��; �?<�>��^;����:�[� �����������;��;���;��;�w?������������l�l��?� ���< �; ��; ��?<�>��^;���:�[� ������_?��;���;���;���;���?��������������l�l����   �  �:  � �u ��������� �Z��Zk�Z�>�Z�>�Z��۪U���������V���� ���  ��  ��  �� �� �     �  �:  � �u �� ������ �Z��Zk�Z�>�Z�>�Z��۪U������������zp�o|��=�Ϋ��:�����? �  �;  ��  ��  ��  �� ������ﻮ^������z��^���׫�������������k��j��jp?�:��?� �� �  �;  ��  ��  ��  �� �?����ﻮ^������z��^��׫�������������o>��k:Щo?����?�?�:�?��
  �  �: �k� �]� �� �;���? �����������������wU�翪�?��_��� �� _: _� o: 0k� �� ��      �  �: �k� �]� �� �� ��?? ������������������wU�翪�?��_�����np��|�=_��6�:�:�� �  l9  ��  ��  ��  k� �������[��n������������﷮����������p��p��=Щ�=Щ����t��9t��?��
  �  l9  ��  ��  ��  k� �������[��n����������������޷������p�|�j|�jp�jp:o|;��?� ��    �� �U= pZ� lou������7���?�_m7�j�5���= �w �� ��  �� �� �� ��
��g�������fU�&�9�?�?�� �U= pZ� lou������7���?��m7�j�5���= �w �� �� �����������
����>�_���  ����*���       �  p7  \� ����\��ְ�:�����W � ��  ��?��[>��[� �k> �����0�kp�o���:��?� ��?       �  p7  \� ����\��ְ�:�����W � ��  ��?��[���[>��k> �� ������2 ��7�����?��*  �� |U W��]�9p_^�ܟW���y�\��|ުp�� ��� ��. ��> ����j�Vo0Z��~��� ����� ������     �� |U W��]�9p_^�ܟW���y�\ߩ|ުp�� ���  �. ��> �Z� �� ��� �٧@����pU�lj����? �   �   �  \  W5 �_��W5�}_�w��U���� W��^������p�� \�� \�k\�k09k��� �9[��� �� �   �   �  \  W5 �_��W5�}_�w��U���� ���߯�W�� ߥ� ���p�jp�k\�kp9kp�jp9[�����                                  V      QE                � R   � � @                  �`      � P P  (                                                                       �    � Z �  �*XU   ��V   �jUE�   �jU�   ��UUU�  ���   �jUU  ��e�V	  (���U�   �*��                                                                   ���   �jU�  � P�  �UP�
  �VQ��*  ��B��
  H�F�*  
��V�  
X穪  heU<�+  �eU�
   ����                                                                      �     �   ���3   < <��   ���;  / ���  �����3  ���ʮ>  ��� �;    ���;     ��     ��                                                                   �      @0     0<�  �/��=  _�<|��  ������  wU�U�  ��WU��  {�j�  ������  �D   � �                                                                   �@            @             	     @  �  �       @                     @   �   @                                                                                                    P      T�    @uU    PU�    T��:    U���  @U���  @ժ�*  PU��<  P����8  P�(�8  TU(��   T*��"  TU)��*  TU)��
  Pw���
  @U���   ���*    �?�
    ���    @UUU     U�    ���    ���     ��?      �?                                                                                   �*     ���
    ���*    ��*    z���   ���f�   j��  ���;�
  ��ⰰ*  (���:*  ���;��  ��l���  ��a���  �-h"��  ���>*  �����+  ��k��
   ��ʨ
   *���   ����    ��/(     �.      �      ��     ���<     ���     ��    ���    ���?     ��?     ���      �?                                 j�U��Z� ���jYj
 �U�VZi �Vi�je  �U���i  ZUVU�  �Z	@Y  Y� U� i� �  ���
   Y��  � U �j  $ * Z�eB     �     � �   ��                                  �U��Z�� ��jYj�� @�VZi�Y @i�je�V @���i�� @VU�ZZ� @�jY��V  Y�U��i X��UU� 
�
PU�� �A`��� �  P��     @��  ��i �  �	 @   ��% �                                                                )       Z      �Z     Y�	     i�     ��)     Y��Ai)  U��
�Z  j�Z�T  ��i��  �����)  ��f���  �Zje��
 UUVYY� YU��j� Ue�V���                                        �      P�      �V     ��i     PU�  � T��  �Yi���  �j�Z��  X�eV��  i����i ����i�Z �f���i� Xje��ZY TVYY�Vj T��j��f e�V����j�U��Z�����jYj���U�VZi�Y�Vi�je�V�U���i��ZUVU�ZZ��Z�jY��VY�Y�U��ii�Z��UU�����ZU��Y��Yi���U��j�Z��j�Z�eV����i����i�����i�Z��f���i��Zje��ZYUUVYY�VjYU��j��fUe�V����                                 <      ��      <���    ����      �   ����   < ����  �?   �  ������  �� ?�  �: 0;  �?3�?;   � ��   #��   � �®  ��<���  0�򫰮  0����  \ �+  _� �*  W�U��*  �Uպ
  �����
  �����  �Ϫ��  �����   ������  �����  030̿:  �30��:  <���  � �                                                                   � �    0?��    <���   ���   �:�>    �:��   �����   0���   0?+;   0��  ��*��    �����                                                                    
�
    ����   hU�U
  ��VVj%  ��iU��  `U��V�  �VUj@�  `T�  XAUQ�  VPUU"  VTQUU  UTUT	  VTUP	  �EUUQ)  `QUUE%  XUiUE%  XU�UU�  V��U�   �%���   &&��V  ���j   ���    �*      �%      �%      �*      �%      �%     ��*   �%H  � �%   P	�j�                                                                                                         �*     � ( *    U���   `U� �   JQD  @U @
  
U 
  
  
  ZP T  h PU)       (                                 �        �            PU     U      U        *      �*      �     ��      �*      )                                        P  �  T �  B @�  XP�  hA  T   h  U�  �UPU�  �RUU   �UU*   
  �
   �
��   ���
     ��     ��                                                                                       h@*     Xh      Y     �VU     �PU    jU    �(       *      `U      �U     �Z      �j                                      "  P  P( T U	
@ @UPPA� TA  T@  U  U PUUPUU UPUUPUUUUU          U     @U @U D@QDU  @U @Q U PeU   P�ZUP TT(U PU�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                  �?���?          ���    H�Z��	�	���������  ����8��������@ 4��|� "���ҩ"�����8������  ������	���@ 4�8�������	��8������ �����@ 4��N� "ဪ "� "��������	�  ��� �@ 4�i���  �����@ 4����	� ��� �@ 4�8���� �����@ 4��� "ဣ���� ��( 6�z�h`H�
�����轗���h` A� �� ���	��d�  ���L�����'
��㈅�㈅ʽ���轛��d1 4��� 6�ɩ�	�����%����^��<����轛��d1 4��� 6�թ��!�	������>����轛����1 4����	������� � �� �� � �� �����<L���@����轛��d1 4����  �� "��d0 ����  �� "�� �ީ�� �� �� � �� 6�`d A���
��݈��݈��
�	�����P8��d1 4� 6����=�̩��d��

i� #ީ��t�� #ީ����� #ީ�����i #ޠP���  �� "������L������ `d5d9d:��;`d6d7d8`�0�	���dd��0�� � ����
 6��d0 ��d��	�����T


�������� ��d���4���=�� �&�
��O���O���=
�������� �߅d1 4���Ƣ 6ဦ�< 6�` A��� ������ #ީ��2�� #ީ��F�� #ީ��Z�� #ީ��n��  #ީ�����! #ޢ�� ��  ���� "��` A�d����
�*����	 Y����2����@d1 4� "� �@ 4���Х�%�' Y����8i2��
����@ 4� "� �@ 4���ө	��� �) Y����2e������@ 4� "� �@ 4����ѩ���
�) Y����2e������@ 4� "� �@ 4����ѥ� �# Y����8i2����@ 4� "� �@ 4���ש
��� �$ Y����2������@ 4� "� �@ 4���� "� "�2�����	�/��
�����轉�	�)������B�e����i �� ����	0� "���e	��i ���ѥ5� �
��
������ �+i
�����轉�	�)���n�����	�����@ 4�i
�����轉�	�)���n�����	�����@ 4�`H�Z�
�����轉�	�)���� ��i��i �ʀ�z�h`���W���Ò�� �����o���O�ߜ��?������ߗ/�����/���o��ϝ��_�Ϙ?�����O������������9�H88HXXXH8(((#(#8#H#X#hhhhhXH8(#  	      	
   	  
	 	
		
	



QNUPR"X&S*O�P���.��� 


 
(
0
8
@
H
P
P2P2FPFZPZnPn�P��P��P��P��P���� �(�0�8�@�H�P�*(Z+F,Z8 2-02.@2+F,Z/@F0�
8�	0�8�
@�0�8�@�
H�	0�8�@�H�	8�@�@n�-H� 29�:�(�9 �: � �2�  *@n2 2(27827@2FF F(F0FZZ Z(Z0Z88F8@Fn n(n8n(�H��70�78�7@�7H�80�88�8@�8H� ��8��  *(�342(8@82@2 F(F Z(Z0F3HF4HZZ5n6� n8n@n8�@��0�� �� �5@�6@�8�H��5�6��  *(�% 020821@2(FHF#Z0Z$@Z0n1 n8n�$0�H��%(�0@�1H�$�(��#8��0�H��  ;(Z;(�;(�B(C(2!FAZ! nA �!�A�! �A �*�D8
E@
FH
GP
H8I@JHKPL82M@2NH2OP228F28Z28n28�28�28�2(F08�1@�2(n2(�2(�2(��   ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                �
  ���
�
�
����      8     888        �     ���  >>      �     ���  >>      �   �������>>      �   �������?>      �   �������?>      �   � ���  >      �   �� ���* >      �    ��� � >      �    ��� �>      �   ������>      �   ������>      �   ������>      �   � �
��  >      ��* ��
(������
      �   8� ��    8      �#  ����  >  �      �#  � 
�?  >  �    ���꣪�� �����>����    �������� �����?����    ������� �� ���?����                                                                                                                                                                          ����� *������
���
��* 
 
�� �#��8 �#8 �  8�� �#��8 �#8 �*�*8�⨊����( �#8���/��8
�������� �#8����8(� �����"�#8 ���8�� ���� *�#8 �  �8��� ����(�#8�
�  �8�� ����( �#8 8�  �8�
� ����� �#8�:�  �8�+� ������#8�?�  �8��� �����
�#8 ���8��� ����8+�#8 � �*8��� ����8,�*8�*�* 8�� � ��8  8 � 
 :�� � ��8 
 : પ��>�� ����:���>��������� ���?�������� �� �� �� �� ��0�� �� �� �� �� �� �� ����, ��������> :�*8��8?�8 �8�+8�8�?��? �?��;�:+ 8��>������> 8��8��8 �8�8��80 8��8�8 �8��8��8 8��>��    |  �  � �5 �5 p p�\s\s�p�=WU5�= p p p p �     �?  �� �?��� �   �   �   � < � ������� ��                  ?   ?   �  �� �� � �? �� ������� ��  ?<  ?           �? ��? ��� ��� ��� ������������< �0 �                    �?  ?  �  �?  ��  �  � �?  �   ?   �?  ��              �  �� �?����  ?�  ?<  <<  <�  <��?��� ��  �?                <   <�  ?�  ?� �  ?� �� �� �� ��  �   <                  �?  �� �     �� ��� �� �   <   �� ��  �?                  � �?� �� �� �� �� �� �� �� �? �� ��                          �=  �  ��  	�2� 
0  �@�� @p  �;  �         :  �*2�0�3�,�00� 3"����0(���
�8  +�30�  2<  �    ��������������������������������������������������������������������������j����j�����������������������꿪�������������V���j�j�e<�jU��jU���jUqժjUq]U�\sUU������������������*  ��   �����
���
������@U *�@U���CU �_U���l���o�>�o�>���������������������������������/ ���? ���? @����UU�{�T�_�C��ח^���^^�^9T������������������������������������������������������ꪪ���V���Z����U����������������������������Z������������������������U���jU���jU������j�U�j�VV�j�ZV��UiVU��ZU�5x�Up~�U\�_UU|��U�U�Z�_UZU��Wi`U�UXUU ^UU �~UU j�UU V�VU V�ZUVUj��o�>U?��>}���;�����������}���]���]����m��W�m��y�m�冀m�辶��讀����j�����m��_5��UW��W���W�J��S�JU�@�B�� �T�� ��� S��� ��������?�������������Z������������������������U����U��Z�U����U�V��UUU��TUU��@UU�� UU��U���@UU�?@UU�?@U�?@AU�VU�VUZU�VUZU�Z jUUZjEUe�UU�@U� U�V TUU @UU  EU  T  @          �VU��V��Հ���׀���@����@����@���P����P��~�PU�_�PU_�PU_�PU_UPU�_UPU�_UjU�WU_�������G����G]����W��W�����_U��WUU�_eQUyoYQU��VEU�WUEU�WU��_U��}UU��}U�������W����A����E����O������������[�����������U����W����_����������������������? @U�? PUU� PUU� PUU� TUU� TUU� TUU�  U� @U� @U� P� P�   �   �   ���      � � ���� ��U�����������ZU�����ZUU^�bUU^U
�U��������ç���ë�������*�����U���jU�WUjU�_Uj��_Uj�*XUj��aUi�V�Uj�U�UjZUViZUUXjUUXj�WY��jZ����U��_UU���U����_�U}կ�Uտ��U}կ�UQ���UQ���Vњ��V�j��V�j�������������W��k�~��j����j����ڿ�կ�������������_��������������߫���ת��������w����w����w������������������������������ ���? ���� ������������?����������������������������������������������������������������������u����u����u����u������_���_����_����_����_����jU�_��U�_��W���������������������������V����W���WU���WU�o�jU����V����j�������몪����������կ����V��������V��������������jU�����������U    U����U����U����Z�����UUUUU�����������������������������������������������������������������������������U������������������������������������������������������������������������������������պz��U���V����Z����jUU��jU���j����j����j����j����j����j����j����j�������     ���U��_U�����VU����������������������������������������������������������     ���������������������������������������������������������������������������     �WU�����U�����W�������������������W��V��������������������������������������������������������W���������������������������������������������������������������� ������W�jU���������  �?�����WU�������������?���  ���WU��������� ���?�����o�jUU    �������������𿫪VU������� �����=�<�󿦪jU��������?�����=�<�� ���U��������?� �����<ţ�說Z������������_�<�������UUUU���?������_�<�3����U����U��?�����?|�<�3��P������<��������U<�33S������? ���� ����T<�33�<� ���?��<S�������P������ ����<󣪌
(�B�*<3����������<򣪌�(��J( ?2���������<� ��(�J(������������<R����(�?J(����������������ʨ�?J(�����������<��ʨ�?J(��0���𨌌���<򣼎ʠE�O���������LL<�S H�S@E�O������OL@LL<�SUL�STUA�O�����OLALL<�SUL�SPU`�O��P�T��OULL<�SUL�S � ���� ��< <� ��������������������������     �                          �300 0���� �?��� �?����������000� ���0030 ����  � ���� 0�<03��0030 ����  � 0��� 003�3���?� �?��  <�?0���<�?003��� 0  ����  �� � ���� 000�0�00�  ����  � 0 ��� 000  �����? �?���  ��0�?��������� ���?� ��� ����?? <<<0<��� ���0� <<�� � <<<0<��� ���0�<<�� �� � < <<<0���  � � �<� �3 � < �<0�?��  �� ��� �? � �  < <0��� � � �<� ��  �  < �<<��� �� <� ���  � ��?�������??<� �����     ��      ���      ���>     ����     �����    ���j    �o
Wj    0�WU    0����    0��5�    �r5�    �Wr5�     W��i     W�Ui     _�UU    ���W�     <��_��    0�?� ���  �_ |�?���^ \U�uUUU^ �Uu��UUy�W�]W�DxpUU�U>pU�_UU���DxWU� �Uy�j�UU�Uy�`�UU�Uy�`�UU�Dx�`���?�Uy�`�]U90^�`����U^�jU���W�_WUZ�? �\W���0 � U��? � ������W�  |UUUUUU  pUUUUU�  �������  �������    W"6�   � W"6   �  \"6   ���_"��5  pUU��^U� |UU�U}UU |UU�V�UU \UUWW]WU= \U�U�W]U5 \U�U�UuU5 \UuU�U��� \Uu�pU ��SU]5pU�����5�U��0  p5 W �0��p5 � �0��p5  ���0  �     ���?           <         ; �      �: �      � �      ���      pU�7      \Ue5      ���      ���      �� �      ���      ]s	�     _%�     ]s%�?     �%\�    CU%�    �W�_U    \��~U   ����zw7  ���?j�W5  |]�����?  WgUU��_5 ������_5��zU����5���^Uտ�5��WUU�Z�5�W����5�� ����6��� ���W;��5 0��U7��5 0���?���5 0W�Uլ��5 0W��֬�z5 0W�����{� W�^�  ��U���  �U�����  0�UU�?   0�__���   �����_�   \��0�U�   W����UU  W�u���e �eU���YU �UVu��UU pUeu��UU �U���U�  \�W? ���  �j} �U�  �� ��  �*� � � �W��  �� �UY�  �V� pUV�  Wi� \�U�  W�u���:  WU�33ϵ  �W�=���  ��W5W��    ��?��*          ��        ��      �>      _U��     �pU��   �Ϭ���   p�����   pU����   �Ww���    �]���    �]��:    �߲�:�  ����0{  ���'��s  ��%��;�  ��	�W�  �U���>� zV��z�:� ~���� r5 ���Z r5 W��V r5 _UUU z5 |U�� z� ��  � z�0 TU�= zU��UUU�� ~U��U���� rU�ͪ���� rU��� 8� rU�PU=� zU= WUU?� zU5 W��3� zU5?���3� zU57� 3� �U57@�3� �U57W��<� �_5?��?�? ��? �?<  �3��� �  ��  �� �  � ������*   _���j   \U�U�0  \U�U   WU��U=   WU�U��  W��W�<  �U� �_�  wU5 <\� �_U� �| �UU��� pUUU�3? pUUU=�?3 ���U5�?3 0���?���� 0��030    ���03<     ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ��# ���ة��  ��� � � �
� �ߍ& ��" � t ����
 �� �� � �
���� ���� � �0�	 ��� �0  ��XL ��@H�Zx�' )�\�% � ��% �' � ��' �) � ��) �+ � ��+ ��
�$ �(��$ �+ �- � ��- �. � ��. �/ � ��/ ��# �� ��� � ��" �$ �% (z�hX@                          �� p� ���
 6�ߍ& �  Z��ߍ& �  A� e� e� ,̢F 6� �� 1� A� I� �� �ߩ ��  ��5 ��L�­  �� �����ߍ& ���R � �ߍ&  �ߩ ��  � �� l� ����ЊL� �����. P� �� �ŭ  ) ��  ����� &���� sߩ ��  �� &� �����T Y߭_ ��������� ���  �� ܀4 �έD � �E �  $���� ����� 4���� {ߩ ��  �� � 
����T b߭` ��������� ���  �� �܀4 VϭF � �G �  $����  ����� B���� �ߩ ��  �� 4� ����# kߜ  ��2 �0�3  �֩�  �2 ��3  �� �߮5 �< �9��4�P ��-�Q ��&� 6� ��  � ��ߍ&  h� A� 6��5 L'�LV��D �E �F �G ��( �* �  �� �����ߍ& L��R �& �ߩߍ& � � ��  � �� l� �����L�L� �����8 P� �� �ŭ � �L�í  ) ��  ����� &���� sߩ ��  �� &� ����� Y��# �# ���#  !� "� �� �� ����&�  ��2 �0�3  �֩�  �2 ��3  �� 9� k� ��L é�T �U ��D � �4 � � ����� �˩ �� ��  �� � � �(��  I՜H �I  ]� "�� � ��  Iթ�H �I  ]� "����� �� �  �� �����ߍ& L��R �# �ߩߍ& � ��  � �� l� �����L�L� �����	 P� �� �ƭ  ) ��  ����� &���� sߩ ��  �� &� �����# Y��# �# ���#  ��� � �-��  M� ����&�  ��2 � �3  �֩�  �2 ��3  �� �� k߭4 ���LM� ��ߍ&  ��L ��< � � �5 �E��S � �O ��& ��R �
�B ��C �I �H �N ��P �(�( �
�T ��D ���E �L �J ��Q ��( ��U �Q�F �J�G �M �K � �0��c ��� � � �� �x�� �Ȁ�`Hڭ  )�:�H � ��H � ������B �$�� �(��B �*� I�L�� ��L�� ��L�ƭ  )�<�H ����H � ������B ��� � ��B �� I�L�� ��L�� ��L�ƭ  )�9�H ����H � ������C �T�� �l��C �l�
 IʀM �ʀH �ɀC�  )�9�H ����H � ������C �4�� � ��C ��
 Iʀ �ʀ �ɀ I��h`Hڭ  )�&�H � ��H � ������B �*� I�L�� ��L�ǭ  )�(�H ����H � ������B �� I�L�� ��L�ǭ  )�&�H ����H � ������C �r� Iʀ5 �ɀ0�  )�&�H ����H � ������C �F� Iʀ �ɀ I��h`� �����c ������ ������ `ک� �� �H 
����mB m � ���mC m � � ��'�D � �D � �� �� � �  �����׀ %� �����
�= �*� ��`H� �� ��  �� �  nޢ �0��c ���� �
� �(�	 ��� �0  ��� �(� � #ީ� �4� �O i	 #ީ� �F� � #ީ� �T� �S  �� �d� � #ޜ �� � �6�� �b�  �ޮ  ���' nީ��  ��� �c�  ��� � ���� �����$ nީ��  ��� �c�  ��� ��� ������� �ީ��  �� � ���3L�ɭO ���O ��O �� �4� �O i	 #ޮO �J��&  Հ;�S ��4�R ��-��S 8��S حR i����R �� �T� �S  � ��L�ȩ� �
� �(�	 ��� �0  �� Iթ��� �� h`Hک�	 �� �B � �C � �  �ݭH 
����mB �B ���mC �C �I �B � �C � �  [݀�B � �C �  �O � �H � �I �  �˩�1  4��h`�B � �C � ��	 �� �  �� ��I �O � �H � �I �  �˩�1  4�`H�b  �˭B � �C � ��	 �� �  �ݭD � �E �  ������ �ݭF � �G �  ������ �ݭH 
�� }��� � }���  IխF � �G � �Q �X �K �V �M �W  ������ [ݜ1  4�D � �E � �P �X �J �V �L �W  ������ [ݜ1  4�B � �C � ��	 �� �  [� ��I �O � �H � �I �  �˩�1  4� ��h`Z�a � �0�S�a �c � �c � �c �� ����ޭb �a �� �����ϩ�	 �� � �7�� ȹ7� �ߍ ��1  4���z`Hڭ )� � 


� � 
m m 
���� �� �ߍ �h`H�Z� �x�	�i�� ��5 
��_�� �_�� � �x�� ������z�h`�� �P� � #�� � �5  �`Hڜ������� �̜������� �̩
� ��� � #ީ!� ��� � #� ��h`H�Z���&�����
��	L}ͭ�
��	L}ͭ����	��
L"ͭ�	��
�
�	�
�L��)� ���L[�����L[����0�L[͢����B��
 ���� �	JJ��
�
�	L%��
�	�
�L�ͭ)� ���L������L�����0�L�͢���	�B��
 ���� �JJ��
�
�	L��z�h`ڢx�� �� �� �� � �= � � � � �= ������� ������թ �`�� �� � � �� �0��`�c � � �c � � �c � ��� ��������� �7�� ȹ7� �ߍ ��	 ��  �������1  4� �c 耚`� m � �m 8� � � �7�
�3� � �+� m � �m 8� � � ���� � ����� `�P �X �L �W �J �V �D �Y �E �Z ���L 

� , P 3Ѐ
P Pр 3ЭX �P �W �L �V �J �Y �D �Z �E `�Q �X �M �W �K �V �F �Y �G �Z ���M 

� , P 3Ѐ
P Pр 3ЭX �Q �W �M �V �K �Y �F �Z �G `ڜ �V 
����mY � ���mZ � �B m � �C m � ���� ���� �/�D � �D � � �� � �� � � �  �����΀ %� ���`�W )� �8�V � �	�Y �P�*�!��	�Z �����	�Y ����Z �ְ �����\  �)�V �Y � �Z �  ������ �ݭY � �Z �  \������1  4�Y � �Z �  �������1  4��W ��Y � �Z �  ������ �ݭV 
����mY �Y � ���mZ �Z �  ������ [ݭY � �Z �  \������1  4�Y � �Z �  �������1  4��W `�Y � �Z �  ������ �ݭY � �Z �  $��V ��V �Y � �Z � �O�V 
����mY � ���mZ �  ������ �V �W i�W �Y � �Z � �� �Y � � �Z � �W  ������ [ݭY � �Z �  \������1  4�Y � �Z �  �������1  4�`�B m � �8� � � �� 8�B � � �� �C m � �8� JJ� �� �� 8�C � JJ� �� � ��� ��� � �� � � �	� � � � � �� `� i� �� i�� �� � �� L[ӭ i/� ��X � �V � �W �  �˩�	 �� � 8� � � � �8� � �t�;��8� � �0� 8� � � 8� � � m	 � � i � � �� � ��`� i� �� i�� �� � �� L ԭ i/� ��x��� �� �ߍ ��	 �� � 8� � � � �8� � �t�;��8� � �0� 8� � � 8� � � m	 � � i � � �� � ��`H�D � �E � �P �����  �Ԁ�J �  gԀ�J �  ��h`H�F � �G � �Q ����� �Ԁ�K � gԀ�K � ��h`�s 
���m �s �ȹ�m �s ��s �`� � � ��4� �s 
���m �s �ȹ�m �s ��s � i� � ��`� � ��(�s 
���m �s �ȹ�m �s ��s �� ��`�# mI mL mM mB mD mF `�O 
i����� ��� �ߍ ��	 �� ��� �� �1  4�`���@ � � �= ȹ � ȹ � ȭ= ��� |����ݜ1  4���`ڭ i
� �� i�� �� � �� i/� �� L$֭= 
��Y�� �Y� �ߍ ��	 �� � 8� � � � �8� � �x�;��8� � �0� 8� � � 8� � � m	 � � i � � �� � ���`H�Z�O ����F� �� �H �� � � ��z�c 
���mB m �c �ȹ�mC m �c ��c �� �˭H � � � � ��:� �c 
���mB m �c �ȹ�mC m �c ��c � i� � ��z�h`H�Z�b �2 �3 �L���b �c �] �c � �c � �c �^ �� ����ѩ�	 ��  ������ �7�� ȹ7� �ߍ ��1  4�^ ��v�] 
���m m � � ȹ�m m � � �� �� �  �� ؀�� �ـ �������^ �! ������ �7�� ȹ7� �ߍ ��1  4�����^ �^ �c �� m �c �� m �c ��] �c L��z�h`� 8� � ���/�� 8� � �
�Ɇ����� `Zڜ � �� �� �D � �E �  �����H���  �� �hL�حF � �G �  �����H���  �� '�hL�ح ���X�� �
������L�ؠx� �= ȹ � ȹ � ȭ= ���$�� �� �� ��  ������ H����� �z`Zڜ � �� �� �B m � �C m �  ������R ���  ���L�٭D � �E �  ��������  ���L�٭F � �G �  ��������  ���L�٭ ���X�� �
������L�٠x� �= ȹ � ȹ � ȭ= ���$�� �� �� ��  ������ y����� �z`Zڭ ���X�� �
������Lڠx� �= ȹ � ȹ � ȭ= ���"�� �� � ��  ������ �����Ā� �z`��T ���_ �P  �� �ߩ�P �J �L �`��U ���` �Q  �� �ߩ�Q �K �M �`�= ��'�*���> ���� ���  �� 	ۀ���  ����� `�= �#��@����  ����� `�= �#�l�M��T �W��> ���� ���  �� 	ۀ@�N��U �7� �> ���� ���  �� 	ۀ �I��D ����4 ��J��D ����4 � ���  ����� `Z �˭B � �C � ��	 �� �  �ݭD � �E �  ������ �ݭF � �G �  ������ �݈���> � �= � � � �  |�����1  4�F � �G � �Q �X �K �V �M �W  ������ [ݜ1  4�D � �E � �P �X �J �V �L �W  ������ [ݜ1  4�B � �C � ��	 �� �  [��I �O � �H � �I �  �˜1  4� ��z`�D � �E �  �����I� �ݭ_ ��=���J �L �P �X �J �V �L �W �D � �E �  ������1  4��_ �L �C���_   �)�i�P �A��T �J��( � ���P�D ��
�D �G �x����E ��.�E `�F � �G �  �����I� �ݭ` ��=���K �M �Q �X �K �V �M �W �F � �G �  ������1  4��` �M �C���`   �)�i�Q �A��U �J��* � ���P�F ��
�F �E �x����G ��.�G `�Z
��Q�� �Q�� � � � �B�m � ���i � � ����	 ���� m	 � � i � � ��z�`�
��Q�� �Q�� �1  4��`H�Z� �  �� )��&  �ޢ 6�� �d� �
�	 �� � [ݩ #ޮ  ���� 6� �ީ� � �ݭ �& z�h`H�Z
����� ���� � ��$�-�c��b��]��:�8�0�8�7�  �ޭ? ���� 6�Ȁ�z�h`H�" �  ����" ɴ��h`H�  ����h`H�Z� �c��$��b��%��]��&����� ��� �ߍ �� � �B�� ���� � ��� Ȳ�� �� ��� � z�h`�% � �� ���`�' � �� ���`�) � �� ���`�+ � �� ���`�- � �� ���`�. � �� ���`�/ � �� ���`H�& �% h`H�( �' h`H�* �) h`H��+ h`H�P�- h`H�<�. h`H�<�/ h`)?	�`�������7 }=��7 ��8 �< �`H�
� ��� �8  �7  �6  �h`��	 �
� �"� ��� �0  ��� �R ��)J��0#��7�� �7� �ߍ ��	 �1  4�� ���`ڪ)�JJJJ�  �ފ)�  ���`H�Z� � � �B�m � ���i � � �1 � �	�-@ �����Q�����1������	 0��� m	 � � i � � Рz�h`�Z� � � �B�m � ���i � � �0 � ��A ������U�A ����A �A ���	 ����I����	 ���� Эz�`ڢx��� �� �ߍ ��1  4��`�Z�5���� ���� ��z�`� � "�ʀ�`H�Z� � ��L��� � �
 �@� � � �
�6� Z� ���%, P8. . ��. . ��. 8. ��z� �
��0���
 i0�
 � i � ��Щ� 6�LG�z�h`�Z A� E�H�� �(� �  #ީ � �(� �;  �:  �9  �� �7� � #ީ � �7� �8  �7  �6  �h���G���  ���
 6�� �)�� �P� �J�� #ވ���	 �� �0  ����Ω �� � � �� �n� � #ީ� ��� � #ީ� �n� �b�  �ޮ  ���8 nީ��  ��c� � �  ��� � � Ʉ��n� �ĭ i� �����9 nީ��  ��c� � �  ��� � � �n���� ��� 8�� L��� � �� �ީ��  ��L5�L�� �n�� ���z�`� ��  � ��; �8 ��(�: �7 �
��9 �6 ��8 �; �7 �: �6 �9 ���� `� �� ��  �� � � ���� ���  ���H�F���� 轏�� 轏��X �X � �㽏�� 轏�� 轏��X �X � ��ڢ	 6�� 䀩`ڭX 
���� �� �ߍ ��	 �� �1  4��`ڠ �$�<���� ȹ��� ȹ���= ȭ= 
��Y�� �Y� �ߍ ��	 �� �1  4����`�B � �C � ��	 �� �O � �H � �I �  �˜1  4�`�Z� �����L� �= ȹ � ȹ � ȭ= �!���"�� ��� � � � i� �] �s � �s � �s ��s ��	 ��  �����Z� �7�� ȹ7� �ߍ ��1  4�zL��z�`Z������ �!���Ȁ𠁹 �B��!� ��ȩA� �/�����)� �!��@��"��A��@��!��A��"� ��ȀӜb  �� Iթ�	 �� �B � �C �  �O � �H � �I �  �˩�1  4� ��z`H�Z�B m � �C m � � � �n8� � � � �.8� JJ� �������] L�� �����	�] L�� 8� JJ� ������
�] L�� ������] L�� 8� � � � �.8� JJ� ���� ���] L�� ������] L�� 8� JJ� ���� ���] L�� ������] z�h`� �
�s��o�$ ��h�$ �  �x���\� � � � �C m � �=� 8�C � �(�/�  
m  ���� ȭ i�� ȭ 8��� ���� ���  ���  ��`�  �  ��LL�
m  ��� �^ 轓 � 轓 � �^ � �LC���u��	��_�^ �s��] � 8� � � 8� � ��	 �� �0  ���] �B��	 �� ��7�� ȹ7� �ߍ ��1  4�� � �ύ] �8�] �] ���] �] ���^ �  
m  ��^ �� 轓 � 轓 i� �� �� �B m � �C m � �� �� � �  ������  L<�R `�E )�] �� � ��� ��] ����,��� ���E `�Z� ��I��^ ��] �� �� �^ ��٩�	 �� � �7�� ȹ7� �ߍ ��1  4������ 0"��ʈ��ʈ��ʈ��ʈ�ڭ� �� ��] ��^ �] )
���m � � ��m � � �� ��  v�����^ �^ ��] �� �� �� ��I��^ ��] �� �� �^ ��٩�	 �� � �7�� ȹ7� �ߍ ��1  4���z�`� )���� �M�Lr��� �N�Lr�ȹ � � ȩ�s � � � �t �@�u � ��v ��	 ��  ������ �7�� ȹ7� �ߍ ��1  4��w � i� �x �<�y � ��z ��	 ��  ������ �7�� ȹ7� �ߍ ��1  4�� `Zڜ � �� �� �B � �C �  ������R �� ɂ�� ���] ��,��] � ����z`H� )� �5 �=� �& � h`� �� �� ��  � �� � � � � � � � �* �� �� � ���� �� `�� ���%�� � ﭾ � �� �  ���� �� �� � R쭞 ���%�� � ��� � �� �  ��� �� �� � �쭜 ���X�� ����� � ﭢ � �� �  �� ����� � �ﭰ � �� �  P�� �� ͤ � ��� �� Ͳ � 9� �� �`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
������ 轗��� �� )0�� ȱ������ �� Ȍ� �� �� �� � �L�쬫  ��� ��� � ��� ��Ȍ� �� ���� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
������ 轗��� �� )0�� ȱ������ �� Ȍ� �� �� �� � �� �� � �� )������ ��  ��`�� �ɍ� ȱɍ� ȱɍ� ȱɍ� ȱɍ� )
������ 轗��� �� )0�� ȱ������ �� Ȍ� �� �� �� � Ш� �� � �� )��@З���� ��  R쀊�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
������ 轗��� �� )0�� ȱ������ �� Ȍ� �� �� �� � Ч��  ��� ��� � ��� ��Ȍ� �� ���� 
��e��� �e��� �占 ȱ卡 `�� 
��i��� �i��� �卮 ȱ卯 `H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����Ϊ �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����θ �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� �ê�� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� �Ъ�� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� � z�h`� `� `H�Z�� ���%�� ���� �� �� )?
��)��� �)��� ��  ��z�h`�� �* �� `�� ��� ȱ�� ȱ�� ȱ�� )
������ 轗��� �� )0�� Ȍ� �� �� �� � ��� `H�Z�� ���L��� �� �� I�� )��� �� �ڪ�� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� )�� �� )����
�@����� �� �� �( �� �� ��* �� �� �� �� � ��z�h`H�Z�  ��  �휟 �� ��� ��  �� 9� �� P� ����� z�h`H�Z�� � �
�� � ��� �� )?�� �Q�� �K�� 
������ ����� 轇��� ����� �� �� � �� �� �� )������  ��� ����  R� ��z�h`u8
���8
��&
�� �
�� �
��&
��8p
��&8
�� 8
��p
��p
��&�
�� 8
��u8
���8
��&
�� �
�� �
��&
��8p
��&8
�� 8
��8
��&8
��8
��     � �8
�� ��
�� 8
��&
�� �
�� �
��&
��8p
��u8
���8
��u8
�� 8
��&
�� �
�� �
��&
��8p
��u8
���8
��u8
�� 8
��u8
���8
��&
�� �
�� �
��&
��8�
�� 8
��     �u8����8���&��� ���� ����&���8p���&8��� 8���p���p���&���� 8���u8����8���&��� ���� ����&���8p���&8��� 8���8���&8���8���     � �8��� ����� 8���&��� ���� ����&���8p���u8����8���u8��� 8���&��� ���� ����&���8p���u8����8���u8��� 8���u8����8���&��� ���� ����&���8���� 8���     ��8�0 �8�0���0���0���0���0�?p�0�8�0� 8�0�O8�0 �8�0�O8�0��8�0��8�0�8�0��8�0� 8�0��8�0 �8�0�O�0�_�0���0�O�0�?p�0�8�0� 8�0���0?�0� 8�0���0�?�0� 8�0�O8�0 �8�0�O8�0� 8�0�     ���3��3���3���3�?p�3���3��3���3���3�?8�3� 8�3���3 ��3���3���3�?p�3���3��3���3���3�?8�3� 8�3��8�3�8�3���3���3���3���3��8�3 �8�3��8�3� 8�3�     � 8���8��� �8���8��� �8���8��� �8��� ���� ���� �8��� 8��� |��� ���� ���� ���� ���� ���� ���� ���� �8��� 8��� �8��� 8���     � 8���8��� �8���8��� �8���8��� �8��� ���� ���� �8��� 8��� ���� ���� ���� ���� ���� ���� ���� ���� �8��� ����     � p�0 ?8�0�18�0��8�0_8�0��8�0��8�0��8�0O8�0��8�0��8�0��8�0O8�0��8�0�_8�0�Op�0 ?8�0�18�0��8�0�_8�0�8�0��8�0��8�0�O8�0�8�0��8�0��8�0�O8�0�8�0�?8�0�18�0  p�0     � ��� ��� ��� ��� ��� ��� ��� ��� �������&��8��     � ?�� :�� /�� '��     � u�� `�� P�� :��     � ���     � �
�1� /��1�     �1�t����� 4�D 4�j�z 4� 0���?��_�o����    �D �D �D �D 0�_�o��� 0�   �( �  �    �_�    �

		�
	 �
�



	�			�
	
	 �m�}�w���]����I�  ����  ��1�  ��  {������������������?�J�HIcSCORE$SCORE$CONTINUE$END$PAUSE$SELECTcACTOR$ENERGY$EXIT$PUSHcSTARTcKEY$HUNT$OWEN$DALE$NEWcHIGHcSCORE$SCORE$ENERGY$ccNAMEccHUNT$HEIGHTcc7M$WEIGHTcc12T$ENGINEcc80KHP$ccNAMEccOWEN$HEIGHTcc9M$WEIGHTcc15T$ENGINEcc70KHP$ccNAMEccDALE$HEIGHTcc12M$WEIGHTcc21T$ENGINEcc90KHP$ENTER$PROGRAMcBY$SONGcQI$MUSICcBY$XIAOcLIWEI$GRAPHICcBY$ZHANGcLI$�����������������������������'�2�>�L�Y�d�p�~���������������������(Fd @
PE@0#2((# x�hLF�F�G,H�HlIJ�J�f,g�glhi�llmn�nLoL`H'�'�(()�`lclclclclclclc�5H6�$�%�a,b�b�b�b�b�b�E�iLj�jd�d�)h*+�+H,�,�-�k,lLe�e�&�-�k,l�&$L%$L%(.�.h/0�0H1�1�2(3�3h45/�/�o����/�o����/�o��BC�CLK�KLlL�L,M�M�MLN�NOlO�O,P�P�PLQ�QRlR�R,S�S�SLT�TUlU�U,V�V�VLW�WXlX�X,Y�Y�YLZ�Z[l[�[,\�\�\L]�]^l^�^,_�_�_,D�D�D�DLE8   9   : "88 "99 "::   .8"8.9"9.:":8 89 9: :
D
E 
F(
GHI J(K2L2M 2N(2O  ��  �        ��  ��������pB�B,'����� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                    a� �c�