�  T���������  T�0�#2� �#�0�2GGGGGGGG���������WGGGGG���������U UUU���U UUU���U UUU��������������������������������������������*� �������*��������7�7�k��{�_���������W�z�_�����sos�խz�_                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �0��?�:�����5���u���u���������;�U��U��W?  �                                          ���������������������5���u���u�����������U���U���W������������������������������������������������� ��� �> ��� \U5WU5W�� W_ ��7 �W� |�� �� �� ���  �:  �                                 ����������������_U5�WU5�W���W_�������W���������������������������������������������������������  ?  ����U?��U���W���_��W]���]���\��z_������?�  �                                             ����������U���U���W���_��W]���]���\��z_�������������������������������������������������������� �?  ��  �� �� �� �W= {�? ��? 0�� ���\U��\U5 ��? �� �� ��                                ����������������������W��{�������?������\U��\U���������������������������������������������������? ��� l��������p��p]� 0\� 0\� �U�  ��  �[�UY�UY��j��}����U�  ��  /�  �� ܣ �� ����������o��������������]��?\��?\���U��������[��UY��UY���j���}������U��������������������������    ��? ��� l��������p��p]� 0\� 0\� �U�  ��  �[�UY�Ue5̪���������UU? ��<�����?���������������o��������������]��?\��?\���U��������[��UY��Ue�Ϫ�����������UU���������������������                    ��? ��� l��������p��pU� 0_� 0T� �U�  ��  �[�UW0�V0����������� ����������������������������o��������������U��?_��?T���U��������[��UW���V�?���������������� �� ��: ��� ��� ��� \�� \�? W= W5 p�? �� p�5��V50\U0\���� �� �U� ��? ��: p� ܨ �� ��  ���������������������_���_���W��W�������������V�?\U�?\�����������U���������������������������� ��? ��? �= �U= _u \u5 |U? p� �W �� ��  �� �� �� �: �? k� �� �� ��  p� pU �� ����������������U��_u��_u��U������W�����������������������:���?��k������������������U������    �� ��? ��? �= �U= _u \u5 |U? p� �W �� ��  ��? ��� ��� ��? �� k� �� �� ��  p� �� ��������������������U��_u��_u��U������W������������������������������k�����������������������?  ��  �_ �U u5 _}5 _U9 |U5 ��     �0 �0 �� � � | �� �� �� �� �� � �� ���������_���U��u��_}��_U��U������ �� ���0���0������������|������������������������������    �?  ��  �_ �U u5 _}5 _U |U ��   0 �� �� �  7 �?   �� �� �� �� � �� �������������_���U��u��_}��_U��U������ ��0����������� ������� ���������������������������� 0  00 �0 �� �� p5 0\= �\: �_5 �z	 ��5 ��? �� �� �: �? �� �� �: � � \ �? ����? ��0�����������p��?\���\���_���z�������������������:���?����������������������_������� � � 0 0�� 0 � 0 �0 ?0�� �p� �s� �~� ��% ��� ���?���û������?��0 ��? �� �: � � \ �? ����� ��?���? ��? ��? ?�?����p���s���~�����������������û�������������������������������_�������            �� � �  �0 30 30 �    ��  p�  |�  ��  �] W _� �� �� �� �� <�  �� �����������������������0��30��30��� �� �����������������]��W��_���������������������������        �� � �  �0 30 30 �    ��  p�  |�  �� ܗ W� _� �� �� �� �� ?� � ?� �������������������0��30��30��� �� ����������������ߗ��W���_��������������������������������� ��? ��? �� �_� ��0��0�W� �U5 �W= �� \W \W \] |u �} \� \� \} \U �� ��  � �� �����������������_����0���0��W���U���W������_W��_W��_]��u���}��_���_���_}��_U������������������    �� ��? ��? �� �_� ��0��0�W� �U5 �W= �� \_ \�? |U� �W� \�? \U \� \U \U �� �� �� ���������������������_����0���0��W���U���W������__��_���U���W��_���_U��_���_U��_U��������������     � ��? ��� �?� �� �0< 0< 0< ? 3 �  �� ��  <� � � � ;�: �: �� ��   �   �   � �����������������?������0��0��0��? ��� ����������?������������;��������������������������         � ��? ��� �?� �� �0< 0< 0< ? 3 �  �� ���<����� � ;�: �: �� ��   �   � ���������������������?������0��0��0��? ��� ����������?������������;������������������������������        ��������������������W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�W�����������������������������  Z  Z���^���^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^"  ^"  ^���^���^���_���_UUUUUUUU���Z���Z  Z  Z���^���^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^bU^"  ^"  ^���^���^������������������������        UUUUUUUU�ꯪ�ꯪ�������� �} �}������p�7p�7������7�p7�p������������        ���������������� �  � P�WUU�V��������UUUU��WUUUU��WUUUU��WUUUU��WUUUU��WUUUU��WUUUU���UUUU�������P�WUU�V �WUU�  �����  �  � P�WUU�V��������UUUU��WUUUU��WUUUU��WUUUU��WUUUU��WUUUU��WUUUU���UUUU�������P�WUU�V �WUU� ����������������UUUUUUUUUUUUUUUUUUUUUUUU��������      ����������������      ��������UUUUUUUU����������������UUUUUUUU��������UUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUU��UCyU�W��WCyժ^u�WCy�U^5�WCy�@^5�WCy�@^5�WCy�@^u�WCy�U^��WCyժ^��UCyU�WUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUUUCyUUUUU���UUUUU5@�WUUUU5 �WUU����������������        ���������������� �  ��RU�RUU��RU�RUU��RU�RUU��RU�RUU��������������������������������������������������UUUUUUUUUUUUUUUUU�����jUU�_UUU�UU�UUUU�UU�U�V��UU�U��j�UU�j�Z�UU�Z�V�UU�UUUU�UU�_UUU�UU�����jUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�����jUU�_UUU�UU�UUUU�UU�U�V��UU�U��j�UU�j�Z�UU�Z�V�UU�UUUU�UU�_UUU�UU�����jUUUUUUUUUUUUUUUUU���������������� T  U   P  T  @  P ��������UUUUUUUUUUUUUUUQVUUUQVUQVUUUQVU�UUUU�UUUUUUUUU��������������������������������UUU	 \UUUU����UUUU�  �UUUU�  �UUUU����UUUUU	 \UUUUU	 \UUUUU	 \UUUU����UUUU�  �UUUU�  �UUUU����UUUUU	 \UUUUU	 \UUUUU	 \UUUU����UUUU�  �UUUU�  �UUUU����UUUUU	 \UUUUU	 \UUUUU	 \UUUU����UUUU�  �UUUU�  �UUUU����UUUUU	 \UUUUU	 \UUUUU	 \UU��������U�QUU�FUU�QUU�FUU�QUU�FUU�QUU�FUU�QUU�FUU�QUU�FUU�QUU�FU����������������UUUUUUUUUUUUUUUU      `TUUUUUiTUUUUUiTUUUUUiTUUUUUiTUUUUUiTUUUUUiTUUUUUi������j�������jUUUUUUUUUUUUUUUU      �FUUUUU�FUUUUU�FUUUUU�FUUUUU�FUUUUU�FUUUUU�FUUUUU���������������UUUUUUUUUUUUUUUU  �   UU�QUU�FUU�QUU�FUU�QUU�FUU�QUU�FUU�QUU�FUU�QUU�FUU�QUU�F�����������������<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                    0 < ����< 0         ����      ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�                               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �������������������������������������?                                      0  LUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU5  LU��U��U��U������U�UU��_�����U5  LU���U��W��W����z���z��zUU�z�ުz��U5  LU���ժ�^��^����z��z��zUU��ުz뭪W5  Lի���^��z����z���z��zUU��������W5  L��W��z�^��z�WU�zUU�^��zUU�U��^UU�U�W5  L��UU�^�_U�z�WU�zUU�W��zUU�U��^UU�U�W5  L��UU�^UU��z�WU�zUU�W��zUU�U��^UU�U�W5  L��WU�WUU��z�WU�zUU�W��zUU�U��^UU�U�W5  LU��W�WUU��z��������W��zUU�U�������W5  LU��^UUUU��z���ު��W��zUU�U����z뭪W5  LU��z�WUU��z���ު��W��zUU�U����z��U5  LUu�z�WUU��z��������W��zUU�U�����~U5  LUU��WU���WU�zUU�W��zUU�U��^UU�^U5  LUU��^Uժz�WU�zUU�W��zUU�U��^UU�zU5  LUU��^�ߪz�WU�zUU�W��zUU�U��^UU��zU5  L���z����WU�zUU�^��zUU�U��^UU���U5  L�����zU�WU�zUU�z��z�������U�U5  Lժ�zժ��zU�WU�zUU�z��z�z��ުz�U�W5  Lժ�^U���zU�WU�zUU�z��z�z�z�ުz�U�W5  LU��WU���U��WU�UUU����_����U�W5  LUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU5  LUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU5  �������������������������������������?  �������������������������������������  �������������������������������������   ������������������������������������    �����������������������������������>    𪪪�������������������������������    �����������������������������������     ����������������������������������             3�0   ����� �3                    � 00  ������ 03                         ������? 0030                        �ת�> ���                   0     �ת��  3�                   0   �? �������  <��                   �   � �������    00                   �    � �������                       �    � ������� 0                      �   �  ���ת�� 0                      �   0  ���ת�� 0                      �     �������                            �������?                       +    ���������                        �   ��� ����                          0   ��  �                         0   ��  ��<   �                     0   �?�  ��   �0                     0   ��C� �    �                    �   ���� 0 �                    � �  � <�� � 8  ��                 � �?  ��@ �� �?   ��                � ��  �<@ ��?�?   �>                � � � @ �   �   �                � ��    � � �  �                � ��  � " �  �                �>�O	    � ��     �                ���S      �0�    �               ��T   <0 ��3�  <  L�               �PU   0���3�  0  C�               VU�    � � �3  
 ��P�               [jU*     0��3  
0���               l��"  (  ���3 ����  ��               l�*
  (  �  ��0 ���� P%�               l��   � �:0 ���CUA�               �UU    �0 ��(�> T�                �UU���*  0��� �����V�:                �V���"  0���  (��VV��                 k(*  
  ���: C ��Xf��                  l�**�
   ��Q  je���                  ��V �    p �����                   ��� �   �<L  ���?                    ���*     ��  ���                     ����
           �                       ���
       P  �                       ���       P   �                        �T         �                         ��e        �                         � �   @    �                         � T
        �                           �       @�                           �$       ��                            *       ��                           @%     ����                           0  �   �� ���                           0  �   ����                           0  T
   *����                           �  @
   �**`:                              �    �
H>                              �*     P                            <  ��    @�                            � ��   U�                            ��< Z T��                             �����@���                              �����ZU���                              l������_�                              l@�������                              l@��?��k�                              lTU�> ���                              � T�>  ��                              � T�>  ��                              �  �>  �:                              �  �>  �                              �V  �>                                   [  P>                                   [ P>                                   l P>                                   � �>                                   �V �                                    [ �                                    o��                                    ���                                     k�?                                     �U>                                     k�>                                     ��:                                     ��:                                     ��:                                     ��:                                     ��                                     ��                                     ��                                                                                                                                                                                                                                                                         �                                      0 �? �����30��? 0���            �� �� 00000003  <0030            3� ��< 00000003  0000            3� ���� 0��00�00�� 0�?�            �� �� 00�? 3030  0 0             0 �� 0000 30�0  0 ��             � �? 000�30���? ��<�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ���ة��  ��� � �A � � �B � �ߍ& ��" � t ����+ ��, �� � �+����, ��� >��#  �� �� �� �� �J XL �H�Zx�� ��� *� =�' )���# �$ �% (z�hX@@                                                                                                                 ��ߍ&  j© �J  �� �� �詟�& ���  � 'ĭ� ��� ŭ� � �L� �ǭ� � ��LR��� �� ���J  � m� *� ��  �� ĭ� �(�� 
��N�/ �N�0 �� �/�5 �4 �6 � 	�  �� � \˩� � �� ���  �� @� �� )� F� �Ӝ3  �­� ���L��� � � �� �� �Ѐ z٭� �������  �� �� ���� �� �L�LR� Q٭� ��� �ϭ� Ɉ�BLR��� ��� � � �Ѐʭ3 ��  �� )� @� �� d� ���� �� �L�LR���L���  ��L�Hک��J  � m� *���  �� � � � �(� � ��� �p�2 � � �  �� �� �� �ݩ���  � E� �� �� ������ ީ �J  �� �� ���h`H�Z� �� ���  (����2��� �� ��� �� � �� r׭� �L�� �� \� �� �� d�L�����2��� �� ��� � � �� r׭� �L�� �� \� �� �� d�L����� 7� 7� ��L���������������  7� e� �� \� �� �� dѢ �����L�������������� � �ۀT��1���� �I�
�? �#�? �����? ��? ����? ��? �? ��? �? �
�@ ��@ � ݩ�? �? �0�@ z�h`H� ���� ���� �� ���� h`H� �J  �� �� �� >�� ��� �  Gީ(� �� � Gީ� �<� � Gީ� �P� � Gީ(� �"� �%�1  �ޜ�  �ɿ�< �ޭ� ���"� �(� �%�1  �ޜ� �ة"� � i� �%�1  ��� ���������= �ޭ� ��"� �P� �%�1  �ީ�� ���"� � 8�� �%�1  ��Μ L����L��h`H�Z >���� �� �� �	�1 ��� � �1  �ވ�� i � �� ��ީ� �g� �%�1  ��� � ��1  �ީ�1  �ީ�1  �ީ�� �� � Gީ&�1 ��� ��  �� �� �� �ީ&�1 �� ��  �ޜ; ���D ��C �
�� �  ����Lxƭ� �$�C�; �L���C �C � ڬ Z�C � �D � �$�1  ��� � � �C z� �� �; ���%�L�ǭ; ��L�ǭ� �1 �; i7�� �; � ڬ Z�C � �D �  �ޭ �C z� �� L�����8 �ޭ �
�i� �&�1  �ޭ� i�� L��8�� �&�1  ��Ο L�����8 �ޭ ��8�� �&�1  �ޭ� 8��� L��� � �&�1  ��� L�����J �ޭ �� i`� � � �&�1  �ޭ� i�� L��8� � � � �&�1  �ޭ� 8��� L�����I �ޭ �n��� � � �&�1  �ޭ� 8��� L��i � � � �&�1  �ޭ� i�� L�����L�ũ �� z�h`H�Z� �� �� ڊ
����- 轨�. �� �� �-��������� ����� �� ���� �� L�ǩ �� �� z�h`HZ _ʩ�� �8 �; � �9 �T�:  �ʜ8 �; �U�9 ���:  �ʜ8 �; ���9 ���:  �ʜ8 ��; � �9 �T�:  �ʜ8 ��; �U�9 ���:  �ʜ8 ��; ���9 ���:  �ʜ8 ��; � �9 �T�:  �ʜ8 ��; �U�9 ���:  �ʜ8 ��; ���9 ���:  �ʜ8 ��; � �9 �T�:  �ʜ8 ��; �U�9 ���:  �ʩ�8 ��; ���9 ���:  �ʩ�8 �; ��9 �T�:  �ʩ�8 �; �V�9 ���:  �ʩ�8 �; ���9 ���:  �ʩ�8 ��; ��9 �T�:  �ʩ�8 ��; �V�9 ���:  �ʩ�8 ��; ���9 ���:  �ʩ�8 ��; ��9 �T�:  �ʩ�8 ��; �V�9 ���:  �ʩ�8 ��; ���9 ���:  �ʩ�8 ��; ��9 �T�:  �ʩ�8 ��; �V�9 ���:  �ʩ�8 ��; ���9 ���:  �ʩ�� ��� � �  =ʩT� �  =ʩ�� � ��  =ʜ �S�  =�zh`  ڭ iU� ������ � ��� ��`H�Z�; �; ��
����/ 轼�0 � � �/������; ��z�h`H�Z�; 
����/ 轼�0 �9 �8 �/�m� ��: ��z�h`H�Z� � � � �  ����(�� �� i.� ����L��� � ��� L�� n� )�z�h`Hڢ � ��<���h`HZ ˭� 
����/ ȹ��0 �� 
��/�- ȱ/�. �� 
��-�/ ȱ-�0 � �/� ���Ȁ�zh`HZ� � ���� ȹ � Ⱦ ȹ 

��  ��Ȁ�zh`H�Z��� �� i��   ��� � i� �
���� �   ����3�� �� i� ����� � �� 8�V� �� � �� L���� �� �� i� ����� � �� 8�V� �� �   ��� � i� �
���� �   �z�h`H� �(� � �
� ��  �ߩ
� �� ��  �ߩ8� �� ��  �ߩ� �� � Gީ#� �� �c�1  ��h`H�� �� �� ���� Gީ!� �� i�1  �ީ%� �� i�1  ��h`H�Z� )͠ �݈���8� �� � Gީ8� �� �� i�� �i Gޠ �݈����� )�z�h`Hک8� � �(� �� ��  �߮� ��8� � � ��2  ��� � ����h` o� ��`Hڭ� iB�2 �� � � ߭ i� ����h`Hڭ� iB�2 �� �� � ߭ i� ����h`H�� 
i�2 �� ��  ,��2 ��  ,ߜ h`H��  ��h`H�� �� �� �� ��  ��h`Hڭ9 � ���  ��� � �: � �� �� )�� � ������ H ��h� �ҭ H ��h� ���  ���h`Hڭ: � ���  ��� �� ��� � ������ H ��h� ��� � H ��h� ���  ���h`Hڭ9 � ���  ��� � �: ���� � ������ H ��h� �ح H ��h� ���  ���h`H�Z��P� �� �� �(� �  �ߠ �݈���`� �� �� ������ Gޠ �݈���йz�h`HZ hͭ� � �̭� 
i��  �ͩ$�9 ��:  � b� oͭ� 
i	�� � �݈�� �͠ �݈�� o���  �� ��zh`H�Z���J  � m� *���  �� ����  �Ω�:  b� �ͭ� ��1� �� 
i	��  �͠
 �݈�� o���  �ͩ�9 �$�:  ��L�Т o͠ �݈���� 
i��  �͠ �݈����ݩ� ���  ��� � � �� �� )�� � ������ H h�h� �՜� �� ���� ��� � ��  h̀4���� � >�
 �݈���L� �� � Gޠ
 �݈����۠ �݈��� �J  �� �� ��z�h`H�Z���J  � m� *���  �� � ��  �έ� 
i	��  �͠ �݈�� o���  �ͩ�9 �$�:  �Π �݈���� ��/� >�
 �݈���L� �� �
 Gޠ
 �݈����۠ �݈��� �J  �� �� ��z�h`H� �� )i�2 �� � �� �  MڭI � � ��h`H�� � �� �  �٭ i� ����� �  ��h`H�� )�	�� �� �� 8�� �� � ��   ڭ� )��3�� �
 �� � �
 8� �(��
 8�U�
 ����� �� �� ����� h`H�� )�	�� �� �� � �� i� ��   ڭ� )��5�� �
 �� � �
 8� �(��
 8�U�
 ���$�
� �-�� �� ����� h`H� )� �� �
�� �U�Lӭ� � �� 8�U� �� � ��   ڭ� )��G�� � �� 8�T� �� � ��   ڭ� )��! �ѭ� 8�U�� ��� �� �� )���  dр� 	�� h`H� )� �� ��
�� �U�L�ӭ� � �� iU� �	� ����� � ��   ڭ� )��d�� � �� iV� �	� ����� � ��   ڭ� )��5 �ѭ� �� �� iU�� �	�� ������ �� �� )���  dѩ��� �� 	�� h`Hک���  �� \� �� dѢ �ҭ )�� ���� �ӭ )� �h`H ӭ )�� Ԁ�h`Hک��  (����
 �ѭ� �,�0���
 ҭ� ��"���
 �ѭ� �����
 ҭ� �� �� �� �� d� ���h`H�Z�� �� �� )����L�ԭ� i�� �� �� ��� 8��� �� �� ��  �ԭ� ���;� ڊ
����/ ���0 � �/�� �ȱ/�� �������� L����� �� ������ z�h`H�Z�� �� �� �� �� �� �� �� �� �� ���L��
����/ ���0 � �/������� L�ՠ �/� ȱ/� ȱ/�� ȱ/�� �� �)�� � � �� � �� ��@� 8�U� �� � �ܭ� )��� �� � �� L�խ� 8�
m �� � �� z�h`H�Z��� �� ���Y
����- ���. � �-� ȱ-� ȱ-�ȱ-�� ���   �� ���   ����� �� �� 8�V� ��� � ��z�h`H�Z�� ���l
����/ ���0 � �/� ȱ/� ȱ/�� ȱ/�� �� �� �֭� �5� � �֭� �(� � � �/ȭ �/ �� \� �խ� �� Ҁ ��z�h`H�Z� H� H�0 H�/ H�� �� �� ��� i� �� �� �+��   ڭ� )��LY׈�L ׭ 8�U� ��� � �ح� ��  ڭ� )��U��� 8�
m �   ڭ� )��9�� ���� i� �� � ��� 8�� �� �   ڭ� ����	������ h�/ h�0 h� h� z�h`H�Z���� �� � �
����- ȹ��. �� � �-����� ����  ���� ��LMٍ ȱ-� ȱ-�� ȱ-�� �L]ح ��
� �U�L�ح� 
�� � iU� ����� � � H� H��   ڭ� )��h� h� L���� �� �� �٠ h�-� � �h�-� � � H� H �� \�h� h� ���� �� L�׭ ��
� �U�L�ح iV� ����� � ��   ڭ� )��D� ��   ڭ� ��4� � � �-ȭ � �-� H� H �� \�h� h� ���� �� L]ح� ���� �Lש�� � � � � ��-�� �� ���   �� ���   ����� �� �� 8�V� ��� � �� �� dѩ��  �0 �݈��� �� z�h`HZ� �� � � �����ȹ �U�
��Ȁ���� zh`HZ���� � � ���p� ȹ � ȹ �� ȹ �� ��,�� 
�� �� � �5�� � �0i� �(�� �� �� ��� � ��� � �i� �Ȁ�� �� ���  �zh`H�Z�  MڭI � ���   ڭ� �2  ��z�h`H�Z� 
����/ 轼�0 � �� ��� �/��/�� z�h`H�Z���I � 8� �
 � � � � � � ���舀��
 �U��8�U��� �(�� �I ���� z�h`H� >�2� �� �	 Gީ� �d� � Gީ2� �� �%�1  �ޜ;  �ɿ�< �ޭ; ���� �2� �%�1  �ޜ; �ة� � i2� �%�1  ���; ���������? �ޭ; � ��� �d� �%�1  �ީ�; ���� � 8�2� �%�1  ���; L����L�ڭ; ��L�� >�� �.� � Gީ� �V� � Gޢd ����� >�F� �� � G� ����� �J  �� ���h`H� �J  �� �� �� )� �@� � �(� �`� �  �ߩ� �H� � Gީ� �d� �	 Gީ� �x� � Gީ� ��� �
 Gީd� �� �%�1  �ޜ3  �ɿ�B �ޭ3 ���� �d� �%�1  �ޜ3 �ح i� �� �%�1  �ޭ3 i�3 �����LF����? �ޭ3 � ��� ��� �%�1  �ީ�3 ���� � 8�� �%�1  ���3 L?���L?ܭ3 �!�� �� 	�  � m���J  *� �� d�h`H� )�Llݩ��� �4 ��5 ��6 �� �� Llݭ6 ��6 �6  �ݍ6 �.�5 ��Y�6 �5 �5  �ݍ5 ��4 ��Y�5 �4 �4  �ݍ4  n�h`H� H� H� )�L�ݩ� ��� � Gީ� ��� �4  �ީ� ��� �5  �ީ#� ��� �6  ��h� h� h`�7 )�
��m7 )��7 ����7 )�i	�7 �7 `�Z�0���� ���� ��z�`�  ���� � �� �� �� �`H�  ����h`ڮ� �   7�����`H�> �> �> �/��h`H�Z
��,�< �,�= � �<�$��a��b��c��d�8�7�1  ��Ȁ�z�h`Hڪ)�JJJJ�1  �ފ)�1  ���h`H�1 �a��$��b��%��c��&��d��'iH�2 �  ��� � h`� � �$�1  ��`H�� � �� � �  E�h`H�� � �� � �  E�h`H�� � �,� � �  E�h`H�� � �� � �  E�h`H�Z�2 
���� ��� � � �� m � � i � ��� m � � i �  W� � ڱ� � ���1�
���Q��� ����� �%� i0� � i � � m � � i � ��z�h`H�Z W� � �� � ����U� ������ ���� � � � ��� ���� �� i0� � i � ��z�h`H� � � ��� �(�  ��h`Hڮ �x�m � �"�i � �h`H�Z� � �9 � �: �2 
���� ��� � �)�JJJJJJ�  ��)0JJJJ� �  ��)JJ� �  ��)� �  ������ � � � L��9 � �: � z�h` p� ��`H�Z� � ���  � )��,      ��      ��      � �� � �-   ���- ��� �M �z�h`Hڮ �x� � JJm � �"�i � �h`H�Z�2 
���� ��� � � �� m � � i � ��� m$ � � i � z�h`H� � �� �! ����U�! ������! ����! ��# � JJ�" � �(� )�  � )� � m )i8� �  ��" � )� �8� � � � � H ��� � � � ��" � ��# � �� i� � i� �# �" �� � � ��� � ��� � � �h� H� � LW�hh`H�Z�! �# � � ���1�
���Q�z�h`H�Z���& � �� ���� �� � �� �  �� �ݬ� �r��� ���� ���� �� �� � �� �  ���� �� �� � �� �  ��� �D�	 �� ��L"� �� �ݭ� � �� �  ��� i�� �  ��� �  ��� 8��� �  �� � m� z�< �݈��z�h`H�r�2 � �� � �� � �  E�h`H�q�2 � �� � �� � �  E�h`H� �� ��  ��h`� �J �K �L  �� �� � � � � � � � �* �� �� � ���� �� `�K ���%�s � ��l � �m �  ���s �s �n � x�L ���%�� � ��y � �z �  7�� �� �{ � ��J ���X�K ����W � ��P � �Q �  �L ����e � ��^ � �_ �  m��W �W �R � ��e �e �` � Y歛 ��� �� *�`�M �N�P ȱN�Q ȱN�R ȱN�S ȱN�T )
��v��U �v��V �T )0�Z ȱN����� ȌM �W �X �R � �L��Y  ��� ��N � ��Y ��ȌY �M ���i �j�l ȱj�m ȱj�n ȱj�o ȱj�p )
��v��q �v��r �p )0�u ȱj����� Ȍi �s �t �n � �� �K � �� )�����L �v  ��`�v �w�y ȱw�z ȱw�{ ȱw�| ȱw�} )
��v��~ �v�� �} )0�� ȱw����� Ȍv �� �� �{ � Ы� �L � �� )��@К���K �i  x倍�[ �\�^ ȱ\�_ ȱ\�` ȱ\�a ȱ\�b )
��v��c �v��d �b )0�h ȱ\����� Ȍ[ �e �f �` � Ъ�g  ��� ��\ � ��g ��Ȍg �[ ���� 
����� ���� ���N ȱ��O `�� 
��$��� �$��� ���\ ȱ��] `H�Z�S )?	@�� �S I��-� �� �X �U��T )@��J��� �� �Z �8��Z ��T )0�Z ȌX �U����X �T �X �� � z�h`H�Z�a )?	@�� �a I��-� �� �f �c��b )@��J��� �� �h �8��h ��b )0�h Ȍf �c����f �b �f �� � z�h`H�Z�o )?	@�� �o I��-� �� �t �q��p )@��J��� �� �u �8��u ��p )0�u Ȍt �q����t �p �t �� � z�h`H�Z�| )?	@�� �| I��-� �� �� �~��} )@��J��� �� �� �8��� ��} )0�� Ȍ� �~���΁ �} �� �� � z�h`� `� `H�Z�� ���%�� ���� �� �� )?
������ ����� ��  ��z�h`�� �* �� `�� ���� ȱ��� ȱ��� ȱ��� )
��v��� �v��� �� )0�� Ȍ� �� �� �� � �蜛 `H�Z�� ���L�魅 �� �� I�� )��� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����Ί �� �� �� )�� �� )����
�@����� �� �� �( �� ͏ ��* �� � �� ͆ � ��z�h`H�Z�  ��  ��M �[ ��Y �g  � Y� � m� ����J z�h`H�Z�K � �
�L � ��� �� )?͖ �Q�� �K�� 
��b��j �l��w �b��k �l��x �i �v � �K �L �� )�����L  �孕 ���K  x� ��z�h`H����  �h`SELECTaPLEASE$BEGINNER$SKILLED$PASSWORD$BEGINNER$SKILLED$STAGE$PAUSE$GIVEaUP$CONTINUE$GAMEaOVER$TIME$END$HAHA$OHcc$PASSWORD$CONGRATULATIONS$BYE$PROGRAMMEDaBY$FRANKaGU$�����������������������������#�l�q�v�{���������FINE$READ$PASS$WORD$LOVE$LIVE$JUMP$DROP$TIME$HIGH$WORK$LATH$l�q�v�{��������� ���� �(�0�8�@�H�P�X�`�h�p�x�������������        ���P����p�Ф0����P����p�Ч0����P����p�Ъ0����P����p�Э0����P����p�а0�����`�ȵ0��� �� �0�@�P�`�p�����������к�� �� �0�@�P�`�p�����������л�� �� �0�@�P�`�p� � � �          @HPX`hpx����<;:9  $(,048� � � � �������$�.�8�B�L�V�`�j�t�~������������'�<�Q�j�������� �=�V�o�����������C�l�y������������)�J�g��������!�B�g�������D�m������{ }, ��y� ��}* }* �y( � ��{& w� ��{ w&  ��{, {& {�{$� �w$ w�. ��w u ���{& {& {�{ � � ��y w�� . ��w}� $ * y,�o q o} y ��� 4 ��{ �� ��s  * (0 ��{( * {& , {�y�&� � y�}( , }* }�u" & "� ��u  � � �� � ��y {& y� . �y * �}y ��}*  ��{( } � � �{ }* � {�}( {( } �s s" w�4 �0 ��y$ y$ y. �. ��}( }�{ }� ��} * , }�{ w�. �y w�. 2 ��y$� $� 0 �w y& w� ��{ �(� ��y y* . .�y� * y�$ * �{ }� �{ � {�{ �u { ��� 0 ��w y& w& "� ��{ ( {& , }, �}*  � (�w( {( � �� ��w& &� �� ,�s   �  �4 �w�& , w�& ,  ��s  u } }  � � �4 � �s u  s{ � {�� 2 ��o qy w" � �2 � ��y {( y( } �. * * �u  " } � }* �2 4 �w � "{ }�, � � *�w" w &  � (�. 2 � �y( * y$ &. �y$ y$ ( }. * . �w& y&� &�, *� �w" & "�  � (�. 2 .�  � �Z�_�d�i�n�s� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^_____ ��� ��� ��� �� �� q�� �� ��� ��� ��� ��� ��� ��� ��� �0��     � �� � �� � �� � � � � � q� � � � �� � �� � �� � �� � �� � �� � �� � �0� �     � �� � �� � �� � � � � � q� � � � �� � �� � �� � �� � �� � �� � �� � � � �  � �     � ��!� ��!� ��!� �!� �!� q�!� �!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� � �!�   �!�     � � �!� � �!� q�!� q �!� q�!� �!� �!� ��!� ��!� � �!�  �!�     � ��� ��� ��� �� �� q�� �� ��� ��� ��� ��� ��� ��� ��� � ��   ��     � ��! ��! ��! �! �! q�! �! ��! ��! ��! ��! ��! ��! ��! �0�!      � ��! � �! ��! ��! ��! ��! � �! ��! ��! ��! ��! �0�!      � ��! � �! ��! ��! ��! ��! � �! ��! ��!�!.�! �0�!      � ��! � �! ��! ��! ��! ��! � �! ��! ��! ��! ��! � �! ��! ��! ��!     � ��! ��! � �! ��! � �! ��! � �! � �! �0�!      � ��! � �! ��! ��! ��! ��! � �! ��! ��! ��! ��! � �!   �!     � ��!� ��!� ��!� ��!� �!� ��!� �!� q�!� ��!� _�!� d�!� q�!� �!� q�!� �!� ��!� ��!� ��!� ��!�     � ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!� ��!�     � 
�!� ��!� �
�!� ��!� d�!� q�!� �!� q�!� �!� ��!� �
�!� 
�!� q
�!� d
�!� ��!� _
�!� d
�!� Y
�!� O
�!� K�!�     �.
�!� ��!� ��!� ��!� ��!�@
�!�.
�!�T
�!�}
�!�T�!� ��!� ��!� ��!� �
�!� ��!� ��!� �
�!� ��!�
�!�.�!�     � ��B �� D ��C �� C ��B �� D ��C �� C ��B �� D ��C �� C ��B �� D     � ��C �� C ��B � D �C � C ��B ��D ��B ��D �(�A  (�A     �T�!�.�!�. �!��!�.�!� � �!�T�!�.�!�. �!��!�.�!� � �!� ��!� ��!� ��!� ��!� � �!� � �!� � �!�   �!�     � �
�� /2��     � �� � ��
�     � �� � � � _� �     � ��� ��� ��     � _�� q�� d�� ��� q�� ��� �� ��� ��� ��� ��� ��� ���     � �� ��� �� ��� �� ��� ��� ��� ��� ��� ��� ��� ���     � ��      ��������*��l� �h� �   �h� �   �f� �I� �   �I� �   �f� �   �   


				 �
	�	
 �
�			�


	�


�	����,�H�P�X�:�L�T�^���-�����Y���  �g����c���  ��  k�  ��  +�  ���  Q�  ������#��������w���1�i�y��������������                                                                                                              �� �e�