                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                L)�L�LԀL��L+�Lm�Lx�L)�L��PRESS  START$STAGE $TOP  SCORE $YOUR SCORE $MISS$CONTINUE$END $ONE$TWO$THREE$FOUR$FIVE$SIX$ PROGRAME BY LIHONG$  GRAPH   BY ZHANGLI$  MUSIC   BY HUXUHUI$(��;�/�G�L�U�Z�^�b�h�m�r�v�����H� �� 7ĩ �	�,��2������� ǩ4��9�� ��   �����h`*�H�
��������� ���h`H� �� 7ĩ�Z � �	���2��k���l�� ǭ   ������ �Z �h`g�� �� 7ĩ���� � 삩��(�� � ݂�,��Z��  ���i ��   �����`� �� 7ĩ���� � 삩��(�� � ݂�4��F�� ��4��Z�� �d����2��<��x� kĥ�
��r���r���v���w�� ǭ   �������p�����]  �Lo�ɿ���]  �懥�)��L	�`AUF�� �� 7ĩ���� � 삩��(�� � ݂���F�� ����Z�� ����n�� ��   �����`Hڢ�� �����h`H� ����� �����h`H��Ŝ�"����ś�����Ś��������������h`H� �	���������� ǩo��� 샀�d���� � �� 샭�D�������	 � � ���i��8�� � ����T�ة��]  �< �:��h`�H�H�H�H���������� �h�h�h�h�`H�Z�/���� ���� ��z�h`7�)� 7Ĝ��'���(�� ǭ   �����`��Hd� u� N� �LF� #� �h�`��	��
���D����
��{D��|D��b�轃D� �挩d �L2���6�x��� 24 68 :< >@ BD FH JL NP RT VX Z\ ^` bb`^\ZXVTRPNLJHFDB@><:8642����"��	�d��b���:
��E��E� �`��>���µ���� v�`�H� �	���]��IJJ

��S��� ��h�`�H� �	���(��sE��tE� �h�`���Hid��(�HiU� �ņ���]h�Sh�I`�H u� � 
� �� � ̅�   ����� #� �h�`�\��d���:
��E��E� �`�[��W��� ��`�[��H��� ��`�H��<� �B`� �	���(��5F��6F� �`	l ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              �������������� <             ������������?�            ��            ��           ��           ��          ����          ����          ����          ����            ��          ����          ����          ����            ��            ��            �������������?<             ��������������  ��  �    ��?   ��   �� �? ������ ��?   �?� ��?���������� ��  �������?�����  ���� �   �?���� ����  ������    �?����  ����  ������    ���?���  ���?  �������  ���?�����?�?���?<�����  ���?�������?����?<�����  ���?���? ���?����?<����    �����?  ��������?<����    �?����?  ��?������?<�����   �?� �? �  ��?����?�??0���  ��� �? ��� �����?�?? ���?  ��? � ��� � �� ?  ��?   � � �� ? �(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ������                                ��<��  ���                           �<�<��  �� �                        ��<�<��  �� �                      ��� �<�<��  �� �                    �� �< �<�<�� ��� �                    <  � �<�<�� �?� �                   �?  � �<�<��  � �                  � ?  � �<�<��  � �                   0 ?  � �<�<�� �?� �                   < ? �� < <���  0� �                   < �?��  ? @��  0�                     ? �?�<  TU5|U0<                   �?? ?�<@ _UU5|UU5<                �� <0? ?�<T _UU5|��?<                0 ?<0? ?�|U _�_5|��|               0 00? ?�|U _�_5|�  |�              < 0? ?�|U _5_5|�  �W             < �? ��|U _5_5|��?_�_�              < �?@�_��U�_5_5|UU5_�_�              ? � ?P�_��U��_:�:���5_5�              ? �� ?U�_5�UU�:�:���:�5�              ? 0� ��_5�V��:�:���:�:��              ?  � ��_5��:�?���?�:��              ?  0 _��_5���?�����?��             �?  0�_���:���>�      ��?             �  �_���: ��                         � @�_���: ��                         � P�_���:                             � T�_���:                             �@U�����>                             �PU=�����                             �UU������          �?                 �OUU�ï���         ��U�>                �WUU�ϯ�          �WUUU�               �WU�����          pUUUUU=               �WU�����          pUUUUU�?              �W�����?          pUUUUUU�              �W�����          \UUUUUUU             �������          \UUUUUUU             ������      ��   \UUUUUUU5             �����>     � �  \UUUUUUU�             �����  �? �    \UUUUUUU�             ����� �� �    \UUUUUUU�             ���?�  < � �    pUUUUUUU�             ���  �?  ��  pUUUUUUU5             ��� �?  ��  �WUUUUUU5             ���  �   �   �WUUUUU             ��  � ��   p}UUUU�             ��   � ���   p�UUU                   � �0�     \U��U�                    < 00�      \UUUW                 �? <�00�      �UUU�                 <0�?�00�UU�   �WU�                  0?��O��U_�   �  �U�                  0� U��U�   �   W�                  ��UU��U��   p@��                  � �WUUտ��U  �P��                ��  �WUU����k  �14 �                �0 @�WU�����  L<= �                �  T�W������  =                  � PU��꼪���:   0                � UU���������:  T                 �PUU��:������?   P                 �UuU��:��?��       �                �_Uu���:�� � �     �U?�?             �_U����:��     �     |U�?�             �_U����:��      �     pU� �             �_U����?�?      0     pU� �             �_U����        0 <   �UU�             �_�����        0 �   �UU�             �_�ϯ�?         0 �   �UU�             �ï         �� 0   �UU?�             ���       ��]�    �UU3�             ��       pU]U�   �U�0�             �� �        \UuU   �uU�0�             ��          WUuU   puU=0�             ��         �UU�U5   _]U0             ��         \UUU_5  �U]U0             ��?         \UUU�� ���W�              ��         WUUUUU�WUUU5              �� ����   WUUUUUUUUUU5�              ��  ����   WUUUUUUUUUU�  ��                 �;  �UUUUUUUUU���  ��                  �  ��_UUUU������                     �� �pU������  �  ��   T          �����0  ������   ���  �  �
@U	         ������?� ���  ���U  �  `%PU!             ���?�  ���UUUU5 � 0  P�T!             ��0����WUUUUUU5 �� �� @             ���0� WUUUUUUU5�   h� �         ������� WUUUUUUU�W�   V  �         ������� WUUUUUUU}UU �U                � � WUUUUUUU]UU5 ` T�             �  �?  WUUUUUUU_UU5 ` P �            �?      WUUUUUUUWUU�   
%         ����      WUUUUUU�WUUU�  Z
         ����   �? \UUU���W�UUU����                  �� \UU�WUUUWUU Z T                 ����UU}UUUU\UU5�U P�                 ��� WUWUUUU\UU5�@ T�                 ��� \�UUUU� \eU�` U�                 ���> p_UUUU� \eU�`  Pd                 ���> �UUUUU� WiV�  Pe                 ���> �jUUUU5�UZVՃ*@PY                 ���� \�UUUU5�U�V�#�  �                 ���� �WVUUU5_�U�# T%                 �����_VUUU�\UU�K dU&                �����0 \VUUU pUU�U ��%                ����� pYUU� �UU�T 	V	                ����� pYU�  �_իPA	�                ����� pYU?   �U��PU                  �����  pY�    ���� T�                   �����  pY=    ���>%
                   ���z5  pY    ����(                    ���{5  _�        �P                    ���z5 ��        �P                    ���{5           ��                     ���z5            *                     ���z5�                                  ���z5<                                  ���z5                                  ���z�                                   ���z�                                   �����                                   �����                                   ����5                                   ����5                                    ���                                    ���                                    ���                                    ��                                                                                                              �                                       ����������?� �?�           ��0 30 � � ��  ��           �0 30 � � ��  ��            �0 �003 ��??�?� ��            �0 30� �� ���   ��            ��0 30 � ��0   00              �� ���?���� ?� �            �                                                                                                                                                                                                                                                                               Q  ����   ����   ����       �      �      �   �      �      �            0      0      0 �     ��     ��     �0                       ������������������������0@  P  @  P  @  P 0 U  @   U  @   U  @ 0 T  U   T  U   T  U ������������������������pUUUUUUUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������������������������������������������������������������������         ����         ����_EUEUEUEUEUEUEUEUEUE����^UUUUUUUUUUUUUUUUUUU����          ����@@@@@@@@@@����^UQUQUQUQUQUQUQUQUQU����^UUUUUUUUUUUUUUUUUUU����         ����         ����^EUEUEUEUEUEUEUEUEUE����_UUUUUUUUUUUUUUUUUUU����      ����������@@@@@@p@@M����_UQUQUQUQUQUQu@@]����^UUUUUUUUUUUUu@@]����      t�<�����      �?��?�����^EUEUEUEUEUEUE'   �E����^UUUUUUUUUUUUU' T�U����       '@� ����@@@@@@@'PA�@����^UQUQUQUQUQUQU'TP�U����_UUUUUUUUUUUUU'T �U����      '   �����      '   �����_EUEUEUEUEUEUE�����E����^UUUUUUUUUUUUU_UUU�U����       ����? ����@@@@@@@@@@����^UQUQUQUQUQUQUQUQUQU����^UUUUUUUUUUUUUUUUUUU����         ����         ����^EUEUEUEUEUEUEUEUEUE����_UUUUUUUUUUUUUUUUUUU���� ��?        ����@qU�@@@@@@@@����_U]UUWQUQUQUQUQUQUQU����^UW�W]UUUUUUUUUUUUUU�����U\5       ������ p5       ����^�: �zUEUEUEUEUEUEUE����^�0 �pUUUUUUUUUUUUUU�����: �:       �����5 �u@@@@@@@����^�5 �uQUQUQUQUQUQUQU����_�5 �uUUUUUUUUUUUUUU�����5 �5       �����5 �5       ����_�: �zUEUEUEUEUEUEUE����^�0 �pUUUUUUUUUUUUUU�����: �:       �����5 �u@@@@@@@����^�5 �uQUQUQUQUQUQUQU����^�5 �uUUUUUUUUUUUUUU��������������������������?������������������������:������������������������:������������������������:������������������������:������������������������:������������������������?Q������������������������?������������������������:������������������������:������������������������:������������������������:�*                     �:�*                     �>�*                     ��*��������            ��*���<<����            ��* �<<��            ��* ��<<��            ��* ��<<��             ��* �<<��            ��* �<<��            ��*�?����            ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*                     ��*    �               ��*   ��|              ��*   ��_=  0          ��*   �UW=  0          ��*   �UU=  �          ��*   �UU=  �          ��*   �WU  0          ��*   �_�  0          ��*    ��              ��*    �?               ��*                    ��*                     ��*                     ��*                     ��*    ��              ��*    W_              ��*    _U              ��*    ��  0          ��*    l�  0          ��*    o�  �          ��*   ���?  �          ��*   ���>  0          ��*   �j�:  0          ��*   �j�:              ��*   �j�:              ��*   ����              ��*   ����             ��*   ���u             ��*   \5�U             ��*   �?��             ��*                     ��*                     ��*                     ��*                     ��*  ����           ��*  ����          ��*  <��           ��*  <��3�            ��*  ���3�          ��*  <��3�          ��*  <��3�           ��*  ?����           ��*                     ��*                     ��*                     �>�*                     �:������������������������:������������������������:������������������������:������������������������:������������������������?     ?� ��W�W� W�  [� �[�����������.頻�w���W������? �? ?� ��W�W� W�  [�  [� ����������������� �� ��  wU �� ?� ��W�W� W�  W�  W� ���������������������  W� �U� ��?      ?� ��W�W� W�  W� �W���������������j�ߪj�W���W��� � 03  03  ��  \�  \�  p5  �  �  �  �  �  �  �  �  �  �   �   �  �  k  k �o ��  <  �  �  �   <                    �  �  �  p  \  W5  �?  �:  �:  �:  �:  �?  W5  �:  W5  �             ��  pU? \U�\UU\UU5pUU5�VU:��� ��                     �*   �* ��* �"       �* �U� �U� �U� �i� �i� �Y� �U� �U�  �*  ?� ��W�W� W�  [� �[��������������쪪;�k��w��Wp����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         @ @      @ @  @ @      @@ @  @  @  @  @ U@U                        U@U @  @  @  @   @    @   @      @  @      @ @        @                                        @    @          UUUU @ @ @ @ @ @UUUU      UUUU      UUUU      @@ @@ @   P @  @ @    @@@@  �� �u]p�\�5�  �7  �?  �7  �?  �7  �7  �7  �?  �7  �7  �7  ����?  �������7|�7��7��7��7��7�������� �? � �  ����?�@��j�@�@�@�@��j�@�@�@�@��j�@�@�@�@UUUUUUUU�������������RUU�FUU�UU�VTU�VQU�VEU�V �V��V��V�VUUUUUUUU���_���^���^UU�^UU�^UU�^U�^UE�^UQ�^ T�^jT�^�T�^�T�^�T�^�V�V�V��V��V �VEU�VQU�VTU�UU�FUU�RUU������������UUUUUUUU�T�^�T�^�T�^jT�^ T�^UQ�^UE�^U�^UU�^UU�^UU�^���^���^���_UUUUUUUUUUUUUUUU������������UUUUUUUUUUUUUUUUUUUUUUUU    ��������                ��������    UUUUUUUUUUUUUUUUUUUUUUUU������������UUUUUUUU�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�V�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�T�^�����������������VUU�  ����������������                        ����������������UUUU    ����������������                        ���?������������UU��  �����������������?                        ����W@UPWUAWTSPCU@UUU�T�@ê^ ��z ���     �        ����U  UU@UTUUPUU      @�PU�zUU��UT�����<  �           ����U�AU@�PP�TT�UU�U@U�P?���� ��� ���@����  �           ����WUUUWUUUWUUUW���W���W���W���W���W���W���W  WUUUWUUUWUUU��������UUUUUUUUUUUU����������������������������    UUUUUUUUUUUU��������UUU�UUU�UUU���ժ�zժ�zժ�zժ�zժ�zժ�z�  @�UUU�UUU�UUU���������WUUUWUUUWUUUWUUUWUUU����WUUU����WUUU��������������������������UUUUUUUUUUUUUUUUUUUU����UUUU����UUUU����������������        ����UUU�UUU�UUU�UUU�UUUժ���UUUժ���UUU�����������������������?����ZUU�VUU�VUU�VUU�V��ռUU>���������������        �����������������ꀪVU��VU��VU��VU��VU��VU��WU��  �:  �  ����� ?� ��W�W� W�  [� �[��������������쪪;�k��w��Wp����     ?� ��W�W� W�  [� �[�����������.頻�w���W������? �? ?� ��W�W� W�  [�  [� ����������������� �� ��  wU �� ?� ��W�W� W�  W�  W� ���������������������  W� �U� ��?      ?� ��W�W� W�  W� �W���������������j�ߪj�W���W��� � ?� ��W�W� W�  [� �[����������>���޻�������ܫ�?W�� W  �   ?� ��W�W� W�  [� �[����������������ߪ�?���7 ��  p�  ��             ?� ��W3�W����0[��[��������������쪪;�k��?����W3�W����0 [� �[��������������쪪;�k��w��Wp���� 03  03  ��  \�  \�  p5  �  �  �  �  �  �  �  �  �  �                       �  p���_WUU���_  p�  �                 �  p  p  p  p  p  p  p  p  p  \  W5  W5  w7  �  �                 �  _  p���_UU�p���_  �                              �  \  k5  �:  �>  �   <   �   �      >   �   �       �   �  �  k  k �o ��  <  �  �  �   <                           /   �   �   �      <   �  ��  ��  \�  p5  �                           <   ?  �  �  <  ? �� p�  p�  p�  �:   ?   �  �  �  p  \  W5  �:  W5  �?  �:  �:  �:  �:  �?  W5  �  �  �  �  p  \  W5  �?  �:  �:  �:  �:  �?  W5  �:  W5  �                             ��\�_5�W� �?                                         ����WUU��W�? �?                             � �WWW�U\�� �U�<p����}��������?�w�:���03  �0                                 ���XU�<�����}��������?�w�:���03 �0     �? ?p����U_� WW5<�U����}w7�w7��w7������ 0� 3                                 ���<U%����}w7�w7��w7������ 0� 30                        �� `)X���  �� ��>� ��  03  ��  ��               � �X`	X`%� ���  J&  �� ��>� ��  03  �� 3                                   
��%h	 �� �/ ��� ��  �  3  3              
  �%��%`	 &X	 "V ��  � ��� ��  � �3   �                  <  ��? p��puupuu5pUU��uU= ���: |5 �W9 �U �U  �; ��  <  ��? p��puupuu5pUU��uU= �� �: �|5 W9 �U6 �U �U  �  �       <  ���Wwp]]\]]WUU|U]�W�  �0 \=� l�� �U? pU ��  ��  <  ���Wwp]]\]]WUU|U]�W�  �  \= l�0 �U3 pU pU ��  �?                  �  �� p� pi \Z5�\Z:̜�:?���5��uݜ�]ճ�^=���                 �  \:  ��� �����U?�����i���ii��iZ��i��0k�5���                  �  �Z �j pi3\�53��5���6\��6w]�6Wu�6|������?                 �  �5 3�� 3�� �UZ�ZZ�ji�iiץiW�i\�����                 �?  ��  � ����� ����� ��; ��: �� � �??   �  |=  {� ��� ��: ���������>������;� �?                                    �  _ �^; ���  ����� ��: �� ��� ��� ��� ��?�  |=  {�  �� ��> ��� �����������>? ��   �                    0  ��� �: ���?�������0ï��0�;��0��3�03� �      �   �� �:��� �� ���� �� ���;� �� ��00 0  �                            0��03030303030��                                    ��?��0��0� �0���0�0�0���?�                                    ��?� �0� �0���0� �0� �0� �0���?�                                ��?�0�0��0��0��0���0� �0� �?�            Q  ����   ����   ����       �      �      �   �      �      �            0      0      0 �     ��     ��     �0                       ������������������������0@  P  @  P  @  P 0 U  @   U  @   U  @ 0 T  U   T  U   T  U ������������������������pUUUUUUUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUUUUUUUpUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������������������������������������������������������������������                   ����                   ����                 ����                ����    @        ����                ����                ����                ���� @              ����                 ����                  @����                  ���� ������    ���������� p@@@@  p@@����p@@    p@@M���� p@@    p@@���� p�<�    p�<����� �?��?�    �?��?�����  '   � @   '   � ����  ' T�     ' T� ����  '@�      '@� ����'PA�     'PA� ����  'TP�     'TP� ����  'T �      'T � ����  '   �  @  '   � ����  '   �     '   � ����  �����      ����� ����  _UUU�      _UUU� ����  ����?      ����? ����                  ����                 ����                  ���� @                ����       @        @ ����                  ����                  ����N ��?              ���� pU�              ���� \UU              ���� W�W              �����U\5          ������ p5             �����: �:              �����0 �0     @        �����: �:              �����5 �5         @    �����5 �5             �����5 �5              �����5 �5             �����5 �5              �����: �:              �����0 �0             �����: �:             �����5 �5              �����5 �5              �����5 �5              ��������������������������?������������������������:������������������������:������������������������:������������������������:������������������������:������������������������?d�������������������������������������������������������������������������������������������������������������������������
                     ��
                     ��
                     ��
�?��??��?            ��
��<�<�?            ��
��<�<��          ��
��<�<��          ��
�?<�?�            ��
�<<?��          ��
�<<?��          ��
���??��            ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
    0               ��
   �=�              ��
   |�W            ��
   |�U            ��
   |UU  �           ��
   |UU  �           ��
   �U�            ��
   �W�            ��
   ��               ��
    �               ��
    �                ��
                     ��
                     ��
                     ��
    ?�               ��
   ��W              ��
   �W�              ��
    ��             ��
    [�             ��
   �[�  �           ��
   ���  �           ��
   �            ��
   ���            ��
   ���              ��
   ���              ��
   쪪;              ��
   �k��              ��
   w��              ��
   Wp�              ��
   ���              ��
                     ��
                     ��
                     ��
                     ��
  ��?����            ��
  ������� �         ��
  ������ �         ��
  �ÿ���?            ��
  ��?���� �         ��
  ������ �         ��
  �������            ��
 ��������            ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                   ��
                   ��
         �           ��
         �           ��
                   ��
                   ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     ��
                     �������������������������������������������������������������������������������������������������������������������������                                                                             ���  <��?�?<<   ��<  <�<��<��<<   ��<  <�<��<���<   ��<  <��������<   ��<  <�<��<��<?   ��<  <�<��<��<?   ���  ����< ?<<                                                                                                                                                                  �                 00                 �                                   �                 00                 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ���آ t ���d���� � �����������  ��� � �� � �� �ύ& ��"  7ĩ�� d
�� ��L`�       ^�n�~�������������������.�>�N�^�n�~®¾�����������.�>�N�^�n�~ÎÞ�                                                                                                                                                                                    �?����<�?<?� <�?  ��� ��?�� � <�� < ��?�� � ? < <� � ��3�<<�?����� < � < <� ��� �<<<���<�< ��� �  ?�����?<��?��<�<<�? �? ��00�?<?��?�����?�������?����<�< < <����?��<���������<��������� ������������ � ��3<<0 ?0<<���<0<0�?<0<0<0���������� � < < < <<<<<���<0<<�<<<���� � � � �������<<?�?�<�<<?��<0�0�3�??<?0��<<�<�<�<��<��?�������?� � ��?��<�<�<�<�<��?�?�����<��<�<����<�<���?�<��?�������������<0<0<0<0<0�<���<0<0�������<�<�<��?�?��?�<0���0<?���<0��������� � ?������                HZ�H�@��m��������8��HJJH

�zh8����m�� ����ɪ�8��i0��i ����h�zh`H�i0��i ��_�����8������h`H�H�H�H�H������ k�h�h�h�h�h`�H�Z�ڮڦڦ� ��8��JJ�8���� � ����� ����h�h�h�h�z�h(`Hڭ  �� �������%���h`��������?_ow{}~���������������������H�  ����h`�H�Z�ڦڦڦڦ�
��`���`�� �â �  q�- �� q�- ��� Ā��iɠ���iɠ������h�h�h�h�h�z�h(`Hڪ)�JJJJ Ŋ) ��h`HZ� ��$�#�0i��:8�0��A08�7�i �Ȁ�zh`�H����� L��Z�H�H�H�H�H�H�H��H��Hi�H�i �H ��8��JJ�8�����m��i ��������?������6� ��ȭ��h�h�� �������� ��m��i ���hh� h�h��0�� �����������ݬ�������
�h���h�	��h�h�h�h�h�h�h�zh(`�� �2��.HZ�Z�Z� ���������
������� �h�h�zh`�H�Z�H�H�H�H�H�H �à �ȍ���-�i��i �� � y�����m��i � ����h�h�h�h�h�h�z�h(`� �#��H���hH�Z�ڦڠ �������Lv�L�L~���� �Ȁ����LYȥH�H�Z�
�������������	8������	�� ��������*�e��i ��e��	i �	� �������	���8����	��������
�8����������������8h���h������
�������	��������h�h�z�h`ڦ
����	��.������`H�� �� h`�  � `H�Z�H�H� H�H�H�H�H�H�H�H�H �Ì�JJ�NN� ����:����:�ȱ���:����:��8�����h�Hڭɀ�
��8�
���Hȱ�����he��e������� ��h�+� � � qʍ �� �3� m������ q�ڮ� y�����
������P��r� m�����m ����8� � �8� �	� �m ��H q� y�h��,���� qʍ �� �� � q�ڢ ��� �� ������ �L.�h�h�h�h�h�h�h�h�h� h�h�(z�h`Z���z�`Hڦ��	���Q����h`�ڮڮڍZ�)���=%ˑȱ�=(ˑ8����Z�JJ�����

������	��
�M��z�

�����JJ����z��ȭ�h�h�h��h`?���H�Z�H�H�H�F�H� �

�ȱ�z��Z�H��hHڍ ǭm����m����hhh�h�h�h�z�h`��d % 4 O B 
 z  0 
7 p 
   � � ���7�kĺ���ŀŕ������vǀȗȦȭ�q�y�,�                                                                                                                          ����# X � �� �� ����Z � �� ��L�ͩ�Z � �� � %� � �� �� �� �� Qͩ2 2�L�̩����� �ũ2����� ��`H�Z�搭�������:�����:��� ���:������(z�h@�Ѝ&  ��h�
h�h�h��H(L}�H�Z�' )��c��� � 	��# �$ �% (z�hX@������`�����d����`�����
����L�ͥ��� ��L � � ��d����`����� � ��d����`�����	 � ��d�`����� � ��d����`���`����d�Lu���L���� �L���� �L���� �L���� 1�Lu�L�� NΜ�` NΩ����` NΩ������ ��������`d� NΜ�������� ������d�d�`�� �Ȝ������������������
��'䍖�'䍟� ��d�����
��i�������� �3䙺�3���������΅���������������d���`d��� �ȩ��������������d�d����� ������d�d�d�d�d�d��� �` �ȜH`� �	�H�G���H���ʽI�}�X�~�gH)�h)�JJJJ� �ۭ���JJ

��� ��h�Ƈ��л`څ{��| ܥ|�:



��` �` �� � (� �� 
� �� ��` n� "� �� �� �� �� ��`���"�������� �ݥ����  ������ ��`�H���� #�)��d� \� � ��L.� 0� (�����������
�������h�`��	��
��k�����
��cЅ�dЅ�b��kЍ �挩P 2�L��@���Ĉ� 24 68 :< >@ BD FH JL NP RT VX Z\ ^` bb`^\ZXVTRPNLJHFDB@><:8642����"��	�d��b���:
���Ѕ��Ѕ �`P�����&��H� �	���(��&х�'х �h�`���� v�`�H� �	���v�}IJJ

��X��� ��h�`��Hid��(�Hid� �ņ���vh�Xh�I`���d�L�ѩ������8����`���
d�L�ѩ���斜�`����d�`����`���d�`�����`���来��
�d���`����%枥��P�)�����
����L�d����`ڭ������������Wҍ�d��]҅����e�������i ���Ň�	���i��������`��d����`���L!ӭ��}���~��H)�h)�JJJJ��H ��h�����|i���i�������� ���]���}���~��H)�h)�JJJJ��H ��h�����.i�p�i�q����� �Ӑ��]  � Ҟ�����L!���Й`���L����L�ӭ��}���~��H)�h)�JJJJ��H ��h��i���i�������� ���[���}���~��H)�h)�JJJJ��H ��h�����,i�p�i�q����� �Ӑ��]  � c�ƥƥ��L����Л`H��e���p�$��8匐�p���e���q���8卐�q�8�h` �� 6� � �� ��`� ����
���
�L0Ԟ�����`��� gԭ�� �֭�� �֭�� �֭�� �֭�� �`�  rԢ  ��`ڽ�� ��	���� ���L�Ԟ��`��� #�)���ԝ�� � ��L�� _���`!#%� ��������������� �������������`ڢ ������]��͖���� ���
���������͟�0� ���
���������



%����L]Պi���� ��֍�L]���Ж #�)���֍��`ڢ ������T #�)�9��͖�����������͟0���������



%����L�Պi���� ��Ս�L����П #�)���Ս��`"!����- 4׽��%��������������� jڥ���������������`� ���K���F���A�g֝����������������� m֥���������������)�ƇL\�懥�����Ы`ڠ �������L�g�
���օh��օi g L�������`" !�־ֶ��ֲ��ֺ��� ��` ��` j�` +�` �� ��` �� ��` �� ��` �� ��`� rԢ ��``� R� 
�`� R� 
�`� R� 
�`� R� 
�`ڽ��"��������������� �� k�������`ڽ���������� �� kݥ����`ڽ���	����Lh׽�������� �� y�����$�����������L�ש����::���`��)�L� ���@���������� #�)�d�L�ש�����e�����������L�ש��L����ж`	ڭ��������	 � {����`����� 4�L3��� N�L3��� `�`��i����ʽJ؅]  �`�����ʽJ؅]  �`����������ʽJ؅]  �`�����������������
��:��L����
����L����
����L�ح�:��` �� � #�`���/����������)��敭�JJJJ��� �� yݥ����`�JJJJ�������8�0�
L"ٜ�`������������������"� m�L]��	 s�L]��L]�� �٥�����������`� ���`� �� |��`���	��0���`� �� ���`�����0���`� ���`��� +�L���� ��L���� j�L���� ��`��)��e�)��ň�挥�)���L�٥�)�e���`��)��8���ň�ƌƊ�8劅���)�e���L*ڥ�)�e���`��JJJJ��8劅�ň�ƍƊ�8�



����)e���Liڥ�



����)e���`��JJJJ��e�)��ň�捥�)��L�ڥ�



����)e���` ���d�d�� �p �ڭi�����L�ڥpi�p�qi �q�i�ɠ��L��`H�Z
��G��H�� �	 �z�h`�JJJJ����8�0	�
����`d�`��	� �H���h�L�� �ڥ��L�۽��}���~��H)�h)�JJJJ� ��ڭi��i� �ŎH�������I���X���g�����L�۩L�۩ 
����p���q��:
��p�ȱp� �h���	�L�`H��{��| ܥ|�:H�|�}8�|�&��"



m��~



m�h



��h���h`Hڢ �{�|��8�|���{�|�h`���� �ܥ�� :�`����B �ܥ��8��JJJJ��i��)ň����)��L�ܥ�



����)e���L�ܜ�`������)���������� �� k�`d���)�0.�������� �� kݥ��C��)����������L��'�������� �� kݥ����)���������`ڭ�����  ݥ�� �� ��`������)�?����d�Lj������� �� yݥ��!��)��JJJJ���Ljݭ��� �� y�`����d�`����`����d�`����`����	�&�����`d�`����d�`����`H�Z �⦔� ��pi�p�qi �q���pe��p�qi �q� �p��z�h`����������� �٥����������)��i��`�ɿ�%JJJJi8��L3��� �⥇��� �� ��`ڭ����� Nޥ�� �� ���`������)�?����d�L��:������ �� yݥ��!��)��JJJJ���L�ޭ��� �� y�`����������� �٥����������)��i��`���*JJJJ����8������� �⥇��� �� ��`ڭ����� ߥ�� ���`������)��p��:����)�0 ���� �� yݥ��Q��)�������Lm��0d�L�߭��� �� yݥ��)��)��������������� �� yݥ��
��������`�������� �ݥ������� �ݥ�����)���L�����)���`��)���� �߭���������� +ڥ����������)��i��`ڭ����� े� ���`������)��m��)�0&�������� �� yݥ��N��)�������Lpୟ������ �� yݥ��)��)��������������� �� yݥ��
��������`��)���� �߭���������� jڥ����������)��i��`������ƀ���Ɓ`�Hd� \ѥ����� 0� (�h�`�H \� �� �� �� � &� V� ��   ����� 0� (�h�`�P��d���� :
���Ѕ��Ѕ ǩg��g��� ��`�2��t���:
��s��t� �`h�p�x��������[��W��� ��`�[��w��� ��`�[��H��� ��`�H��<���� ����`� �	���(������� �`��  ������L����� �]  � � �� ���Z �L��������L�⭍��̭���
�	���� �׊���𳭍����	���� ݩ��Ld�	������� 4ފ	���� �ީ ��L��	���� �ߩ��L��`�)�����`d�`��
���p��q` �⩠��d�d��JJJJi
�� ��` ��8���d�d��JJJJ��ƕ�H� ��h�`�pe��p�qi �q� �p �ڥpi�p�qi �q�i�ɠ��`��e�m  e�m�e�`H�Z����� ���� ��z�h` �B���ƀ�J� � � � � � � � � � � � � � � � � � � � � �΁���R���ւ�Z���ރ � � �b����(�j����0�r�����8�z����������@���Ĉ�H���̉�h����.�p����6�x�����>����F���ʑ�N���Ғ��Ғ�V���ړP���Ԋ�X���܋�`����&�{�W�3������	
		""""""""""""""""""""$                  %$ +,-+,-+,-       %$             +-   %$               %$  +,-+,-+,-+,-   %$                  %$    +,-           %                  ####################!""""""""""""""""""""$%$())*%$(*%$(*%$())*(%$()*()))*$()*()*%% ####################!""""""""""""""""""""$%$./0%$./0%$./0%$./0%$./0%$0.//0%$.////0% ####################!""""""""""""""""""""$%$12313%$%$123123%$12312313%$123%$123%$123123% ####################!""""""""""""""""""""$%$444%$444444%$%$4444%$4444444%$44444%444% ####################!""""""""""""""""""""$%$555%$555555555%$555%$%$5555555%$55%$555555555% ####################!���&   ��ύ& `���&  ��ύ& `���&  ��ύ& `���&  	��ύ& `���&  ��ύ& `���&  ��ύ& `���&  ��ύ& `                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           L�L��L`�LI�L�L��� ��� �� ��� � � � � � � � �* dWd_� ���Xdc`�����;� ���4� �5�  D��;�;�6� R�����H� ���A� �B�  ���H�H�C� �����J������ ���� ��  ������-� ���&� �'�  ������ ���-�-�(� �c��� �� `�`���ȱ�ȱ�ȱ�ȱ�)
��=���=���)0�"ȱ����XȄdd �� �L��! l�� �
�� �d!��Ȅ!d���1�2�4ȱ2�5ȱ2�6ȱ2�7ȱ2�8)
��=��9�=��:�8)0�=ȱ2����XȄ1d;d<�6� �� �� �])��	���d> ��`�>�?�Aȱ?�Bȱ?�Cȱ?�Dȱ?�E)
��=��F�=��G�E)0�Jȱ?����XȄ>dHdI�C� к� �� �])��@Ы���d1 R򀠤#�$�&ȱ$�'ȱ$�(ȱ$�)ȱ$�*)
��=��+�=��,�*)0�0ȱ$����XȄ#d-d.�(� й�/ ��� �
�$� �d/��Ȅ/d#���Z
�����[����\�[�ȱ[�`�Z
�����[����\�[�$ȱ[�%`H�Z�)?	@�K�;��%K�K� ���)@��J��K�K�"�8��"��)0�"Ȅ ����� �d �K� z�h`H�Z�))?	@�K�);��%K�K�.�+��*)@��J��K�K�0�8��0��*)0�0Ȅ.�+����.�*d.�K� z�h`H�Z�7)?	@�K�7;��%K�K�<�9��8)@��J��K�K�=�8��=��8)0�=Ȅ<�9����<�8d<�K� z�h`H�Z�D)?	@�K�D;��%K�K�I�F��E)@��J��K�K�J�8��J��E)0�JȄI�F����I�EdI�K� z�h`� `� `H�Z�X����Y���X�_�Y)?
�����a轱��bd` %�z�h`d_�* dW`�`�a�Sȱa�Mȱa�Nȱa�T)
��=��P�=��Q�T)0�UȄ`dOdR�S� �dc`H�Z�_���L���M�V�S;�V)��V�R�P��T)@��J��V�V�U�8��U��T)0�UȄR�P����R�TdR�S)�K�Y)����
�@����K�K�V�( �K�W��* �W�O�O�N� %�z�h`H�Z�  l�  ��dd#��!�/ �� � �� �� �����z�h`H�Z�� ��� �d^�])?�^�D�� �>�^
��%��2�1��?�%��3�1��@d1d>� ���])����� ��]��� R� ��z�h` j�� j
�� w(�� j�� j
�� (�� j�� j
�� w�� �� �P�� ��� �
�� j(�� ��� �
�� �(�� ��� ��� ��� ��� �P��     � �(�� �(�� �(�� �(�� �(�� �(�� ��� ��� ��� ��� ��� �
�� �(�� ��� �
�� �(���� ��� �(�� �P��     � w�b� w(�b� �
�b� w
�b� �<�b� �
�b� �
�b�  �b� �(�b� �P�b� ��b�  �b� w�b� q�b� w�b�  �b� q(�b� d�b� q�b� w�b�     �  �b� ��b� ��b� ��b� ��b� ��b�  P�b�  P�b�  P�b�  P�b� d��E� q�b� d�b�  (�b� w�b� q�b�  (�b� ��b� ��b�     � w�b� ��b� ��b� ��b� ��b� ��b� ��b� ��b� w�b� ��b� ��b� ��b� ��b� ��b� ��b� ��b� ��b� ��b�  P�b�     � ��b� �(�b� ��b� �<�b� ��b�  �b� �(�b� ��b� �<�b� ��b�  �b� ��b� �(�b�  �b� ��b� ��b�     � ��b� �(�b�  �b� ��b� �(�b� d(�b�  P�b�  P�b�  P�b�  P�b� �(�D� �(�D� �(�D� �(�D� ��b� ��b�     �  (�b� ��b� ��b�  (�b� �(�b� �(�b� �(�b� ��b� ��b� �(�b� �(�b� �(�b� ��b� ��b� ��b� ��b� �(�b�  P�b�     � �P�D� P�b� wP�D� �P�b� �<�D� �b� w(�D� j(�b� w(�D� �b� w�b� �P�D� �
�b� �
�d� �
�b� �
�d� �(�D� �
�b� �
�b� �
�b� j
�b� �(�D�     �P�"� �P�"� �P�"�hP�"� �<�"� ��"� �(�"� �(�"� �(�"� �(�"� �(�"� ��"� ��"� ��"� ��"� �(�"� ��"� ��"� �(�"�     � ��� /��     � j��     � �� �~� w~� �}� �|� w|� �{� �z� wz� �y� �x� wx� �w� �v� wv� �u� �t� wt� �s� �r� wr� �q�     � Y��     � T�� Y�� d�� q�� �� ��� ��� ���     � d�� q�� �� ��� ��� ��� ��� ���     � ��� ��� ��� �� _�� K�� ?��     � ��� ��� �� _�� K�� ?�� /��     ���������	�,��f� �   �f� �I� �   �f� �I� �   �Y� �F� �6� �   �F� �l� �6� �h� �   �h� �h� �h� �f� �f� �   
	 �

		 �
	�	
 ��				


�
�

����	��!�{�  �  ���y�  ��W���  /�  ��  1�C�O�����Q�1�C�O������W�c�������������                                                                                                                                                                                                                                                                                                                                                                                                                                             �� �(�