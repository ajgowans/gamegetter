(�����������������������������������������                                   �? �                  �              000 �                  �              �? �                 �?             �� <  �                 �            � �    �                 �          � �?�?   �                ��         0 ���   �               ��<         � �����  �              ���         � ���  �              ���         <  ��? ��             ����            ���� �             ����          �  ����            �����          0  0����            ����?          <<��� �           ����         ���� �          ������         ��� �         ��?�����       �  <���  �         �??�����       0� �  ���  �        ����������       0� �   ?  �        ���������       03 3     �       0���������       03�� �0  �      �?���?��?��       �0�0 �0  �      �?�0�?����        0�� �0  �     ���  �?����        0���0  �     �? �  �?���<��        0�0     �    �� �  �?�����        0 3     �    ��  �  �?������        0 �  ��   �    ��  �  �?������        0  0    �  �?��  �  �? ?����        � �0    �  �?��  �  �?  ����        ���0 ?    � �����  �  �?  � ��        �<���    � �����  �  �? 0� ��          <�   ������  �  �? <� �           3���   ���� ��� 0� ��? ?� �           33? 0   ��� ��� ?� �������           �<� �?   ��� ����?� ��?����           0<3� �   ��� ����?� ������           00�  �   ��� ����� ������           0�  �   ��� ����� �� ���3           0��    ��� ���? � � ���           0    ��� ��� � ��?���           0 �  ��� ��� � ������           � ��   �������  ��?�����             0�   �������  �������               0�   �����?��  ���?����               0�   �����?��  �?�?��?��������������  ���������?��  ����?TUUUUUU��UUU � 0UUU�������    � ��       |  0 ?0   ����� ��   0� ��CUUUUUUU�O]UU1  �\UUU����? �� � <�  ��CUUUUUU��]UU���� �U���� �� � ?�  � ��������_����ª� �0����� �� ��?�  � ��������𮪪ʪ��?�����? ���?�?�  ��������� ����?�� 0�����? ������?���������T����?��� 0������ �������?�       �A��   ����? ����� ����� �����       \P�?    �0 0 ��������? �����       U�    ��� � ������� �����      �A��    �0 0    �������� �?��?      \P��     �� 0    �����?��  ���     �U�?      � �    ����?��?  ���     pA��          ����?��?  ���     P���?   �     �����0 �?  � ��    �U�� ��  0 0    ����� �?  0 ��     p@��𺫮   �   ��� � �?    �<     P����������   ��� �  �?    �<    �T�� ����><�3��   ��� <  �?    �     p@��?�����������   ���   �? <  ?     P�������������   ���    �? ? �?    �T��������        ���    �?�? �?    p@��? �?����:        ���    �?� �?    P�� ������        ��� �? �?� �   �T�� �����        ��� �� �?� �   ����   �����        �������?�  �  �Щ�? � �����       ��������? �  _ U�� �  �����       ��� ����� ?� �PU��  �  ����       ��?������ ��  \ TU�? �� �����       �������� �?  ���� ��������       �����?��  �?   ��� ��������       � �� �?��  �  @���   3  <����       ���? �?�?  � �T���     ����       ��� �?�?     �J���    �0����  ��  ��������?����� ������?  �����  pU  ���TU���?UUUUU @UUUUU  ��������� ������?  ���?     ��        �����TUU� pUU���?  ���?    � <       �0����   �U5  ���?UU���?U0PU}UU�UUUU  ���?   �U5  ���?UU���?0U�TUU�UUU � ��OUUU�UuUU���?UU���??T}UUUU��TUU �� ��SUUUŪzUU���?�����?
?�WUUUUU���*  ? ��TUUUŪzUU���?�����?�?fUUUPTY-���    �?����ʪ������?�����?�?_UUUUAU�����0     <������������?�����?��UU PUUu�����   �������������?�����?�cUPUUUTUZ���?   �������������?  ���?�cUUUUTQ=    0   �������������?  ���?�XUEUUWUTTU��?  �       ��  ���?  ���??DUPU��UQE_�    �    ��  ���?  ����?FQT� �PU�CU  �         ���?  �����QU  �0 U �3��2         ���?� �����U�    LP ��0 �         ���?� ����#AE1    p W �� ����        ���?�����cUQ    �W�V�_� ���        ���?0����XEQ     �Z�@5 ���        ���?p���?XE     ��j} � ���8        ���?p���?HA�       ��_T� ��8        ���?p���XQ�       ��[P�0 �<�        ���?� �?�VQ5       ��k@5����        ���?  �?�VQ5       ��U � <0�?       ���?  �?� RU1       ���VT� �0�       ���?  �?��UU1       ���ZP= �        ���?  �?<�UU        ��j@           ���?  �?�UU        ���U�            ���?  �?�UU        ���V1  �          ���?  � �ET   ��
 ��Z  0          ���?  � `EU   L� 0���   �         ���?  � `E   �X
 0 �;   W��        ���?  �0`QU  �? � 0 �  � UU������������?  �0hQT�   �  � �    PUUUUUUUUU���? ��<XQA5p       � �W           ���? ���XQE5p          �jU          ���? ���hQU5�           ��ZUU         ���? �� LkAE12          0����ZUUUUUUUUUU���? �� \�aE�       �  ������ZUUUUUUUUU���? �? |[aA�   <   O   �����������������? � �B�  �S �U   ������������������? �  �A0  0U1 ��   ��*����������������? ��  LA�@_E1�     �
���������������?���  \b�\�]T1     ����������������?��� U��0QT<       ��>��������������?�?pLZ��ST       ��3          ���?�?p\X�uTU�       ���          ���?�p�E%�E]T}       �>�          ���?�p�WdQU�       �          ������@WUUW\��?                 �����    UW@UDT�                 ����� ��?�U5UpUUU�     0  � 0       �����?@MA�TUM\EQ�     �  ��� <      � ����|1UUUWUE�QQ�     �  �����      <�����WUUUU_G_QUDU<       �����     �?�����TQUUUOUUUUUUU�       �����    0 ����WUUUQDQU�fVU�     �����     ����� UUUU��UT dUUU�     �����   �  ����? �U1�CU�UUAPUUTU  �� ����     �?���?� ? ��VQUaQUEYUUT� ���<       ������� <UUP /TQ$QE� ����?       0 �? ���� SUUUQ�TDUQU���?����       �� �����UU�_UU� W UUU������     �� �?  ��� �5�UU5\UU< cUU0 ������    � ��  ��� �5�Y�|TU 0E���������    0 �?   ��? �5 S5 pUU  OU ��������    0 <�   ��   <  �� * ��?    ���?    ���    ��           �                 <�<    ��                           ��<    ��                          �?<    ��            X                  ?    �            �                 ��    �                               �     �                                      �����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ������&�h�,����ԍ  U��.�p����6�x���������ĈƈȈʈ�N���]�҉�V���ڊ�^�⋠�f�$�ST$TIME$STAGE $GOOD LUCK$MIND THE TRAPS$ WHAT A PITY$  WATCH OUT$           $      $PAUSE$GAME OVER$CONTINUE$SELECT LEVEL$END$EASY$NORMAL$HARD$GAME OVER$HIGH SCORE $YOUR SCORE $C$   TRY AGAIN   $V���Y�^�e�����������ЀÀԀـ�������	�~�o����P���ԃ�X���܄�`� #     ������Ɓ́ԁہ���������!�,�7�@�I�T�_�j�w�������������Ȃт܂������ $ $ $ " " "           	 
 
 




   
   �?  �� ��������������������??���p��\��W5��W5  �       �?  �� ��������������������?��W�W�5�\�  \�  ��     �?  �� ����  �0�0��2���  ?���p��\��W5��W5  �       �?  �� ����  �0�0��2���  ��W�W�5�\�  \�  ��     �?  �� �?�� ����,��,�0 <�  �  �  �?  \�  W�  ��      �?  �� �?�� ��0��8��8�0 <�  ?� 7W�5_p5|�_=�\��     �?  �� ����� �?0�8�8�< �  � ��\��\p�|�_=p5p�?�     �?  �� ����� �?�,�,�< �  � � �  �?  W5  W�  ��      �� ���?�<0 0�3Î��������?�5 ��� ����?�����     �?  �� ����  �<0�8 ������0����W��\p5���?               �   �$  �  �  �   � @ �  �@  �   � @ �  �   �   �   �����        ���0  ��0ê�ó��γ��γ��ί������������?������     �� �    0� �� �� ������ó������?�:������ 00< ��� �� �    0� �� �� �������<�3σ�����?0���� 00< ��� �     � 0  ���        ?<    �?   �     ����    �    ??     ?     �   � <        ��     ?�  �     ?<��   �    ��   �:  �:  �:  �:  �:  �:  �:  �:  �:  �:  �:  �:  �:  �:  �:  �:                     ����    ����������������                     �:  �:  �:  �:  �: ��:  �: ��: ��: �� ��                      �:  �:  �:  �:  �:  ��� �*  ��� ���  �� ���                                        ��    ��: ��: ��: ��:  �:  �:  �:  �:  �:                      ���     �� ��� ��� ��� �:  �:  �:  �:  �:      �  0   �     �  �:  �:  �:  �:  �:  �:  �:  �:  �:  �:                     ����   ������������ ���                     �:  �:  �:  �:  �:  �:  �:  �:  �:  �:      �     �      �                     ���?  � ������ ���?��                      0  0  0  0  0  0  0  0  0  0  0  0  0  0  0  0                     ����                ����                     0  0  0  0  0 �0   0   0   0    ��                      0  0  0  0  0  ��              ���                                        ��      0   0   0 �0  0  0  0  0  0                      ���              �� 0  0  0  0  0  0  0  0  0  0  � ���                ��� 0  0  0  0                      ����     �     ����                         �  0   �     �  0  0  0  0  0  0  0  0  0  0                     ��
   �  �   �  � ���                     0  0  0  0  0  0  0  0  0  0      �  0   �  0   �     ? ��3 ��� ��� ��<��?�/�?|0�7 �����L�(?<.�?�������?@��  �   � �� 0�: ��� <<� � ����à���>3 ��<��0������ �  � �� ��<  �   <   �   ? �< �<� �<����?�?�?������?�����? �?  �� ��W�5\�?� ��  w� �7�p�|�v��_=�V�2�jç�?������  00��00  0 � ���� 0   ���      ��������    3���� �/����> 3.�VUU� ��  � ���?���� ��WU� ��W]� ��Wr�������<<�� 2 �3�� 2 �3�� ��?<��  ̻p� ��N�p�   |�p�   �/�     ����������WVYe�u�^�����z���U�UV٤[�Uժ�������e�դ[�Uժ�꤫���UV٤[� ������      �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              &   �          ��                       �<        ���                         ?         ��                        ��� �� ?   �?�?�?� �?� ����   �3���?���   ���?��� ?��������    �3��3��3�   � �? � 0�?������? �� �3<�3��3�   ��?� �?�?��������   �3�3��3�   ��?� ������������  ����3��3�   ��?��?�� ������������0�3��3��3�   �����0� �?��������� � �3��3��3�   ��� ��0��?�������? � �3��3��3�   ���� � ?��������  �0�3��3��3�   ��?� ���?��������  ������0�   ��?�<������������� ���??�?�   �?� ?��0��� ?���< ����� ����  ������?�?�  ��<�� (a                          �                                     ���                                    ��+                                    ����                                  ����                                  ������                                  ������                                 ������                                 ������                                 ����;                                � ����:                         ��    ������>                         |4    0������                        �@�   0 ������                        |TU   0 ������                         U�  �� ������                        ��_�  0� ������                       ���:  0� ������                       � P��:  �  �����                       |U��>    ������                      ��R���?    0����   ��    �������������? C�������   ?����   \U   UUUUUUUUUUUUUU  PUUUUU�   <�������, ���              ��     �   <���?UUU  \UU             �      �  0���?   `U   UUUUUUUUUUUUU_UU�_UUUU�   ����   `U   UUUUUUUUUUUU�UU��CUUU�  0����SUUUaU]UUUUUUUUUUUUUU_UUUUi=UUU�  00 ��TUUU��^UU������������UUUUUU����
 � �?UUUU��^UU�����������YUUUUV���*    �����������
�����������WUUUUPUe5��?     ����������
����������sUU  TEUU����� 0   ��������������������XTUUU������  �����������          XUAUUUAUT      �����������          VUQU�UUU<�  0  �     ��             QT��UTEQ�W5  �  �     ��             �QU� �oTU�P�   �                    `E�  �DE@�  ���                   `UA=    T �� � �2                   HPQ    \����3 ��/�                   XUT    �U�U�W=� ���                   VQ�      �V=P� � �"                  V�      ,�Z@5� � �+                  R1      ���W � < 0+                  VT5       ��VT? 0>                 �UT       ��ZP��� 0�?                 �UT       ��j@5� ��                 �TU       ���U �0 0��                 `UU       ���VT 0��                 `UU       ���Z�  � �                 `UU        ��j0  �  �                 `UU        ���U  0  �                 `U   � � 0���    �                 XQU   � * ��:   � �                 XQE  �� �  �  �U�?�                XTU  � �   �  <@U����������       ZU�    *  0 �    TUUUUUUUUU       VTP�       ��� �U                   ?VTQ�           �ZU                  'ZTU<           ��VU                 �ZPQ�          ����VUUUUUUUUUU       �fXQ,       �   ������VUUUUUUUUU       �VX#     ��    ���������������
       <�PE(  �T p�   �*��������������
        cP  LU �?   ��
�������������
     0  SPD8P�WQ<     ����������������     0  �X 2�pU�      ���������������     < GU25L      ��������������     � �V�u�U     �  �� �               VaAU�      �  �>0 �               |QIaQUE�      �  �0                \�YET��      �  ��                � �UUU�UW��      � �                  �_EU�PU<      �                 0��UMD\UUU3       ��       �?     PSDP=UUSWEQT0     0  ��?       0�     _LUU�UU|@TT3     0  �3��?      �    �UUUU�W��WTQ     �  ����?     ���    0UTUU�SUUUUUUU=     �  �����      �   �UUUUQTUE��U��    �  �����    � �    CUUUU�fU YUUU=     �����    < ��    |U��PDfUUTUU�   �? ����?     �    0� e�UTUXTUQVU�? ���       � ��     �  OUD�UITE0�����        �     0�TUDUT�<QUTUu������?      ���      ppUU�WUU0�@@UUU������?     �? �      ppUUWU�XUUL������?    �  ��       ppV� U�  DQ��0�����?    ��       p�T \U�  �SU �?�����?     �        � �  �??�
 ��   �����    �<<                 �%                 �                 ��                 �?                 �                 �                  �                  ��                  �                  ��                                    �?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ���آ t ���d���� � �����������  ��� � �� � �� �ߍ& ��"  �é�� d
�� e�L`�       ^�n�~�������������������.�>�N�^�n�~®¾�����������.�>�N�^�n�~ÎÞ�                                                                                                                                                                                    �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  HZ�@��mHJJH

�zh8����00�/��m�ɪ�����i0��i ����zh`H�H�H�H�H������ *�h�h�h�h�h`xH�Z�ڮڦڦ� ��8��JJ�8���� � ������i0��i ����h�h�h�h�z�h(`Hڭ  �� �������%���h`��������?_ow{}~���������������������H�  ����h`xH�Z�ڦڦڦڦ�
��`���`�� �â �  _�- �� _�- ����i0��i ����iɠ���iɠ������h�h�h�h�h�z�h(`Hڪ)�JJJJ �Ċ) ���h`HZ� ��$�#�0i��:8�0��A08�7�i ��Ȁ�zh`xH����L��Z�H�H�H�H�H�H�H��H��Hi�H�i �H ��8��JJ�8�����m��i ���ﭩ���I������@� ��ȭ��h�h�� ��������)�i0��i ��m��i ���hh� h�h��0�� �����������ݬ�������
�h���h�	��h�h�h�h�h�h�h�zh(`�� �2��.HZ�Z�Z� ���������
������� ��h�h�zh`xH�Z�H�H�H�H�H�H �à �ȍ���7�i��i �� � g�����m��i ��i0��i ����h�h�h�h�h�h�z�h(`� �#��H���hH�Z�ڦڠ �������L[�Ld�Lc���� eȀ����L>ȥH�H�Z�
�������������	8������	�� ��������*�e��i ��e��	i �	� �������	���8����	��������
�8����������������8h���h������
�������	��������h�h�z�h`ڦ
����	��.������`H�� �� h`�  � `H�Zx�H�H� H�H�H�H�H�H�H�H�H �Ì�JJ�NN� ����:����:�ȱ���:����:��8�����h�Hڭɀ�
��8�
���e�ȱ������e�������� ����+� � � _ʍ �� �3� m������ _�ڮ� g�����
������P��r� m�����m ����8� � �8� �	� �m ��H _� g�h��,���� _ʍ �� �� � _�ڢ ��� �� �������i0��i �L�h�h�h�h�h�h�h�h�h� h�h�(z�h`Z���z�`Hڦ��	���Q����h`�ڮڮڍZ�)���=ˑȱ�=ˑ8����Z�JJ�����

������	��
�M��z�

�����JJ����z��ȭ�h�h�h��h`?���H�Z�H�H�H�F�H� �

�ȱ�z��Z�H��hHڍ �ƭm����m����hhh�h�h�h�z�h`��H 4 Y B 
 �  0 7 z 
   � � ����*ă�����S�hŘŪ���[�e�|ȋȒ�_�g��                                                                                                                                                �������ύ& x�d�# ��Xd9 �� � J��ύ& x�d�# X �d9� r�d9 � � �� �  r� �����$d'dddddd nͭ��
 ��  r������� /�LLͭ�� �:�d: �ĭ���� � ��5�������d ذ  �� �ЀH���h �Ҝ��'� � �� �� �� ��L���$0L�� 0����L�� h���L��L��d<d=d9����������P�6���������6� r�d'dd!��" �� b� K� i� ѩ�( x� r� �ѩ0�&�d%���1 ��d)d* 	ѩ� ��� �� �Щ�9����`Hڢ � �P��E�� 	�F��.��������������-��������
����� �P�&��������E 	�F��0��/�P�h`H�Z�H�H�ȍ������
��i��ȹi��� ��#ȱ� �ȱ�+ȱ�5ȱ�7�8�B����ȱ��8���� ;������� ��i��i ��Ѡ��+ȱ�5ȱ�7�8����"�5�+� ��5� ��+�::�5�+� �ʆ+���� ���P��F���� �P����F��h�h�z�h`H�Z�(���. 	ѩE� ��� ���E����ڮ����� }π ��� �ͨ��Pz�h`Z���1 	ѩE� ��� ������
������D���:���;�Ө�P� �˘z`�Z���
� �蘤���	��� �� �>� ���	: �� �.� �� �8�
: �� ��� ��	�8�
 �� ���� z�`ZH��P� � �� ȹP� ��i
��P� ���P� �h� �hz`H�Z�+� �( 	ѩE� ��� ���E���
�訹P� ���P���z�h`HZ� ����� �	� � i�1 ���i�����zh`HZ 	ѥ#����� ������� 	ѩ� ���i��#���!��"�� �������!�"�� �!zh`H�  ee6m# e5e�h`H�Z� �� �� �	� d�P�1 �����F�2ȥ��
� �� ���m�� ��i ��ɭi���z�h`H�Z�H�H�H�H�������H���� hť 8� S�h�h�h�h�z�h`H�Z�H�H�l����� Sť Sť S�h�h�z�h`H�Z�5H�H�H�H�H�
����ȹ���d��� hť5 8� S�h�h�h�h�h�5z�h`�Z��d�)�
���8�
�e�؊JJJJ� ����i����إ��z�`H�Z�H�H�H�H�$������I��ȹI�� �Ơ���ȹ���i����� �	 ���i��$ ��h�h�h�h�z�h`H�Z�%��	� �, Ӏ'��	��� Ӏ�&��	� � Ӏ����� �z�h`H�Z������&�/�%�0��*�
�%�/�&�0d* c֥,� �a OԮ�)�*��8�
�)� �1�*�,��i
�)� ��*���:�)� ���*�
�)� �Ȅ* ��� �Lԥ*� �	�) ��� �V �֥&���8�(�&���e(�&��%��8�(�%�e(�% �֥%��&� ԭ��1� �	 �ե'�� "�z�h`Hڭ�)������8��i���	�������)
i���)���������h`H�Z�*� ��+��-�+�-�,��.�,�.�
��+::� ��e-�)�*�+� ��,��.� �� �i
�*��*�d*z�h`�Z�)���P� ���L����� L����	��'� L����	��'� L����=dd�� c�%�/�&�0 c֥,��.��(�������e(�(� �P��L�������t�*� �� �j�)��
� ������� �N�)8�
�2�)��� �=�):�2����	�.�)�2���#�)i
�2�2 ��� �����'�)� �P���� z�`HZ�H�H�H�H�����1��B��,8���
��8���@��ȹ@���.
����ȹ���8�
��I��ȹI���
�� ��ȹ �� ��h�h�h�h�zh`H�Zd'��2�P�2��
� ���� ���i ���� �����1 ��z�h`H���/� ���-��.���0� ���+��,h`H�Z�+H�,H�-H�.H�/H�0H� �	�%�/�&�0 c֩
��+::� ��e-� �ש��+� ������-� ��� �թ�; ��d;�,� �W�.� �r� �׭i� �թ�; ��d;�i��i
� �� �թ�; ��d;8���� �� �թ�; ��d;�>�.� �8�i�� �� �թ�; ��d;��i
� ���i� �թ�; ��d;h�0h�/h�.h�-h�,h�+z�h`HZ��H��H���%�������8���������� T������h��h��zh`H���������������
�P)����P�1h`H�Z��=�%�/�&�0 c֥,� �p�.�l�
��+::� ��e-�� �U�E�Q���L����� H�P)�ɀ�h�4hi�dd�P���Pd� �
�� c������  �P� ~������  �8d=z�h`H�P��� �o��� �g��� �_�� ����  �dd�� c� �P�1 !٠�;�����3� ����+�-��	�.��
��������dd ~詂��  ��h`H�
�� ������ ������ ��� ��h`H�Z��H��H�����P�/�R�0�N��\8���9i M�M��� 6ڎ�)����)�jjjj����)�jjjj���"�)���� �ِ�������������h��h��z�h`H�Z�����M��
� ������ �� �5��8�
���'����"��i
�����	� �����	����8z�h`� ������ �
�����`HZ� �P�-�����
���
���� ��zh`H�Z���L+ۭ��
� r������L+ۭ��>�������������{ R٭��V���������� �P��	��P��� R٭����7���� �� �ܩ���#���� �� �ܩ����	������P� T������ ��z�h`HZ�5H��5���6i �P� �P�� ~ۀ�� ~���F���5��� �P��F�� ѩ�' ��h�5zh`H�Z�H�H�+H�+�P���H��:H�P�1 %� �Մ�
� ���	��+  ��+���+  ��+��� �8�+�
�+  ��+i
�+���
�+i
�+  �h�+h�h�z�h`HZ�+�P���	������P�1 %� ��zh`H�H�H�+��
� ��



i ��



�h�h�h`H��8��� �߀B� � �߀9�� �݀0�� 	ހ'�� �ހ�� 4߀�� �߀�� 7݀ �ܥ;��@�dd c� ��h`H�H�H�1H�%��&����1 ��h�1h�h�h``H�����7��8J�7h`HZ�E�P	��Pz���� =���� ��� �������������h`HZ� �P	��Pz����#� �3�F�4�!e3�3�e4�4������������ ������
 �������h`Hڭ����� =����� ���X �S���� E�F ��A���� ��4 E�/����8�3�0�3�4� �4� ���������� ��� ��h`Hڭ����� =����� ���p �k����8�3��3�4� �4 w�Q 8�L���� 8�? w�:��*��� ��8�3�0�3�4� �4�����3i�3�4i �4�� ��� ��h`Hڭ����� =����� ���} �x��(�� ��k�38鐅3�4� �4 ���3i0�3�4i �4�L���� ��? ��:��*������3i��3�4i �4����8�3�0�3�4� �4�� ��� ��h`Hڭ����� =����� ���} �x��(��8�3��3�4� �4 ��^8�3鐅3�4� �4 ��L���� ��? ��:��*������3i��3�4i �4�����3i�3�4i �4�� ��� ��h`H���� =� ��h`H���� =� �h`H��� �	�� �߀ ���h`H� � �ِ�����h`H�Z���P Mਮ� 6ڎ�)����)�jjjj����)��z�h`�Z��H�H���"�/��&�8���
����ȹ���
���8�����z�`H�Z�3H�4H�� �6ڠ �3�����J�������)��)� �3�3i0�3�4i �4�ʀ�h�4h�3��J�#�����3i�3�4i �4�8�3��3�4� �4z�h`H�Z�� �6� �3)�3ȱ3)�3��� ��3i0�3�4i �4ʀ�8�3�0�3�4� �4ʀ�z�h`H�Z�3H�4H� �3)ϑ3 -�3)�3 -�� �3)�3ȱ3)��3 -����h�4h�3z�h`HZ�3H�4H� �3)�3ȱ3)��3 -� �3)�3 -� �3)ϑ3h�4h�3zh`HZ�3H�4H� �3)�3ȱ3)�3 -� �3)?�3ȱ3)�3 -��3)�3h�4h�3zh`H�Z�3H�4H� -�3)�3 -� �3)?�3ȱ3)�3 -� �3)�3ȱ3)�3h�4h�3z�h`H�Z�3H�4H� �3)?�3ȱ3)�3 -� �3)?�3ȱ3)��3 -� �3)?�3h�4h�3z�h`H�Z�3H�4H��3)�3 -�3)�3 -� �3)?�3ȱ3)�3 -�3)�3h�4h�3z�h`H�Z�3H�4H -� �3)?�3ȱ3)�3 -�3)�3 -�3)�3h�4h�3z�h`H�Z�3H�4H -� �3)?�3 -�3)?�3ȱ3)��3 -� �3)?�3ȱ3)�3h�4h�3z�h`H�3i0�3�4i �4h`HZ����
� ����� ��

e��i ���3�iF�4��� �
�х���$��
��� ����
�#����� ����e3�3�e4�4zh`HZ����� ����$�L�̤5�d5 ��dd�� c� �ш�� �� �ܠ� ����zh`H�Z�H�H� �P��M�%�IZ����  �dd�� ~� �ј� :�P��d1 �� �� �����1 �� �ܠ �������d1 ��z��EЧ �ܩ��h�h�z�h`H�Z�H�H�H�H �é0��2��
����ȹ�� hť 8� Sť'd'� �Ci
����ȹ��� ��R� hũ��x��
����ȹ�� hŢx ������a��,��Z��
����ȹ�� hŠ �ĭ� �7 ����,��Z��
����ȹ�� hŠ �ĭ� �	 �����Сh�h�h�h�z�h`H�Z�H�H�H�H��	
�� ��ȹ ����� ����� m���h�h�h�h�z�h`d9H�Z�H�H�H�H �Ģ �h����
����ȹ�� hŠ �� �ĭ� ������h����
����ȹ�� h�� �� �� �ĭ� ������h�h�h�h�z���9h`H� �	� ����� ���� �� ��r�����d���� �� �� ��������� �� �� �� �é��T� �� �橀��  �d ��:��h`�H�H�H�H��������� ��h�h�h�h�`Hک �2:������h`H��H��=��� R٭��������h��d=h`HZ�H�H�H�H�H �é,��2��
����ȹ�� hŭ��0�����0�����0������������d���K��
����ȹ�� hŭ� Sŭ� Sŭ� Sũ��\��
����ȹ�� hť Sť Sť S� �ĭ��� ��� ��h�h�h�h�h�zh`HZ�H�H�H�H���

�d������&  �Ʃύ&  �ĭ����� �� ��h�h�h�h�zh`H�Z�� �� y � �����z�h`H�Z�� 8�� � � ����ذdddz�h`Hک �F�eJf����h`Hک �*��������h`H�Z� r� �֠��) :�'����1�����1���3��1�� �� �����1H��'����� �1 �� ����h�1��ө  r�z�h`HZ��
� ������ ������ ���zh` �é8��<��	
����ȹ�� hũ8��L��

����ȹ�� h�d�<��,��
����ȹ�� �� �ĭ�����&�� �ĩ$ �ĩ<�d�� �ĩ$ �ĩL����� �� �ĥ�8������`HZ�H�H�H�H���2��
����ȹ�� hũ<��A��
����ȹ�� hũ<��P��
����ȹ�� hũ<��_��
����ȹ�� hŜ��A��2��
����ȹ�� �� �ĭ��� ����3�2��$ �ĭ�� �
���P�����
���_������A���� иh�h�h�h�zh`H�Z�H�H�H�H �é����� ��ȹ �� �Ʃ��>��� ��ȹ �� �� �ĭ���� �� ��h�h�h�h�z�h`�� �`H�  �����L���Z�9�>�'�:�6�6����5 �ѥ5�$����7�6��:�;��������=�	 uڀ�P�6�<�<�
�x�d�# X�z�h@�Ѝ&  ��h�
h�h�h��H(L}�H�Zd<�' )�&���������� � 	����'��<��P�# �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    L�L��L]�LF�L� �P�Q�R �� �� � � � � � � � �* d�d�� ����d�`�Q����y� ��r� �s�  A��y�y�t� O�R������ ��� ���  ��憥�Ł� ��P���J�Q����]� ��V� �W�  ��R����k� ��d� �e�  ���]�]�X� ���k�k�f� 
���� �� ]�`�S�T�VȱT�WȱT�XȱT�YȱT�Z)
�����[轉��\�Z)0�`ȱT�����ȄSd]d^�X� �L��_ i�� �
�T� �d_��Ȅ_dS���o�p�rȱp�sȱp�tȱp�uȱp�v)
�����w轉��x�v)0�{ȱp�����Ȅodydz�t� �� �Q� ��)��	���Rd| ��`�|�}�ȱ}��ȱ}��ȱ}��ȱ}��)
������轉�����)0��ȱ}�����Ȅ|d�d���� к� �R� ��)��@Ы���Qdo O񀠤a�b�dȱb�eȱb�fȱb�gȱb�h)
�����i轉��j�h)0�nȱb�����Ȅadkdl�f� й�m ��� �
�b� �dm��Ȅmda����
��=����=������Tȱ��U`��
��E����E������bȱ��c`H�Z�Y)?	@���Y;��%����^�[��Z)@��J������`�8��`��Z)0�`Ȅ^�[����^�Zd^��� z�h`H�Z�g)?	@���g;��%����l�i��h)@��J������n�8��n��h)0�nȄl�i����l�hdl��� z�h`H�Z�u)?	@���u;��%����z�w��v)@��J������{�8��{��v)0�{Ȅz�w����z�vdz��� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ƈ��d���� z�h`� `� `H�Z���������������)?
������轥���d� "�z�h`d��* d�`������ȱ���ȱ���ȱ���)
������轉�����)0��Ȅ�d�d���� �d�`H�Z�����L��������;��)����������)@��J��������8������)0��Ȅ������Ɛ��d���)����)����
�@����������( ��ŕ��* ��捥�Ō� "�z�h`H�Z�  i�  ��dSda��_�m �� 
� �� �� ����Pz�h`H�Z�Q� ��R� �d���)?Ŝ�D�� �>��
��y��p����}�y��q����~dod|� �Q�R��)�����R �����Q O� ��z�h` F�� _#�� _#�� _F�!� _F�!� F�� T#�� T#�� TF�!� TF�!� G#�� K#�� T#�� _#�� T��3� F�� K#�� K#�� KF�!� KF�!� F�� T#�� T#��     � TF�!� TF�!� _#�� d#�� q#�� d#�� _��3� F�� ?#�� ?#�� ?F�!� ?F�!� F�� G#�� G#�� GF�!� GF�!� KF�� TF�� _��3�     � �F�!� F�!� F�!� F�!� �F�!� F�!� F�!� F�!� �F�!� F�!� F�!� F�!� �F�!� F�!� F�!� F�!� �F�!� qF�!�     � qF�!� qF�!� �F�!� F�!� F�!� F�!� �F�!� F�!� F�!� F�!� �F�!� F�!� F�!� F�!� qF�!� F�!� F�!� F�!�     � ?#�� K#�� T#�� _#�� ?#�� K#�� 8#�� ?#�� /#�!� 8#�!� ?#�!� G#�!� /#�!� 8#�!� *#�!� /#�!�     � ?#�� K#�� T#�� _#�� ?#�� K#�� 8#�� ?#�� /#�!� 8#�!� ?#�!� G#�!� /#�!� 8#�!� *#�!� /#�!�     � K#�� _#�� d#�� q#�� K#�� _#�� G#�� K#�� 8#�� G#�� K#�� T#�� 8#�� G#�� 2#�� 8#��     � K#�!� _#�!� d#�!� q#�!� K#�!� _#�!� G#�!� K#�!� 8#�!� G#�!� K#�!� T#�!� 8#�!� G#�!� 2#�!� 8#�!�     � 8�� ?�� 8�� ?�� 8�� ?�� 8�� ?ȧ� T�� ?�� 8�� ?�� T�� ?�� 8�� ?�� T�� ?�� 8�� ?�� T<�� ?<�� 8<�� ?<�� _�� T�� _���     � ?<�� G�� ?�� 8<�� /<�� ?�� 8�� ?�� G�� Kx�� T<�� ?<�� q<�� <�� _�� T�� _<��     � ?#��� GF�� K#��� TF�� _#��� dF�� q#��� F�� d#��� _F��     � �#�3�  F�!� �#�3�  F�!� �#�3�  F�!�T#�3�  F�!�#�3� �F�3�     � ��!� �!��!� ��!�.�!� ��!�T�!� ��!�}�!� ��!�     �     � �
�� /d��     � '
�� %
�� *��     � ,
�� *��     � ?�� 8�� ?�� ��� ��� ��� ��� ��	� ��
� ���     �     �	
�
	�
	
�
�
�	

	�	

	�	

	�	���

		�
	�M�Y�e�q�S�_�k�u�x��  ����  j���  6���  ���  ���  �  X�  ������������`�f�u��������������������2����������� % O  % O     % o  %                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    x� ���