~����.���N�ދn��������>�Ζ^���������)�;�M�_���á��'�Y������!�S�������M����������ˤ܀�����,�<�L�y�����7�?�?�����y�y�����7�7�7�7���?���ÜK�R�\�d�p���=�ۤ��K�=�|�O���ȁ+�ށ��́W���۟���۟���G���˝�G���˝�q���q���q���q���O���O���O���O���_���_���_���_���Ӟ�Ӟ�Ӟ�Ӟ�������������������STAGE  $YOUR SCORE $HIGH SCORE $CONTINUE $END $         OK                               LET US PLAY AGAIN $TIME$    PRESS START $$$
$

$$$$$
$$$$$$$$
$$$$$$$$$$#
$$$$$$$$$$$$$$$$$$$$$$$!$$$$$$$$
$$$$$$$$$$$$
$$$$$$$                    ffffffffffffffffffff`                  `                  `                  `       V          `       V          `       V          `       V          `       V          `       V          `       V          `       V          `       V          `       V       UUUV`       V       U  `   4   3       U  `   3   D    P U  `  4  "4Q U  ffffffffffffffffffff                    ffffffffffffffffffff`                 `                 `                `                a$%           `                 `                 `                 `                6`            5  U#6`           U  SE26`         D3"3#C`         44#D4#V`     E"  DE4#D3`     RU"fU$!""""F`     QU"4U1""""`    "U"D31""""ffffffffffffffffffff                    ffffffffffffffffffff`                  `                  `              ` `              ` `                 `   DDA         `                e                `       f        `                `                `   fffff  P    `   UUUUUP        `                  `                  `                  `                  ffffffffffffffffffff                    ffffffffffffffffffff`                  `                  `              P   `                 `  "            `  3        UP  `               `               `        U       `        U       `               `               `      3        # a%      3          `                  `                  `                  ffffffffffffffffffff          P        ffffffffffffffffffff`         P       `         P       `UUUU3fff`      `                 `                `              0  `   f              `   f             `   f             `   f             `   f  UU        `   f         1   `   f           `   f         0  `   f            `   f         `  `   f         `   ffffffffffffffffffff                    ffffffffffffffffffff` `       P        ` `       P        e `       `        ` UUUUUU        ` P     P       ` P     P          `       P f        `       P f        `       P UUUUU    `       P P        `        P      `       0 P     `        P    V `       P    V! `              V! `           $  f `             f ffffffffffffffffffff                    ffffffffffffffffffff`                 `                 `             UV`   UQ      ` `  U UPU   R ` `  U UP       ` ` UUUUU      ` `             ` `             ` `             ` `         b@ ` `            ` `             ` ` 0            ` ` `$$$$$$    !  ` ` `          !  ` ` `             ffffffffffffffffffff                    ffffffffffffffffffff`        P        `       UUUP       `        P     U ` U$UQ#AUUQUUUUP ` P      P       ` P      P       aP     P      `        P   "  `             "` `              "` eUUUUUUUUUUUU"Dfff `                 `                 a ffffffffffffe  `                  `                  `                  ffffffffffffffffffff                    ffffffffffffffffffff`                ` P              `                ` P              `              `aP         P @   `                `      P      UUPV`      0    Q      `      `          ` U               `      `     P    `    e`    P    `    `          `` U               `    P            `                 ffffffffffffffffffff                    ffffffffffffffffffff`                 `      P           `         QUUP   `       P      P   ` E      @   P   `      P `   P   `        ` U P   `        P`   P   `       `   P   `       UUUUP U `UUUUV             `  UUV             `               @  `        @         `           P      `                  `                  ffffffffffffffffffff                    ffffffffffffffffffff`        P    P    `        `         `        0    `    `            `             ` U    $  f    ` U   $$EUUUUC1  `                  `               0 `                  `                  `                  `                  `   f  f           `                  `                  `                  ffffffffffffffffffff                    ffffffffffffffffffff`                  `                  `                  eUUUU$%UUUU$%UUUUUUV`   e        P     `   f        P     `   e        P    `   f        P     `            P    `        $$  P     `       $%  P     `       P   P     `    UUUP UfP     `       P   P     `                  `                  `                  ffffffffffffffffffff                    ffffffffffffffffffff`             P    `                `       RBEUUQ  V`       P    P    `       P    P    `       P    P   `        P    P    `             P    `       @   `    `          !    `       @       `       @       `       %UUUUP    `  $    @         `                 `       `         `       `         ffffffffffffffffffff                    ffffffffffffffffffff`                  `                  `       ff         `              `     UUP       `         P       ` UUUUU    UUUUUUU ` P               ` P               `                 `                `                ` P U          U  ` P              `                  `                  `                  ffffffffffffffffffff                    ffffffffffffffffffff`         0        `                 eUUUUUUUU 0      U `            U `        `P    U `        `P    U `UUUUUUP `P    U `      P`P    U `    P  P`P    U `      P `P    U `      P `P    U `   P  UP `P    U `   P  UP `P    U ` UP   R"`3$  U ` U  UP     U `                 `                 ffffffffffffffffffff                ���R�R�R�R�R�����r�r����Ƽ������V��f�f�f������r�r����Ƽ������j�Z�V��������Z�ڦ�fڦ�Z��� �* �V�`UU	XUE%XU%VU�VU�VU�VUU�VUU�VUU�XUU%XUU%`UU	�V� �*      �
  Z� �UU`UQ	`UA	XUA%XUE$XUU$XUU$`UU	`UU	�UU Z�  �
     0�� �U�p��p�p_� �W� �U�U�  �?  W�  w�  w�  ;�  ��  �� ��    0�� �U�p��p�p_� �W� �U�U�  �?  w�  ��  �� ��������     ���_U��W�W� s� s��pU WU ��  ��  7�  �� �������?� ���_U��W�W� s� s��pU WU ��  W�  ��  ��  ��  �� ��� ���  ����W=����UU�5\�5\�u]�UU �� ��pUU�UU3���?������� ����W=����UU�5\�5\�u]?�UU3\��5p��UU�UU������:�:��? �� �_ W� w� ��  w�  W�  �� ��_�]u�����: {�  ��  ;� �?���? ��� ��� �W�  ��  W�  W� ����s�_��_�? �:  �:  {�  �� �?�    �   �  �  �5  ��  �U �U �U5 �U� �UU����   �   �   �   �                                   �   0  �  ��0��<?�����                                       � � �3����� ��� �?                                   �  �  �?����?���<���? ?�                                     ?  �� ?�������?������ ��?           �   (   *   . ��
���+��ϯ��������ÿ������+�������� �   �   �   *  .* �..���
���
���>��
:��+8��/���/���+���
����     �
  
� �   � 0�� 3� 3� ��  0 ��   
�  �
     �"���" � �(("� ��#��0"0�"0��0��#�� �((" � ��"�"���� �� ��0�? 0���: �����  ��  �  �  � �� � �  �     ��� �� ��0�? 0���: ��� � ���  �  �  ��  <�  <�  ?   �� ���� ���� ����� �� ��  �  �  ��  �� �� �� �      �� ���� ���� ����� ��  �� �  �  �?  �<  <   �         UUUUPPii��UUUUUT�VUUZ�Z�UU�ZUiUUjU�UUUUU�e�eUUUUUUUU    UUUUA�Vj�P@AAZUUZUijUUUU�iUiUUjUUUU�Z�VUUUUUU��f�UUUUUUUU    ��W���          �?{��?      � pppp������pppp�     �    �      00��00   ����W=����UU�5\�5\�u]�UU��� S�|UUpUU3���?�������      W  �    �    �    �    �    d %     4  4  D  D  W " �    �    d % 4  4  4  4  4  '  ' 
   %  d ! 4  4  4  4  4      '  T   d  4 
 4 
 D  D  D  D   
   '  d  4  4  4  4        ' $ �    d  '    '  '  D  D   
   4 	 d $ '   ' %
 &  '   
       D !
 d  4 
 4  4         '  & #   d # 4 
 4 
 4 	
 4 	 4 	 4 	       d  '  $  '  '      4  4    d       %   4 
 4  4  D  D  d % 4  4  D  D  ' 

 ' 
        d % ' 
 ' %
 '  &   
  %
       d           %    4  4  '  d                         %                                      ��                  ��              �                 �?             ��                 < 0             �                    �             �                     �             0    �?0��  �     �0 �  �?  ? 0    ��0�?�?  �?     �0 0  �� �? 0     ��� � �     �� <    ?  0     0 � � 0 �     ��       0 �  0 � � ���     �   ��   0    0 � � ���     �   ��   �    0 � � 0       �  �       �    0 � � � 0     �  �       ��  0 � � � �    < <  �   �    �  <�0 � � �<    �   0   <�    ��  ��0 � �  �    ��  0   ��    "\� � � � � � � � "*08CUh|�����$/?Qct���������!=Zw����6Y|���+Nq����)Lo����Ad����4Wz���	'	�� ��?  �W�  ��UU  �pUU5  �pUU�  ��WUU  ���UU  ����W  ��� ��  �� �U  �� ��  ���  �  ���0  ���0  �0��?  �@UU  ��U��> �TU�  �<_i�� �PU�  �PUU  ��j�V �PU�  �TUU  � ��V5 �TU�  U� � ��Z5 �TU� �@U� � ��~5 �PU� �@U� � ��� U� U�  � ��  ������  �p���>  �p���  �p ��  �TU	 �p ��:  �PUU �p ��  �PUU �0 ���  U� �0 ���  �0 ��?  ��  ��  ����  �\U�  �WU�5  ��U��  �pU�  �_U�=  ��U��  �pUU����� ������ZUU  �\U��  XTQE	 �� `UU  ��WU������XTQE������VU�  �pU������" ������*XUU  �\UE������bEUT�������UU  �WUP�������EU�������
VU5  ��U ������� ���������XU�  �\U������*VQE%�������HUU  �WU������*VQE%�������UU5  ��UU  �������  ��������b@U�  �pU�RQ�������HU������
�b�VU  �_U	RQ�������bU��������bXU�  ��UU �������"  ��������"��UU  �pU�(��������Q���������b�
VU  �\U!*��������Q���������b��hU5 � �W$* �������* �������"���U� � pU *RQ�������*%�������b��*VU � \U�%*RQ���������������b��*BU5 � W� &* ���������������"��*�Z� ��U	*&*����������������b��*&`U�p��*"*�������
��������b��*"�U�\%�*&* ������������"�
(&*V5�\��*&*RQ������������b��&�X5�W�� &*RQ������������X��)"�bՍW�
� * ����������
*���$��Ս��E!*�����������*F��Q$�*֏��E!*���������������*F��  ��ȏ��  * ������"��*���������%
�آ�(R%*RQ������������������X��%��آ�(R%*RQ������"���"�������X�
� ��Ȣ�(  * ������b���X�����
�"��
&��آ'*FQ$*������b���X�������b��*&��آ'�EQ$*������" �*�������b��*"��Ȣ#�   * ������b����������"��*&��آ'�E!*RQ������bT�b�������b�
(&
�آ'�E!*RQ������" �" �������b��"��آ#�   * ������bE	XT�������"���%�*¢'�Q%*������bE�VT�������b��%�*֏'�Q%*������" ��������b��  
�آ#�   * ������bTQE�������"��E!��Ȣ'*F�%*��������bTQE�������b��j!��؏'*F&*  ������" ��������b�
� ��؅#��("��������bEUT�������"��*&��ȅ'�*&��������bEUT�����
�b��*&��؅���*&��������" ��������b��*&��؅���*"��������bTQE�������"��*"��ȅ���$��������bTQE�������X��*&��؅	 h$ �� ��    � �� �V  &�؅�����������jEUT�����������ʅGQEQ	T�QEUTQE�QEQ�(+  �                                     � <                                     ��  ��� �� ��������� ��3������  �� ���<�0 0��� � � 0 <� 0� �  �� � ��� <�0 0��� <� �0 <� 0� <�  �� � ��� ��0 0��� <�0�0 0� 0� <�0 0�  0 ��� �?0  � � �0 ��  � 0� �0  0�  0 ��� �<0  � � �0 �� � 0� �0  0�  0 ���� ��0  � ���? ��� 0���?  0�  0 ��� ��0  � �� �0  �� 0�� �0  0�  0 ��� ��3  � ���0 ?  <� 0���0  �� � ��� � ?  � ��� �?0 <� 0���  �� 0 ��� < ?  � � ?� <0 <� � ?�   �0 ���? <  � � ?� � �0 � � ?�   ��  ��� �� 0  ��<���������<��  � <                                      �                                                                                                                                                                                                                                                                                                                         ��           �   �  �     �? �?�� <            �   �  �     � �0                   �  �   � � �� <                  �  �     ��� <   ����?��� <<�� �    ��    <<� ��������?� �     ��    ��� ?0����� �     ���   ��� <0� ���� �     <�<�<    ��� �� ���� �     �� ���   ��� �� ����� �     � �0 0  ��� �� �0� �� �     ?� ?�0 0 < ��� �� �0  �� ��    ?� ?���? �� �?��? � �? �?���?��?  ���? �?0�      �  �      0�?                         � �0      0 0                         � �      �                          �? �      ��                                                                                                   ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���آ t ���d���� � �����������  ��� � �� � �� �ύ& ��"  7ĩ�� d
�� ��L`�       ^�n�~�������������������.�>�N�^�n�~®¾�����������.�>�N�^�n�~ÎÞ�                                                                                                                                                                                    �<<<?�<<<<<�  �������?  �<< <�< < �?  �<< <� <<<�   �0<�?    �?< < � <<<�  �<<< �<<<<�  �?<<<< ���  �<<<<�<<<<�  �<<<<�? <<<�  �0<<<<�?<<<<  �<<<<�<<<<�  �<<<<< <<<<�  �<<<<<<<<<<�  �?< < �< < �?  �?< < �< < <   �<<< <?<<<<�?  <<<<<<�?<<<<<<  �������   ?   <<�  <<� � <<<0  < < < < < < �?  0<<�?<<<<<<<<  <<<�<<?<<<<<<  �<<<<<<<<<<�  �<<<<�< < <   �<<<<<<<?<<�?  �<<<<�<<<<<  �<<< � <<<�  �?������  <<<<<<<<<<<<�  <<<<<0�   <0<4<3<3<3<3�  <<<<0�0<<<<  <<<<�����  �?<<  � <<�?                  HZ�H�@��m��������8��HJJH

�zh8����m�� ����ɪ�8��i0��i ����h�zh`H�i0��i ��_�����8������h`H�H�H�H�H������ k�h�h�h�h�h`�H�Z�ڮڦڦ� ��8��JJ�8���� � ����� ����h�h�h�h�z�h(`Hڭ  �� �������%���h`����������ow{}~���������������������H�  ����h`H�Z�ڦڦڦڮ	�
��`���a�� �Ü	� �  q�-  y���� �����iɠ���iɠ������h�	h�h�h�h�z�h(`   Hڪ)�JJJJ Ŋ) ��h`HZ� ��$�#�0i��:8�0��A08�7�i �Ȁ�zh`�H����� L��Z�H�H�H�H�H�H�H��H��Hi�H�i �H ��8��JJ�8�����m��i ��������?������6� ��ȭ��h�h�� �������� ��m��i ���hh� h�h��0�� �����������ݬ�������
�h���h�	��h�h�h�h�h�h�h�zh(`�� �2��.HZ�Z�Z� ���������
������� �h�h�zh`�H�Z�H�H�H�H�H�H �à �ȍ���-�i��i �� � y�����m��i � ����h�h�h�h�h�h�z�h(`� �#��H���hH�Z�ڦڠ �������Lv�L�L~���� �Ȁ����LYȥH�H�Z�
�������������	8������	�� ��������*�e��i ��e��	i �	� �������	���8����	��������
�8����������������8h���h������
�������	��������h�h�z�h`ڦ
����	��.������`H�� �� h`�  � `H�Z�H�H� H�H�H�H�H�H�H�H�H �Ì�JJ�NN� ����:����:�ȱ���:����:��8�����h�Hڭɀ�
��8�
���Hȱ�����he��e������� ��h�+� � � qʍ �� �3� m������ q�ڮ� y�����
������P��r� m�����m ����8� � �8� �	� �m ��H q� y�h��,���� qʍ �� �� � q�ڢ ��� �� ������ �L.�h�h�h�h�h�h�h�h�h� h�h�(z�h`Z���z�`Hڦ��	���Q����h`�ڮڮڍZ�)���=%ˑȱ�=(ˑ8����Z�JJ�����

������	��
�M��z�

�����JJ����z��ȭ�h�h�h��h`?���H�Z�H�H�H�F�H� �

�ȱ�z��Z�H��hHڍ ǭm����m����hhh�h�h�h�z�h`��d % 4 O B 
 z  0 
7 p 
   � � ���7�kĺ���ŀŕ������vǀȗȦȭ�q�y�,�                                                                                                                          �	L��Ln�L��x�d�# X � ��)��& ��� �X� �� �d � � �ĩύ& ���d!��H��������������d���$��  �d$  ��H� 갷�ǭ��� ����!�� �� �ϥ�
�	�����˭��
 �ĭ���d�
�C���� j� �πF�� �� �π:�� �� �π.�� �� �π"��L�� �� �π
��L��~ͅ�ͅ   �ϥ�	��L�̜�i�jφϊϊϔϘϜϜ�H�  ����h`H�H�H�	Hd��� ����  �8��i�i�� ��ک �	�#΅�$΅ � �ͩ *׭  ��� �ͩ �	h �� v������  �h�	h�h�� *�d���d h(`%������������������������������������������������������������������������������������������������������������������� �
���� ��������������������������������� �����
� ������� ���*��������������������������� �������������������������������������������������������������������������������������������������������������������`Hڥ�����  ��� 	�����h` �` � � �` �` �`H����d����  �h`H�� $� '� �ϥ��	 $� '� �h`H��� !� � � �d�	��� �h`H�  ��Lx̩����������� �����=������� � !� ��h@�Ѝ&  ��h�
h�h�h��H(L}�H�Z�' )� 	�P�# �$ �% (z�hX@Hd 7ĩ��<�� � ǩ *ש��h`Hڢ �:��:��
���h`H�Z�H�H������d!d"��H  ׭H��M�  ��F U� �ϥ��	��
���ݭ�
�
 �ĭ�
��d
��L��~ͅ�ͅ   �ϥ�
����h�h�z�h`				!�HZ�"�Sх�Tх���"�"�2�d"zh` �� 4�����HZ�Hd���y��)�
��"��1�h��:���������6�����-�������������������������� ҭ����Й���������h�zh` �Ҁ�  ө������H�Z�H�H��H��H 3׭������ 6׭��
�H�iȅ�i �h8�
��

m�

m�� �ұ���)�JJJJ�)��h��h��h�h�z�h`He�� e���h`HZ�H� �������



H�)�h��)�������� -׭����	H� �	�� 0�h�	h�zh`HZ�H� ����)��)����� -׭����	H� �	�  0�h�	h�zh`H���������  � [�h`H� � ץ�����D)����d�2 $� ������	 $� �������� 1� >������ 1� Z����� ��h`H�Z Wװ*���F����F�� <������ T� <׈��z�h`H�Z Nװ,�ɠ��F�	���F�'� 9������ E� 9׈��z�h`H�
��y�JJ�h`H�
��y�J�h`H�Z Hא���
�G�� ?�z�h`H� Kװ Qאdd�
�G�� B��h`�Z��d�)�
���8�
�e�؊JJJJ� ����i����إ��z�`H������ Z�h`H�H�H�H�H�H�H�	H�H� �	 ;� P�h�h�	h�h�h�h�h�h�h`Hڜ��� 0��i�����h`H�(�� �� j� ��h`H��H��H�����<�� 6שP��� �ũ`�� j� ǩh��� �� ��h��h��h`H�Z�H�H�� ���� j� �H�H����  � ŭ  ��'� *��������i��i �hi�h���hh�
 *�h�h�z�h`H�Z�H�H���2����i�� A���	�e���h�h�z�h`H�Z��)�2�����*�����"����������
�����������z�h`                                                                                                                               L`�L��L�L��L,�L�LN�LF�L�L��L7�L`�LZ�L#�L��L��Li�L
�L��Ld�L��L��Lb�L��L��L
�L��L��L�L��L��L�H�Hd ddd�=���!���������x��Z������� �� �� � W� z� 	� ��

e� ���
����dh�h`H�Z�H�H��:
�� ����� 
٢ � �������i��i ��i��i �����h�h�z�h`H�Z 7Ĝ���� �� �حi������z�h`Hڮ�H)�JJJJ i��i�h) i�h��h`Hڦڦ�
��(���)�� �h�h��h`H�Z�H� �	� 
٭������ �٢ ����� �؀� C� ������h�z�h`Z��H��)



��ȱ)�JJJJm�z��z`H�i��i ��i�h`H�م�مh`HH�dd� �F�eJf����h`H��� � >�h`H�ɠ�� �� >�h`Hڭ�:
�����F轾��G�E��D 7��h`H�Z�H��:
��6���7��� ��

e����ȱ��ȱ��ȱ��ȱ����
��h�z�h`Hڢ ������8��������h`H &������� kĊm� �� >� &� '�h`H� &������� kĭ:���� �� >� &� '��h`H�H�9ɠ�5����� �٭��%��H
i����� ��h:
��


�� ��h�h`H�Z 7� � �D)�8 �߰3��F��* ����� �� 7� � ���F���� ڈ��� �� 7� � �z�h`H�F���E)�� ޭ��F�E)�m��Eh`H�Z 7� � �D)��: �߰5��F�'�, d���� �� 7� � �ɠ��F�	��� �و��� �� 7� � �z�h`H�F���E)�� �ݭ��F�E)�m��Eh`H�Z 7ޢ ����� 7�z�h`H�Z �߰
�G�� ��z�h`Hڢ�G���E)�JJJJ�� ޭ��G��)



H�E)�EhmE�E����h`H�G���E)�JJJJ�� ޭ��G��)



H�E)�EhmE�Eh`Hڥ�� 7ޢ E���� 7��h`H� �� 
��d�
�G�� b��h`H�G���E)�JJJJ�� �ݭ��G��)



H�E)�EhmE�Eh`H�Z����d�� b�:���z�h`Hڭ����� �٭���:H
����8���-��)


m�� �ɰ���


m�h



��h����h`H�Z�H�H�H��	��)�L�ݽ���������H)�h)�JJJJ� �ܭ���5��HJJJJ)
��`���a��hH)

�hJJJ)
e���ȱ� �h�h�h�z�h`HZ�H�H��H 
٭������ �٭��
�H�iȅ�i �h8�
��

m�

m������)�JJJJ�)��h��h�h�zh`H��i��8��������h`H����8����	i����h``HڥH�H�H��	�F���G���EH)�h)�JJJJ� �ܭ���$�DH)

�hJJJJ)
e��p���p�� �h�h�h��h`HڭD)�������������	��h` �ހ� ߀� "߀� A߀� `߀� q߀�H���� �� �D�
 �߀��Dh`H�������D�
 �߀��Dh`H�������D� �߀����h`H�������D� �߀����h`H����D� ��h`H����D� ��h`H�,D�
��-D�D��D�Dh`H�E)�	�F: �߀h`H�E)�
�F �߀h`H�H�E)�����h���G�� �ݭ��8�������h`H�E)��	�G: ��h`H�E)��
�G ��h`H�H�E)����h���F�� �ݭ��8�������h`H�Z�H� ��

e� ݹ:�����  � �� � �� ݽ�)p�0��@��`� � �� �� �� �� ���
��h�z�h`H�Z����� ���� ��z�h`HZ�������)�� ޭ�����)�m������zh`HZ�������)�� �ݭ�����)�m������zh`HZ�������)�JJJJ�� ޭ�����)



H��)��h}����Лzh`HZ�������)�JJJJ�� �ݭ�����)



H��)��h}������zh`H�<��
��=��������h`H��)���<��
��=������������=������h`H��)����� ^� ��� ��� �h`H��)����� �� 7� K� ��h`H��)�	��: n�h`H��)���)p�p������ n�h`H�ZH��)p�p���)�������)�����h������ �ݭ��8������z�h`H��)��	��: ��h`H��)p�p������)��
�� ��h`H�ZH��)p�p���)����h������ �ݭ��8������z�h`H�Z�H� ��

e� �����h�z�h`H�Z�H�
��

e���)����� y� ݩ���  �h�z�h`H�Z����ڭD)�!������0��,��(��3��7�z�h`��t���F���G���E������u���F������v�����w���G��� �F���E)�� ������������)���E)�m�����H�Z�H�
��

e���)� ݽ�)����� � *� �� �����h�z�h`H�Z�H�
��

e���)����������������h�z�h`H�Z�H�
��

e���)���)���A��H����h�z�h`���F���::�G���)�JJJJ��E)�JJJJ��� �8�ɽ�:�F�π�������)�� � ޭ��F𱀚H�Z�H�H�H� ��

e���)�=�����)p��������� ����)p�`�
 ݩ�����:� ����
��h�h�h�z�h`H�F��:����+�F�'����G��:�����G����8�h`H� 7ޢ������ ���H��H� ��	�D��������  � 7ޭ��d� �ܭ����� 7� �����  ��������$������  �d$�H� `ש �� ���h`H�Z�H�H�H�H�
��

e����)������� ������h�h�h�h�z�h`H�Z�H��H��H� ��

e���)�"��)p�0��@��`��������� ����
�ɀ %�h��h��h�z�h`H���� ������������������8�h`H������  � ݩ
����H��H����� �٬�� �:h��h����=���� ݩ{=����h`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             L-�LE�Lj�L��L��Lr�L��L1�L}�L��L��LD�L��L��L
�Hڥ#�_d 7ĭH� r� �� e�d� *� 7� @�$� �� �H��$�d��� *����  ��� �Ād�� *���������h`Hک  �� �����d���	�� ������h`H ��  � |� @� *�h`H�Z�����������Q�������� ���y��������z�h`Hڮڮ����� �ŭ� �ŭ� �ŀ�� �ŭ� �ŭ� �������h`Hک=�������������������� �������h`H�H�H� j�+��� �ŭ� �� ��h�h�h`H�H�H�H�� j� ���� ��h�h�h`H�H�H� j�4��,� ǩ j��m��m� ǩm��H ��h�h�h`H�H�H� j���\� �� ��h�h�h`H�H�H� j���L� �ũ �h�h�h`H�
�����轘���h`Hڭ��� ���������h`H�Z�H�
��

e�������h�z�h`H�Zdd#�� �� 7Ģ � �
�������� j� �ȩ j��g� ǩ j� ���i� �ũύ& ��� *��� h̀��  ��� �ĩ���#z�h`H�Z�H� ��

e���H)�hH)��������:���� �h��
��h�z�h`H�Z�H� ��

e���H)�hH)�������h��
��h�z�h`Hک �	� �����	 j� � X�o������d����� � '� X�������� � '� X� 7ĩ��T� � '��  �< X�:��h�`�H�H�H�H�����
 j� �h�h�h�h�`Hک �/:�������h`�Z�/���� ���� ��z�h`H�H�H�H�H�Hd 7� ��  ��'ɿ�� �ĥ��� �  H��d�  � H�ҥ� ��� ��8h�h�h�h�h�h`H���<�� j� �ũ(��n�� j� �Ţ  �h`H�	H� �	� ��h��8��
�h��j�� j� �h�	h`H�	H� �	� ��h�i��8�i���h�i��j�i� k�h�	h`Hd � 7� �� 7ĩ ��P�� j� �ũ2 *ש �� ���h`                                                                L�L��Lc�LL�L�L��L�� �P�Q�R �� �� � � � � � � � �* d�d�� ����d�`�Q����y� ��r� �s�  G��y�y�t� U�R������ ��� ���  ��憥�Ł� ��P���J�Q����]� ��V� �W�  ��R����k� ��d� �e�  ���]�]�X� ���k�k�f� ���� �� c�`�S�T�VȱT�WȱT�XȱT�YȱT�Z)
��4��[�4��\�Z)0�`ȱT�����ȄSd]d^�X� �L��_ o�� �
�T� �d_��Ȅ_dS���o�p�rȱp�sȱp�tȱp�uȱp�v)
��4��w�4��x�v)0�{ȱp�����Ȅodydz�t� �� �Q� ��)��	���Rd| ��`�|�}�ȱ}��ȱ}��ȱ}��ȱ}��)
��4����4�����)0��ȱ}�����Ȅ|d�d���� к� �R� ��)��@Ы���Qdo U񀠤a�b�dȱb�eȱb�fȱb�gȱb�h)
��4��i�4��j�h)0�nȱb�����Ȅadkdl�f� й�m ��� �
�b� �dm��Ȅmda����
��������������Tȱ��U`��
��������������bȱ��c`H�Z�Y)?	@���Y;��%����^�[��Z)@��J������`�8��`��Z)0�`Ȅ^�[����^�Zd^��� z�h`H�Z�g)?	@���g;��%����l�i��h)@��J������n�8��n��h)0�nȄl�i����l�hdl��� z�h`H�Z�u)?	@���u;��%����z�w��v)@��J������{�8��{��v)0�{Ȅz�w����z�vdz��� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ƈ��d���� z�h`� `� `H�Z���������������)?
������轖���d� (�z�h`d��* d�`������ȱ���ȱ���ȱ���)
��4����4�����)0��Ȅ�d�d����  �d�`H�Z�����L��������;��)����������)@��J��������8������)0��Ȅ������Ɛ��d���)����)����
�@����������( ��ŕ��* ��捥�Ō� (�z�h`H�Z�  o�  ��dSda��_�m �� � �� �� ����Pz�h`H�Z�Q� ��R� �d���)?Ŝ�D�� �>��
����p�(��}���q�(��~dod|� �Q�R��)�����R �����Q U� ��z�h` q<� � �<�!� q<� � �<�!� qZ� � Y�!� �x�!� �<��� �<�!� q<��� �<�!� �<��� �<�!� �<��� �<�!� �Z��� ��!� �x�!�     � YZ��� q�!� YZ��� K�!� ��!� ��!� ��!� ��!� �x�!�     ���!�h�!�.�!  ��!� ��!� ��!�.�! h�!���!�h�!�.�!  ��!� ��!� ��!�.�! h�!�     ���!�h�!�.�!  ��!� ��!� ��!�.�! h�!���!�h�!�.�!  ��!� ��!� ��!�.�! h�!�     ���!�h�!�.�!  ��!� ��!� ��!�.�! h�!���!�h�!�.�!  ��!� ��!� ��!�.�! h�!��<�!�.<�! }x�!�     � � � q�!� � � ��!� �(�!� �(�!� � � q�!� � � ��!� �P�!� � � q�!� � � ��!� (�!� _(�!� �� � �!� �� �     � ��!� �P�!� T� � K� � G� � T� � d(� � (� � T� � K� � G� � T� � dP� � � � q�!� � � ��!� �(�!� �(�!�     � � � q�!� � � ��!� �P�!� � � q�!� � � ��!� (�!� _(�!� �� � �!� �� � ��!� �P�!� T� � � � T� �     � � � T(� � ?(� � T� � � � T� � � � T(� � ?(� � � � d� � T� � d� � _� �     � �P�!� �P�!� �P�!� �P�!� ���!� �P�!� �P�!� P� � �P� � �P� � �(� � (� � �P�!� �P�!� �P�!� �P�!�     � ���!� �P�!� �P�!� �P� � �P� � �P� � �P� � �P� � �P� � �� �     � ?�� ?�� ?�	� ?�
� ?�� ?�� ?�� ?�� ?�	� ?�
� ?�� ?�� ?�� ?�� ?�� ?�� ?�� ?��     � �
�� /���     � _� � d� � q� � � � �� � �� � �� � �� �     � /�3� 2�3� 8�3� ?�3� G�3� K�3� T�3� _�3�     � ?(�3�     � K� G� K�     � T� O� T�     � ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���     ����������OA 4    ( H h � � � � �    ����������_�?�/�   (    	
	�
	�
	
�
�
�	�


				�
				�	
�
	�


	��������������~���  ,�����  p���f���  8���  ��  ��          R�d��������R�d����������� �+�0�5�=�}�������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �� �O�