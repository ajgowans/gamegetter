 ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������?���������������������������������������C���������������������������������������T��������������������������������������?U��������������������������������������_U��������������������������������������WU��������������������������������������UU��������������������������������������U�������������������������������������U�������������������������������������_U�������������������������������������WU�������������������������������������WUE�������������������������������������UUE������������������������������������UUE�����������������������������������_UUE�����������������������? �����������_UUE������������������������ �����������WUU������������������������� ����������UUU�������������������������? ���������UUU�������������������������� ���������UUU���?���������������������� ��������_UUU�� ����������������������? ��������WUUU� ������������������������  �������UUUU�������������������������� ������UUUU���������������������������? ����_�UUUU����������������������������  ���W�_UUU���������������������������� ���U�WUUU����������������������������  ��U�WUUU�kUUU�����������������������?  �U�UUUUUUUUUU������������������������ �_UqUUUU�
 PUU������������������������  \UYUUUUꫪTU������������������������?  �UVUUU��^��U�������������������������   �UUUU������������������������������ �uUUUU�ʪ�����������������������������?�jUUUU��Ϋ���� ����믿����������﾿����[UUUUU�������3 �����������������_UUUUU����:����Ϫ�* �ﻮ����������������^UUUAU����>���������
 ��������������/���U�U����?�����������
࿻����������������V�U���������������
�����������������UU�
D�������?TUUUU����
���������k�9��PUU   ������@UUUYUU�����뺻�����g�U*�?QU    �����    BUUU�������������I)�?UTUP    ���?       @UU�������v�U��OQUUQU                DU*�������޾�e��WQEQUUU           @UUU�������������UUUUPUuUUUUUUUUUUUVUUUUU�:���*�꺯���WUUUUUT�UUUUUUUUUUUYUUU������� ������PUUUUUUUUUUUUUUUUUUU�����j������j��?QUUUUUU UUUUUUUUUU������j������
 ����?@UUUUU����������������꿪�������* �jf%�DDUUUUUUU��������������j�����������UUUUU�UUU�����������U����������
 o�%�DYUUUU}U�UU���������UU������������ ��YfUUUU_U}UU�����UUU�������������� �*��efUUU�WUUUU����jU�����������������
 �+�YUUUUUUUUUU����������������������* ���YfB@DUUUUUU�����������������������  ��_fVUUU  TUU������������������������ ��gYUU�W�iPU��n���������������������*  �UU�E�UU�j ����k���������������������  |UUUU�Ue������������������������������ `UUUUU��
����������������������������
 XUUUU   ���������������������������zUVUUUUUA��������o���������������������Z�UUUUP����W�����Z���������������������V�UUUU�����W�������꼪�����������������UUUUUU YU��U��UWտ��������������������jUeUUU@�����U��������������������������ZUYUUU������S��������������������������VUVUUU���������������몪*��������������UUWUU �����������������*������*����jU�UUU@���  ��������󮮪������*�������XUuUUU�+���������������������*�������(�VU_UUU ���?��������������**�������������U�ZUU@/*������������?/�������*�*�����jU�WUUЃ*� ����������<**����*(�����"�"XբUUU�?�"�������������(
�������(��(V�zUU@���� �����������?�à�*(��(�*�����XZUU������� ������������������� �"�(�(XUU����� "���������<�� �"�

��"(�� VUU@��  �� ����������̢ �� � 
�*����UU��?   � ���������ʀ� 
"
����
�(`UU�����  ����������/ *�� "�� ��bUU�����   ����������� (       *��  *XU@         ����������   � ""�" " V����  �?� ��(�>� �  �� ���    �U����? ����?�(�� �  ��� 
  ��  � `U�O�� ��<�?� ���?� ���      ���`U�� ��?�� � ��?� � � (�  XU��  ��?��������?� �? �?     �    VU�?  ��?�������� � �? �?         �U�  �����?���  � � �?   �    �U�  ��?��?����� �  �?�         `UA�  ���?���?����?� � �?        XU��  �� ?� �����?� � �        X��  �            ���� � �?          p=� ��            ���� �? �?         �A� �?            ���� �? �?           �� �  ��  ���� �� � ����             ���� ��?� ������ �  ���             ���� ���� ����� �   ��              ����� ��� ������   �               � �����? ������ ���              �  ����������� � ��?              �  ���������? �� � ��?              �  �?������������ :���             �  �?����������� ����?             �  �?����?���?� � ����            �  �?������?� � ����            �  �?������?��  �+����           �  �?��� ����?��� �����?�           �  ���?�    ������ �����            ���         ��� �? �?            ���          �� �� ��         �� �               � ����         ����                    ���00        ����?                    �? �?�0      ����                     �� 0��<    �������                    ��   �?   �����0���?                    �   �?  ������ ����                   �   ��  ���������������?               �  ��� ������������������?                  � ����������������������                 ���������������������������            ����������������������������           ������������������������������          ��������������������������������        ������ �<���? � � ���� � ���      ��������������?������������������    ���<<���������?�����3���������������  ����?����� �������3��������������? ����3�������������<���������������?���<<������<�������� ��������������������������������������������������������������� �<�������  0����� ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������?0�� ���   ����?�?�?����������������?�����<<��?��������������?��?�����<<������������������������?����?���������������������������?��?�����?���?���?��������������?��?��?�����?���?��������������������?��?�����?����?�?���������������?�?����� ��� ����� ��������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            TUUUUUUUUUUUUUUUUUUUU                                                           TUUUUUUUUUUUUUUUUUUUU                                 ��                       TUUUUUUUUUUU���
�VUUU                               $dUPU��                   TUUUUUUUUUUU
U�U�Z
 �                              @ZUUUeUUU                   TUUUUUUUUUUB&�ZVUUUU                               	TPF@                        PUUUUUUUU  �
TU�                                * ��
                      TU    @UUUUUU�jUUUUU                                                           TUUUUUUUUUUUUUUUUUUUU                                                           PUUUUUUUUUUUUUUUUUUUU                                                           PUUUU  DPUUUUUUUUUU                                                           TUUU        @UUUUUUU                                                           TUUU    DUUUUUUUUUUU                          EQA                              TUUUUD@TEUUUUVUUU                      @        �                        TUUUUUUUUUUUU��UUUUUU                               ?                         TUUUUUUUUUUUUU\UUUUUU                                                           TUUUUUUUUUTUEQUUUUUU                               @                          TUUUUUUUUUUUUQUUUUUU                                                           TUUUUUUUTUQUUUUUUUUU                     �    <                             T��UUU?@@TUU{UUUU                     ?     �      ��   �                   TU  @Q  Q�^WUU�                     A R`(
       �  �                   TU�UUUUUUUUUUUU�CuUU�                   TUU     ��     � �  �                    PUUUU���_UUUU�UWU�                   TU    ����    �                      TUUUUUU����WUUU�:PuUU                       < ����    ��                     TU�W�UU���WUUUU�UWU                   T��    <  �    �^                      <TUUU=  �WUUUU�zQ}U                          <  �    @��                       @UUU����TUUUU���U                      ���V���� �  ����                      ���������WU}WU���_W                       ����?���s ���W                         �3����]U�n�UW                       U��=  �|@� ��~��                          6��WUw_��U                      @UUU����   7��UUu                          ���sU���UUUU�                     UUUU���jUUU����w                   T     �� UUUUU�UU~u                   TU  ����pUUUUU�U�~u                       �_Ѓ�zUUUUU�U�~u                    @��P��*�WUUUU�U�~�                     ��_������UUUU�U��u                   T����ߏ�����UUU�U��u                    ������� �jUUUW��u                   ����p�ի*W[��WUUW��u                   ����Oui��U�����W���                   ����\]jU�rU��j���W��u                   ����e�^��\U�檰��W��u                   ���?e��_=\}�����W��u                    ��i��W=W����������                   TU�Sꩯ^�U�����������                      �ڪ�z������VWU����                   TUU�����w��: �VWUUUUu                      S� ����: �V_UUUUu                   TUU�� ���������_UUUUu                     Ф������ꪮZ]UUUU�                   TUդ����ꪪꪫjuUUTu                     0��﫪���?����U�Ru                   TUM��ꫪ������U��
u                     L��着� �<��j� ���p                   (PM������� ���������                   �
_������������������                   ��W������ �����z�����                   �����W��������o�����                    �����  �
 ���W_UUUu                     ����SU@  ���WWUUU�                     ����G  h ����_UUUu                    �����  � ����wUUU}                    p������j��{�UUUU                    p���������*����uUUUU                    p������着�����uUUUU                    ���������
 ���}UUUU                    �������몪
���vUUUU                    l��_�������?�j}EUUU                    \�������� _�j5UUUU                    ���T|TQ�� �*�vTEUQ                    ���U}UU����*?�_=@UU                    ���A�
�ꪪ���_5TTTU                    ��� ?������+���UTU                   ��?�_"��ꪪ*���?@UU                   ���տ���ꪪ*���?  @A                   ��������ꫪ����?TE                   ���_����������W�  P                   ������?������_�@@T                    ������������W\�  @P                    ��������������AD                    ������������0  TP                    �� P���������� DT                    ��  ���������W?�  D                    �?  ����������� @                   Ԩ�UU����������                      ���  ��������� �?                      ��?��������?�<                      ��  ��������? �U�                      ���  ��~߿���; k�                     @��UU��������{�ZU<                     <� P���}����?�z �@                   T TU ��������?��U�                         ��������?�{                        @�������?�lU >                       ���V���?��  :                    @  ��U������V :                    T ����������jQ :                         ��j�꾪�j��:                    P@ ��_U���j��:                    P @ ��������ïj���                        ���V����ïj���                      @  ���������ڪ��                     D ��^U�����۪��                    P    ���j���������                      @ ���Z��������?                         ��zU��������                         ����ή�� ���                          ����Ϫ��  �                           ����Ϊ��                               ����Ϊ��?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �?����<�?<?� <�?  ��� ��?�� � <�� < ��?�� � ? < <� � ��3�<<�?����� < � < <� ��� �<<<���<�< ��� �  ?�����?<��?��<�<<�? �? ��00�?<?��?�����?�������?����<�< < <����?��<���������<��������� ������������ � ��3<<0 ?0<<���<0<0�?<0<0<0���������� � < < < <<<<<���<0<<�<<<���� � � � �������<<?�?�<�<<?��<0�0�3�??<?0��<<�<�<�<��<��?�������?� � ��?��<�<�<�<�<��?�?�����<��<�<����<�<���?�<��?�������������<0<0<0<0<0�<���<0<0�������<�<�<��?�?��?�<0���0<?���<0��������� � ?������    ���                      ����������������  � � `X	[9`�,�6�,�6�,�6�@�J�T�J�T�^�T�J�T�J�h�J�T�J�T�^�T�r�|���|���������������̃փ���J�T�������&�0�:�D�D�N�X�b�l�v���������������������������ƄЄƄڄ����������������������UYYYYWVYYYYXUJYYYWVYYYYYXUYYYYYWVYYYSXUIYYYWVYY
YYYXUYYYYYYWVYLZYYSXUYY) YYWVTYYYYSZ UYYY$#$YZZ[[YZZ[[YZZ[[YZZ%&ZZUYYYZZVYYY	XU)*Y&WVYYYYYXUYYYJYWV(+YJYXUYYYSYWVYYYLYXU)*YLYYYWVYYYYSSSX*YYYYY	W[[YYYYYX[[[Y) W[[[[YYYXT$*YYYWTYYYY)TYSJY[[TYYYY[[ !YUYYYYYYYYWVYYY	YYYXUYYYYYYWVYYYYYYXUYY	YYWVYYYYXUYYYYW����������������ÅɅυڅ������������
�����!�'�-�3�C�I�O���Z�`�f�l�w�}�������������������ʆՆۆ��������	������$���4�N�����T�����������n������������
@ �
p �
` � �
p � �
@ 
` ���
p �
@  �
` �� �
p �
` ��0�
` �
p ���   � �� �h �
@ � �
�   < �
 �
� �
h � �
@ �
h � ��� �4 �� �� ��  0�� ��X ��` � T� � � �X �T �( � �
� �
(   �� �( �( | �T �� X� � 8 X x � �T ��8�X�x����@0�� �*�4�>�H�R� �*�4�>�H�R� �*�4�>�H�R� �*�4�>�H�\�f�p�f�p�f�p�f�p�z��� �*�4�>�H�R� �*�������������ʈԈވ�ʈ���������$��.�8�B�L�V�`�j�t�~�����������8�������������������OPYYTYMNYYTYQYYYYHOPYYTYMNYYTYRYYYYJQRY'YLTOPYYYYTYMNYYYYYTRY	YTQY'YT'&YYYYYZZYYJJYYYYYYTTYYLLYYYYYYOPYYMNYYQYYYYRYYYQYYRYYYYYYYYYYYYYYY	YYYOPYYQRMNYYOPQYYYMNOPYYOPMNYYMNQRYYRQ          L�L�M�S�Y�d�y���Y�������������Ŋ��L�Њۊ������Њۊ��-�L��-�=�H�S�L�����^�i�t����������ʋ�������Ջ���L�L� �L��L��&�L�6�A�G�M�L�L�L�L�L�X�L�L�L�L��
P �
p �
@ 
` �
p 
`  � �
@ 
P 
` 
p �  � �0 � �
@ 
p �
H 
X 
h �X � 0�0�
P @ �
` p �
P 
` � � �0 � �0 t �0 p �
@ 
` X �
P 
p X �0 � �
H 
h �( � �
  P �
� ` �  � �
  P ` �
� p @ �   � �� � 0 �  � �( � �
 
( � �
� 
�  � � �D h � �X �
H 
h �
X 0 � �
H 
h �
X�T �4 t �
.L��
���(�2��
���(�2��
���(�2��
���<�F�P�Z�d�P�Z�d�P�Z�d�F�n�x���������������������������ȍҍ܍��������������������܍��"�,�6�@�J�T�^��h�r�r�������������������OPYYYYYYQMNYYYYYYTTTYYYYSYY67YSYYYYR45YYYTTYY)+YYYYY[[[YYOPY[[[YLMNY[[[YTYRY[[[YYYYY(*YYYYYYYYYYYYQY)+YRY[[[[[YTY[ZZZ[YQY[ZZZ[YRY[ZZZ[YYY("*YTYYYYYYYYYYYYYYYYYY)#YYYYYYYYYYYOPRYYYYYMNYYYYYYQRTYYYYYOPQYYY(#$ YYYYYY67YYSY45YYTYSYYBCTYY@ASLYYYSSYYYHSYYYYYY�����%�0�;�K���%�[�f�q�f�|�������������������ȏӏ��ӏ�|��������	���*�	���	��5�@�P�@�P�@�P�@�P�@��`�f�q�w����������������̐������
` �0 �
` � �
` 0 �< P ` �
`   � �D p �0 � �P h �X  � �� �@ 
� �� 
@ X �@ 
� X �  � �X\ �  T� �` �
0 � @ �0 
� � �  � � � �0 � �8 | �
  � �
  �  �
  � @ �X �  � �T �  � �
H 
X 
h �$ L x �
@ 
P 
` 
p �H d  � �:@��~���~���~�����������������������đΑđΑ��ؑ�ؑ⑰���� �
��(��2�<�
�F�P��Z�2�<�
��(���� �
�F�P��d�n�x���������������������������~�������~���ȒȒȒ������������������YYYYYYYYYYYY67YYGG45YYFF>?SY23<=YS01>?YT:;<=TY89T6767YY4545STYYYYYYYYYYSYDEDESTDEDEYT67BCYY45@ASY./BCST,-@AYYYYYYYSDESDESDESDEYYYYYYYKTYKTYITYITYYYYYY!#$ n�n�o�u�{�����������{�������������Ǔғݓ����	��)��	��>�S�^�n�~���n���	��)���n���	���n���n�����Δ��Δޔ��Δޔn��n�n���n�(�n�.�n�n�n�n�n�n�C�n�n�n�n��
P �
` �
@ 
p �
H 
` 0 �@ p X �0 � �
` � �
P   �H d �( � �@ p �0 � �  � �
( � �
� ( � �
( �   �
  
0 
� 
� �
( 
�   � �0 t �
  � 0 �  
� � �
  
� �  0 � � �( � �  P ` � � 
X � �
` �  � 
P 
` � �X  � �
H 
h �X 8  x � �T ��@�h����
!L��        PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUU        UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   �   �UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUU��������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU���������   �   �PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU�PUU���������        PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUU��������        UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������   �   �UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU���������PUU�PUU�PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUU�PUU�PUU�PUU�PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUU�PUU�UUU�UUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUU�UUU�UUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUU�PUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UU�_UU�PUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUU_UUUPUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUU_UUUPUU�PUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�_UU�_UU�PUU�PUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�_UU�_UU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UU�_UU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUU�        UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UU�_UU�        UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUU_UUU        UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUU�PUU�PUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������PUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������UUU�UUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������PUU�PUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUU�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU        PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUU�PUU�PUU�PUU�PUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUUPUUU��������   �   �UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�_UU�_UU�PUU�PUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU�UUU���������  < TU�UT��_T���D��4��<D��<��7D��7�3D��7��3D� 7�7D�3�    ]UEUUEUWGWUEWU WUEWuE�����������   0���:   0���7D��7��3D��7��7D��7��3���7���7��������꫷��믪�꯾�z���_       �����W�����u�� �jE�ZE�VE�UE{] _UEU�EUUE�UE      ��TQ5�TQ=�TQ=�TQ=�  ?�TQ3�TQ3�TQ?�TQ3�  ?�TQ3�TQ?�TQ3�TQ?�  3���   c  k  k  k  k  k  k  k  k  k  k5  k  k  k  kTQ?�TQ3�TQ?�TQ3�  ?�TQ3�TQ?|TQ�TQU  sUTQUTQsUTQ_UTQ_U  _U  ��  k  k��k5U�kU�kU�kU�kU�kU�jU�jU�jU�jU�ZU��U�U�_U�+  ��T�S��_Z�_��_������0�����?������������`i�    �TE�SE�OE�?E�? �?U�?U�? ���+���*� ��� ������0���?�� ���0 꿬������?����*�
�� �����h��������U �OU �   ��:��;���&��*�����p��ԩ����j������������UUUU      ��TQ5�TQ=�TQ=�TQ=� �?�� 0�4�?�<��0��<��0��<��0��<��0���   c  k  k  k  k  k  k  k  k  k  k  k  k  k  k<�30�3�>�3�3�� <�C�3�U=|C���}UL�uUUuUtUuU��_UTQ]UTQ]U  ��  k  k��kU�kU�k��k��kU�kU�jU�jU�jU�jU�JU�RU�T�  ����  ������ ��� ��� ��� ��� ��� ��� ��� ��� ������������  �    TQESQE�� p�
0 �
��
��
��
��
� �
��
��
��
��
�   �  �����\UU�tUUU�UUU�WUU�\UU�pUU��UU� WU� ���   �   ���� ����
��
��
��
��
� �
��
��
��
��
� ��� �  �  ���� �������������������   WUUUW�WU_5_U]5_U}�_UuUUUuUUU����U���U���U������_���o���{���{   �UUU��WU�5_U�5_U��_U�UUU�UUU�������������������p��?p3��z3��z� �{��{;��{,0�{���������������T�WUTUU]tUUU    ���}��U��U��U�� U�����}U�WU�UU� UU�UU�WU�WU����    ����������������   WUUUW�WU_5_U]5_U}�_UuUUUuUUU����U���U���U������_���o���{���{   �UUU��WU�5_U�5_U��_U�UUU�UUU����������������� � �D}UD�WD�WD�WD��D��D��D��D��D��D��D��D��D��D��D��D��D��D��D��D��D��D��D������ ���û��  �  �����U�UU��U�"�W���o-"�n���o-"�n���o-��n�|�o�W�n}�_ouUWmuUUmuUUm���_���U}U�Ws��^sW�~s���s���sW��s���sU������sU������_UU�����WUU�����T�_U��U���_T�T��U��U��CU��]U�z}U�^�U�_5��_5��_5��_Ք�WT��U��U� _=�|��<<��?�|>���  �3  �����C���M��M�����_U��U���W_W��^W��^���^���^���^���S�_W��^W��^���^���^���_���WTUUUU�UUU�WU]�U��zU���U���W5º~M���M��?�������c�����n����zU��UUUU�WUU5_�U5~UU{UU�U]�~_U �jU���U��W������w�������p��>��^� ���0�5n�-���°����p��𲕯��U��U���]շ�UU���U��UUU��p�W��U��Wu��_U��W��~���{߾�_���W���U��_U��UU�Uu�WUU�UuU_UUUU�UUU�WUի_]5�zU���U=<�u�U��W��^à�^��~3 ��=��5���լ�_U�_UU�UUU�_UW�^]U�~U���U5 �W���~��� ��
�����5��~�˫_U�UU=_UU�WU�WUU\�_�p|ͳ���� ���S��_x�\�?3p��ps�]_�]}Wr}UU]uUUUuUU_UUU]U��su���U���U��_=���/�}0�7 �����M�(=.��������U��U �p �P �P �P  Z@  Z@  Z@ �P �T �T �T �T �t �P �P �P  Z@  h  h  h  Z@  Z@ �P �P �T �T �T �T �t �T �P �P�  �  � � � � � � �  �  �  @)  @)  �  �  � P
 P
 P
 P
 P
 P
 � � � �  �  �  @)  �  �  �  UUUU]UUUUW]UUUUUUUUUUUU]UuUUUUUUUUUUUUUUuU��UUUUUUUUUUUUUUUWuUUU   �T�T�d�d���������d�d�T�T����� � �T�T�d�d���������d�d�T�T�����UPUTTUUPATAPPTAAUPUTTTTUPUTAAPPATAUUPTTUPU �  p  � 0��p7�>;��;ܵ^7|w�=��7W����]u���������������?�  ��� ��i�w� �� �w5 ���?�Yj��Yj����?�w5 �� �w� ��i��� �  0�<�<���?����ii�V�sV�ͬUU:�UU:sV���V��ii������?<�<0�    �0����ii�V�pV��UU:�UU:pV��V��ii����0         � �aI����V��Ye`UU	�UU6�UU6`UU	�Ye�V�����aI �             0`	@���UU�Ye`eY	�UU�UU`eY	�Ye�UU@��0`	          ��|p=���6|]u=�޷>\[�5|��=p��p[�p}}��W����� �  �  �   � �� ����]������z�:��� ��  ��  �;  �     0�    7�  @7��p;��]u�:����:���� ��_  �ii?   ��    0    �    �   �  �� �3�p�Wp_W���W�W�W�W����p_Wp�W�s� ��   �   �   ��    \��   ��uY���}���=p�uuu�5ܹ�uݹ�\��wo�����wo��\��wo��ܛ�wߛ�|W�u}W�p�w�u�7��u��? �w�   �      0     ��  WU  ��  WU������UUU��U�W���U}��]�����U�?���?��W��\�U]�\ת^�\ת^׬�U���W������몮�\׫_�\��\׬� ��� ��\� \��� �� ?   �   7 �?���������7_��_����7�������� w  �   ?        �        ��           ��         �          ��          ��          �5 ������? p�          �5 �������� p�          ���UU�WU�?|�          �V�_U�VU�W��W�     ��  �j����VU���[��   ?��|  �����U�ZU����  ����_� �����eg�����?  ����_���������ٟ�����?�����\_������jU���U���������\]u�����VU��^UU����u��\]uU����VUUٟUUU����Uu��\]}U�z��VUUegUUU���~U���\_}����_���Z������^�����_}��������_�����_������������W�\U�����_�������������UW��������������w��Z��UW�_���w���?��������Z��WW���������?��������Z��_�o��������� �����z�Z�������������� �������Z�������������   ������ZU���_U�~�����    ������kU�_�U�����     �����������������     ����ޯ�_����������      �������_���������?       ���z��_���������       ������_���������        ����_}������?        ������^_��^����         �����^WU�^���         �����^WU�^߫��         �����^WU������          ����^WU�����?          ������WU�����           ����UU�꭪�           ����UU�ꯪ�            �����UU�z���            𫪿�UU����?            �����UU�ު�             ��~�UU����             ����UU����              ��WUUU��>              ���_UU���?              ���~UU���               ���UU���               ���WU���                �����>                �ꯪ�?                �������                 ��_ի�                 ���_��                  ����>                  ����                  ����                   ��_�                   �_ի                   �~��                   ����                    ���?                     ��           �  �  �5  w7 pww\]]w�w7wWu7w�@77� 7� 4  0  �    0    ��   �UU?  ��_ ����\��W5\�]uw5��p7�  @7�    7    0�  ��:[��[��W�����Z
��Q0�                 �  �:  +�  �  �  +�  �:  �                          �?  �� ���@�  �  �  �  �@�� ��  �?         ���પ�@..  �  �  �  �  �  �  �  �  �.  ��@.પ����l9[�[�k���?�P   TU  UUU ������� ��  �           P   TU  UUU ������� ��  �        U UUU���� ���  �?                U UUU���� ���  �?        <   <�   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   ��   �<   < 0   0   0   8 ,  � .  � �  � �  � �  � � �� o���n�~ý��Þ � �  ( ( ���������?�������������ö������ö������ö������ö������ö���� � �  < <  �  �� �����Z�>�V�>�UU��UU��UU��UU��V�>�Z�>���� ��  � �?���������������  �  �  �  �              0  �  �    ��       �UU      \Ye5     �WUU�    |i�Vi=    Wj�Z��   ��Z�j�V  ��Z�j�Z  peUUUUY  lUUUUUU9  l�jT�Z9  l�QE�[9  [�F�^k�  [z��W��  �^�Z�W��  �WU[�U��  �UU�zUU�  [UU�_UU�  [U�UU�U�  [�PW�W�  [5T]u\�  [U^�Up�  �C�^�V��  ;P�_�Z�  �W�W�k�� �U]�UU�uU���~UU�v���UU��0 ��UU�� � �W���� � �UUUU? � |�_�_= � |����= � ���/�� � ��((
� �<��� �<���? �_� �������   W���W�    TUU�    l@UU9    �VUU�    �[UU�     �UU:      �       ��    �           �_�           �W�         �W��W         ���|=         |=���         _���       ��?��_� � �? ���?  |�?W p��W=    �U�U �U_U    �Wu� �_]�     u�   _]�      p]�   Wu      �]U �Uu      �]U5 \Uu      �WU� WU�       WU� WU�        WUU�UU�        WUUUUU�       �WWUUU��      �VWUUUՕ      �V������      �V�U}U�      �V}UUU}�     � [�U�w�     �[�UUU��    ��]Uu��0    ���WUUU��?    ���UUUUU�    �P�jU�j�    ��W��U���    ���׵�^��j    ���_�����V    �Um]UUUuyU     SmwUUU�y�      m�UUUwy0      ��zUUU�:?       ��WU���        �3oU��;        �3oU��;        ��U��?        ������         ���W          �U�U          �U}U          �UUU          pUUU          pUUU          puU]          �WU�           �U>            �U            ��            �<            �             ��             �              <         ������   �UUUUUU  |U����U= �W��UU�_�pe�u�W]_Y\Uu����]U5\UmYYeeyU5\U[���z�U5\�V�Z�W�W5\�VU�jU�W5\�zUUUU�W5\��^UU��~5Wm��UU[y�Wk��^�Z��W���^�����W���_���{�W���Wժ�z�\���UUZ�^5\ՖjUU��W5�U�uUU]�U7\U��UU��U5�_����__�?�Y��o��^e���my�Wg�YUsmy�Ue���s�ͪj�YUs�W�Ue�������� ��>  �[�  ��  �[>  ��  �[  ��    �       �    0@P`p��������  0@P`p��������  0@P`p������������������������������������������                                          ���ة�� ���  ��� � � � � � � �ύ& ��" � t ���� �� �� � ����� ���� � U�X�d� �# L �H�Z�� � � �P0� � �� �� :�z�(h@H�Z�' )��� ��� K� ^� �# �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                                         ���  � h�  � � � � ��  �� �� ��  �� � �.��� �� � �  k� #� -�  � qǩ ��  ������� ���� $� f�ɠ��i��Lt� aʭ� ���
� ���I {� |� �� `�)�� A� �� έ� ��� ��� ����� �
��8��Lt� �� Z� � ���h�� � � qՀ k� � ߭� ��� hح�M}��m �� � ��LY���������� �ͭ� �������� LY� �ǭ.�L7�L� ��� � ��  �� �� �� M�L  ��� ��LB� �ʭ� ���
� ��� {� �� �� �� �� �խ� ��� d� ���- Z�-)� �� � ���Lbí� � � 0ŀ	 �� K� �� �� �� �� &� �؜������ ���Lr�L�í� �����	�-)���-)�	 ]� k� m�`H�Z  � ����  ����(��� #� �� ����4��� #� �� ����D�� #� �� ����P�� #� �� ����`�� #� �� ����l�� #� �� ����x�� #� �� ��
����� #������  ����0� ��  �� ��z�h`�� �������-)�$��-)���-)���-)�	 �� q� ��`H�Z��� �� � �� �� � �/� ��X� ��� �� � �� � �-���z�h`H�Z�  ���������  �� x�  ��G���������� #�	������ #� ������� � #�  ���� ���  �� ��z�h`H�Z  �@����� i #�X���� #�2 x�� ��� �� z�h`H�Z� �����\������ � ��� � �� � f� �r� x�� ��d� ��� � � �� ��\��� f�� � � �� ����]� f� �D� x�L�� x� x� ���� ��\� �� i� � f� ��]� �� 8�� � f� �T� x�Lǩ���  (�< x�� ���ύ& z�h`H����� #��� #������  ]���  ]�#�� #�'�� i
 #�h`H�Z �� ��  �� ��  ���<�� #�
��\�� #������  ]���  ]��.�.�������  #���  ����
���. �� �z�h`H�� )��-)� kȀ
�-)� k�h`H�Z�  ������� ��	� 8�� L]����� ��	� i� L]����� ��	� 8�� L]����� ���	� i� L]����)� ��L�Ȯ ��Lyȭ 8�� � 8�� L]����)� ��L�Ȯ ��L�ȭ i� � 8�� L]����)� ��L�Ȯ ���Lyȭ 8�� � i� L]����)� ��L�Ȯ ���L�ȭ i� � i� L]���� ��L]���� ��Ly���� ��L����� ��L����� ��L����� ��L����� ��L���� ��L/���� ��L\����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L�����L��z�h`H�� ���0� 8��%� 0!� ������ �� � �� ��h`H�� ���� ������ �� � ��h`H� � �ʩ��h`H� 8�� � 8��  �ʭ i�  �ʭ i�  �ʭ 8��  �ʭ i� � 8��  ��h`H�Z�
��� ����(��4��E�Ґ� �Ґ� L|˽��� 轀�� L|˽t�� �t�� L|˽^�� �^�� ���z�h`H�Z�  ���i��L���^�
 x�� �� ������ � �������
 #�  ������L���� x�� �� �� �����z�h`H�Z� ���4� � � 8��� � �� �	����� �⩁��  (�z�h`H�Z� � �A�	������� 8�� �� � �� �0�� ��ݩ�� ��� � z�h`H�Z� � �9�	������� )�� 8�� ��� 8�� �� � ��z�h`H�Z� �� � �4�	������ �� � �� �0���� ��� � ���z�h`Hڢ � � �) �5 �A �M �� � �s �[ �g �� ��
0ة�� � �Y �Z ���	�
���,� �)�*�+�h`H�Z�
��� ������'��3Lν��� ���� L�ͽ��� 轰�� L�ͽ|�� �|�� L�ͽҒ� �Ғ� � ��Y �
.�Y �����$�� ȱ�) ȱ�5 ȱ�A ȱ�M ��Y L��z�h`Hڢ �� �00�g 8��%� 0!�� �"�[ �%�g �&� �#�s �$ ���	�L��h`H� � mΩ��h`Hڢ �� �0!�� �"�[ �%�g �&� �#�s �$ ���	�Lq��h`H�Z� �� � �LXϽs 8���g 8� 0�0LXϭ 8�g 0��� 

8���[ 8� 0�0LXϭ 8�[ 0��� E� �� � �� ���� � � �05�������'�� i
 #�����X� �ȍ ��	�L��z�h`H�Z� �� � �Lнs 8���g 8� 0�0LЭ 8�g 0��� 

8���[ 8� 0�0LЭ 8�[ 0��� '� E� �� � �� ���� � � �05�������'�� i
 #�����X� �ȍ ��	�Li�z�h`�[ �%�g �&� �#�s �$�� �"� � ����`� �� ��	������ � ����`H�Z� � �
00�M 8��%� 0!� ��) ��5 ��A ��M � ���Y �L��z�h`H�Z� � �
0!� ��) ��5 ��A ��M � ���Y �L��z�h`H� � �Щ��h`H�Z� ��� �
� �L���� 4�L����L'���L��� ��L����L?���L��� ��L���� ��L���� �L���� �L���� �L���� �L���� ��L���� +�L���� +�L���� +��Y �L�z�h`H�Z�,�,)�L�ѭ� ��L���� ��L���� 2�L���� j�z�h`�*����A ���A 8��A ����*��A Ɉ�� �*�	�A i�A `�)����M ���M 8��M ����)��M �T�� �)�	�M i�M `�+����M �t��M i�M ����+L�ҭ*� ��)� � ��L�� ��L�ҭ)��� ��L�� ��`�A ���A 8��A ����)`�M ���M 8��M ����*`�A �|��A i�A �� �)`�M �t��M i�M �� �*`�M 0�M i�M ��M 8�d�;0� <�`�M 8�x0L�ӽM ��L~��'�L~��9�L~��B�L~��N�L~��W�L~��`�L~��f�L~��o�	�A i�A �M i�M L�ӽA �8�L���@�L���H�L���P�L���X�L���`�L���l�L���t�L��Ɉ�L��ɘ�	�M i�M �A i�A �A ɰ��M 8�x0�'0 <�`�M 8�x0LaԽM ��LL��'�LL��9�LL��B�LL��N�LL��W�LL��`�LL��f�LL��o�	�A 8��A �M i�M L�ԽA �x�L���p�L���h�L���`�L���X�L���P�L���D�L���<�L���(�L����	�M i�M �A 8��A �A � ��M 8�x0�'0 <�`�M 0�M i�M ��M 8�d�;0� <�`�M ��	�M i�M `�M ���M 8��M � <�`�M ɠ��M i�M � <�`�M � �	�M i�M `�Y ,�M ʝM �A ʝA � ʝ �) ʝ) �5 ʝ5 �L<��Y `H� �t�� 8�� �� �� h`Hڭ ���L�֭ ���L�֩ �� � �3�������� �֭/���SL�ֽ5 8���M 8� 0�0L�֭ 8�M 0���) 

8���A 8� 0�0L�֭ 8�A 0��� ������dL��������SL�����	 SЭ	�#�?L�����
 SЭ
�<�+L����� SЭ�d�L����� SЭɖ�L�� [�A �'�M �( <խ8������� ��� � ��� � �/�	�Y �L���h`�� ��#� �@Lz��h0Lz׭ �20Lzש��/Lz���%� �DLz��h0Lz׽M i*�� �0�Lz׽5 8���M 8� 0�0Lz׭ 8�M 0���) 

8���A 8� 0�0Lz׭ 8�A 0�����/`H�Z� �� ��"������������
�� g�LZؽ5 8���M 8� 0�0LZح 8�M 0���) 

8���A 8� 0�0LZح 8�A 0��� [� <խ �� � �� ���� � � �05�������'�� i
 #�����X� �ȍ ��� � �	�Y �L��z�h``Hڢ �Y 0L�ؽ �
� ��L���� �L���� 4�L���� \�L���� ��L���� ��L���� ��L���� ��L���� ���Ll��h`H�� ��  �L���� p�L���� )�L���� �h`Hڢ �� � �轋 � �轋 � �Lm٢ ��� �\�[ ��g �� ��s ��� �D�[ �$�g �� ��s ��� �t�[ �$�g �� ��s �h`Hڢ �� � �轋 � �轋 � �轋 � �L&ڢ ��� �A i�[ �M i �g �� ��s ��� �A i�[ �M i �g �� ��s ��� �A �[ �M i�g �� ��s ��� ��� �A i�[ �M i�g �� ��s ��� �h`Hڢ �� � � 轋 � �轋 � �轋 � �轋 � �Lۢ ��� �A i�[ �M i2�g �� ��s ��� �A i�[ �M i�g �� ��s ��� ��� �A i�[ �M i�g �� ��s ��� ��� �A �[ �M �g �� ��s ��� ��� �A i,�[ �M �g �� ��s ��� �h`Hڢ �� � � 轋 � �轋 � �轋 � �轋 � �L�ۢ ��� �A i�[ �M i�g �� ��s ��� �A i�[ �M i�g �� ��s ��� �A i�[ �M i�g �� ��s ��� �A i�[ �M i�g �� ��s ��� ��� �A i�[ �M i�g �� ��s ��� �h`H�M � � �܀�h� ��h`H�M � � �܀�@� �܀�`� �܀ɀ� ��h`H�M �0� �܀�P� �܀�p� �܀ɐ� ��h`H�M �0!� �܀�<0�> �܀�d0�f ��h`H�M �0!� �܀�:0�< �܀�b0�d ��h`H�M �20�50L�ܽA �
�A 8�d�L ��h`�� � �L;ݽ �
� <�L;��� c�L;��� ��L;��� ��L;��� ��L;��� ��L;��� ��L;��� ��L;��� ��`�A i�[ �M i�g ��� �� ��s ��� `�A i�[ �M �g ��� �� ��s ��� `�A 8��[ �M �g ��� �� ��s ��� `�A i�[ �M i�g ��� �� ��s ��� `�A �[ �M i�g ��� �� � �s ��� `� �������A i�[ ��A �[ �M �g ��� ��s ��  /�`H� ��) 


��A 8� �� 8�A ��M 8� �� 8�M ��� ��+��6��A�L�ޭ�l��tL
߭�I��1L�ޭ�F��.L�ޭ�C��L�ީ�� Lߩ�� Lߩ�� Lߩ�� Lߩ�� Lߩ�� Lߩ�� Lߩ�� h`Hڢ �� � �L`��� ��L`��� ��L`��� ��L`��� ��L`��� ��L`��� ��	�L��h`Hڢ �� � �L���� ��L���� ��	�Lo��h`�g 0�g i�g ��g 8�d�;0� E�`�[ ɰ� E�	�[ i�[ `�[ �� E�	�[ 8��[ `�g 0�g i�g ��g 8�d�;0� E�`�g 0�g i�g ��g 8�d�;0� E�`H�� � �Ls��� ��Ls��� u�Ls��� ��Ls��� ��Ls��� ��Ls��� ��Ls��� ��Ls��� �h`�[ ɰ� �g 8�d�;�[ i�[ �g i�g � E�`�[ ɰ�#�g ��g 8�d0�[ i�[ �g 8��g � E�`�g ��g 8�d0�g 8��g � E�`�[ ��#�g ��g 8�d0�[ 8��[ �g 8��g � E�`�[ �� �g 8�d�;�[ 8��[ �g i�g � E�`� �g �[ �� � �s �� `H�Z�� ���C���� ���  ��� � ��$�'��(������m � ��� �� � z�h`Hڭ� ���1�(8��&� 0"�'��(������m � ���h`H� � ����h`H� � ���h`H�Z�� ���J� � ��$�� ��� ������m � ��� �� ���� � � � ���� z�h`Hڭ� ���1�� 8��&� 0"�� ��� ������m � ���h`H� � `���h`Z� x�� ��z`� ��� ��`H�Z�8�0Lb�
��G�� �G�� �� ��!����?�� ���� �JJ��0	��
��8�	�-�� i� � i � �!�!� �Ȁ�� � � ����!�L��z�h`H�Z�
����� 轃�� ��������?�� ���� �JJ��0	��
��8��-�� i� � i � ��� �Ȁ���� �����L��z�h`H�Z�%8�0L��"
��9�� �9�� �$� �#�!�&��&�?�� ���� �%JJ��0	��
��8�	�-�� i� � i � �!�!� �Ȁ�� � � ���#�!�L/�z�h`H�Z�8�0L6�
��7�� �7�� �� ��!����?�� ���� �JJ��0	��
��8�	�1-�� i� � i � �!�!� �Ȁ�� � � ����!�L��z�h`H������<0������h`H�Z����� ����
�����,�� �� � � i� � i � � G�� �ߩ��� L��
��� � � i� � i � � G�L���"���� � � i� � i � � G�(������� � � i� � i � � G�����  ]���  ]����z�h`� ��$�� �����	�����������8� i� �-� i� �0�
� ���'�� i
 #詂��  (�`H����� #���  ]���  ]�h`H� � f���h`H� � ����h`H�Z��� �� ��U� �� �� � �� ����z�h`H��� �� U� �� ��U� U� �� �� �� � U� ����h`H�Z� �@� � � �-����� ���z�h`H�Z�/���� ���� ��z�h`H�Z����� ���� ��z�h`�  ����`Hڪ�.�




���)�& �h`H�Z ��
��1�� �1�� � � �@� � � ����(��� i0� � i � � i(� � i � ���Ωύ& z�h`H�Z
������ ����� � ���$��a��[��d��*�8�7��  z�Ȁ�z�h`H�Z�)�JJJJ��  z�)��  z�z�h`H�Z� H� H� H� H�� �[��$��a��%��d��&��*��'����� ���� ����?�� ���� ��� ��R�� ȱR���-�� Ȳ-�� ��н��h� h� h� h� z�h`� �� �� ��  �� �� � � � � � � � �* �� �� � ���� �� `�� ���%�� � ��� � �� �  ���� �� �� � �꭯ ���%�� � ��� � �� �  X��� �� �� � 뭭 ���X�� ����� � �� � �� �  )쭯 ����� � ��� � �� �  ��� �� ͵ � #��� �� �� � z�� ��� �� K�`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
������ ����� �� )0�� ȱ������ Ȍ� �� �� �� � �L물  ��� ��� � ��� ��Ȍ� �� ���� �͍� ȱ͍� ȱ͍� ȱ͍� ȱ͍� )
������ ����� �� )0�� ȱ������ Ȍ� �� �� �� � �� �� � �� )������ ��  �`�� �ڍ� ȱڍ� ȱڍ� ȱڍ� ȱڍ� )
������ ����� �� )0�� ȱ������ Ȍ� �� �� �� � Ы� �� � �� )��@К���� ��  �ꀍ�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
������ ����� �� )0�� ȱ������ Ȍ� �� �� �� � Ъ��  �� ��� � ��� ��Ȍ� �� ���� 
������ ����� ���� ȱ��� `�� 
������ ����� ���� ȱ��� `H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����λ �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� �ƪ�� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� �Ԫ�� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� �᪭� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� � z�h`� `� `H�Z�� ���%�� ���� �� �� )?
������ ����� ��  �z�h`�� �* �� `�� ���� ȱ��� ȱ��� ȱ��� )
������ ����� �� )0�� Ȍ� �� �� �� � ��� `H�Z�� ���L��� �� �� I�� )��� �� �몭� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� )�� �� )����
�@����� �� �� �( �� �� ��* �� �� �� �� � �z�h`H�Z�  ��  윰 �� ��� ��  #� z� )� �� ����� z�h`H�Z�� � �
�� � ��� �� )?�� �Q�� �K�� 
������ ����� ����� ����� �� �� � �� �� �� )������  �� ����  �� ��z�h` ���� ���� ���� ���� ���� ��� ���� �G�� ���� ���� ���� ���� ���� ��� ���� ���� �(��� q���� K��� d��� q��� ���� q��� ���� ����� T��� K���� C��� K��� T��� q��� T��� C���     � K�� ���� ���� �������.���� ���� ���� ����.��� �(��� ⠧�� ���� ���� ���� ⠧��.���T����     � ��� ���� ���� ���� �
��� �槕� K��� C��� K��� Y��� ���� ���� ���� ����.������.���h������.��� �������.���h���T���@���     �.x��� ���� ���� ����.��� ����  �� �
��� 
 �� �
��� 
 �� �
�� 
 � �
�� 
 �
�� 
 � �
�� 
 � Y��  � Y
�� 
 � Y
�� 
 � q
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � ���  � �
�� 
 � �
�� 
 �     � �
�� 
 � �
�� 
 �
�� 
 � �
�� 
 � Y��  � Y
�� 
 � Y
�� 
 � q
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � ��� ��� ��� ��� ���.�� ��� ��� K���     ���   ��
�� 
 ��
�� 
 ��
�  
 �O
�� 
 �?
�� 
 ��
�� 
 �h�  �h
�� 
 �h
�� 
 ��
� 
 �
�� 
 ��
�� 
 �
�� 
 �     � �
�� 
 � �
�� 
 � �
�� 
 � q
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � q
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � q
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � �
�� 
 � q(��     ��
�  
 ��
�� 
 �\
�� 
 ��
�� 
 �\
� 
 ��
�� 
 ��
�� 
 ��
�� 
 �\
�  
 ��
�� 
 �\
�� 
 ��
�� 
 ��
� 
 ��
�� 
 �\
�� 
 ��
�� 
 �\
�  
 ��
�� 
 ��
�� 
 �O
�� 
 ��(�      � ��� /d��     � �� � �� � �� � �� � �� � �� � �� � �� � �� � �� �� �� �.� �     �     � � � �} � �| � { � _z � Ky � ?x � �w � �v � �u � t � _s � Kr � ?q �     � � � �} � �| � { � _z � Ky � ?x � �w � �v � �u � t � _s � Kr � ?q �     ����%�  �O   �O  % �     % �d  % �    �    � �
	 �
�



	�	

			
�
	
	 �

		�����������g���{�k�  +�  ��  ��  ��7�=�������,�/�7�F�P�������PRESSaSTARTaKEY$$SCORE$7777777$READY$GAMEaaOVER$STAGEaa8$STAGEaa9$STAGEaa:$STAGEaa;$PAUSE$7$8$9$:$;$<$=$>$?$@$*a:$dddddddddddddd$SCOREaa7777777$PROGRAM$ESONaCHU$MUSIC$L[W[aXAO$PICTURE$Y[aBAN$L[aZHANG$CONGRADULATION$CONTINUE$���#�+�1�<�E�N�W�`�f�h�j�l�n�p�r�t�v�x�~�z��������������������� � @ �ȸp���X���跈�	�I�p���ɬ	�I�����(���˭��C����p������˭��˭��H���ȶ�Ժ:���I���ɕ	�I���ɖ	�I���ɗ	�I���ɘ	�I���ə	�I���ɚ	�I���ɛ	�I���ɜ	�I���ɝ	�I���ɞ	�I���ɟ	�I���ɠ	�I���ɡ	�I���ɢ	�I���ɣ	�I���ɤ	�I���ɥ	�I���ɦ	�I���ɧ	�I���ɨ	�I���ɩ	�I���ɪ	�I���ɫ ��� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       a� ���