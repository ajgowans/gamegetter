�m ���v �/�� ��r ��t ��u ��e ���f �f �l �e �k  �ۭf �r� ��f �u ����u �� �� ��� ���� ��� �f �f �l �e �k ��r ��u ��t  ��Λ Λ �� �l �� �k �� �u ��r ��t  �ۭ� �D� ⭳ �� � ����� �� � �f �l ��u �e �k ��r ��u ��t  ܭe i�e �k  �۩�u �� 8��� �k ��r ��t  �ۭ� ��  ���^  T�< ���L�                  ��m  ���t ��u ��r ��k ��l  �۩�r ��k �(�l  �۩L�l ��k �!�t �=�u ��r  �۩��l ��k ��t ��u ��r  �ۭ  ��� �v � �m L �                                                                                                                                                                                                                                                                                                             H� �v � �� ���f�� � �� ��Y� �  � �� �� ��P�q ��p � 㭊 �s �P�q ��p  p�
�� ���w �w � �  ��� � �� �� K�h�v L���  ��00  ��?�?������0  0030  �������� ��  00�0  �������� 3�  �33  ��?��������?3�  003<  ���� ���� ��  0030  ��0�� ��� 0  ��00  �������?���                                                                         �  � � �            �                �                 �  � �              �      �             �      0             � �  �  �       ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?   ?��������?�?   ?����������?   ?��� ����?   ?��� ����?   ?��� ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                                  �   �     �� �? �?   � �U� p��  �WU \� p� �UWUU� \UU� �_UU W� \U �UWUUU\UUU\UUU WU\U �UWUUU5WUUU5\UUU WU\U5 �U\UUU�WUUU�\UUU \UpU5 pU\UUUUUU�W�\U��  \U�U5 pUpU�WUUU\�pU?   WU�U� \U�U\U_� \���    WU�U� \U�� pUs� W���� �UU5�U� WU�� pUs��U5|UU �U_5pUUWU�� pUsUU5WUU p�\5pUU�UU�� pUsUUUWUU p�p�pUU}UU�� \�pUU�WUU _��pUUUUU�� \�pUU= |�� �UUU�pUWUUU�� W�pUW5 p5  �UUU�p�\U�U���U�p�\� p5   WUUUs�pU5W�UU5p�pU?p����UUUUs5pUW|UUU5p�pU�\UUU�UUUUs5�UW\UUUp��UUWUUU}U�U}5 � W\UUUp� WUUUUUU� �UU5 < W\UU� p5 \�WUU�W�  WU5   WpUU= � p5|UU=\5  W}   ����    �����  ��   <         �   �    �  �   ��  ?�W  W��  p5 �W�?  p\5 �5pU��UUU p5 \UU� \5\� ��\UU=�UUU� p5 \UUU= W5\� �UWUU��UUUUp5 \UUU� W5pUpUUUUU}UUUUp5 pUUUUW�pUpuUUUUUUUUp5 pUUUU\�pUp�UUUUUU��Up5 �U�_UpU�U\�UU�U�U�U\5  W=pUpU�U\�U�W5WpU\5  W�UpU�U5W�U \5W\U\  W�U�UW�U�U \5W�WU\  W�U�UWUU�U \5WUU� \  W�U W�UU� W \5WUU= W  WpU WUUU� W W5WU� W  WpU WUUU� W W5WuU W  W\U \UUU5 W5�U5W�U W  WWU \U}U5 W�UWW�W�� W�U�  \UsU5 \UUUWWU�WUU�UUU�  pU�U \UUUW\UuUUUUUUU5  p��U pUUUWpUUUUUuUUU  �� W �UU� W�U}UUU}UUU  �� W  _U= �  W�WU��UU�    � �  ��    � �� ��                UU                            @UUjUU                           UU��UU                         PUU��UUU                        UUU��VUU                       @UUU��VUUU                       PUUU��VUUU                      UUUU��VUUU              $     @UUUU��VUUUU                  0 PUUUU��VUUUU      �          @=TU�ZU��VUUUU                  � UU�jU��ZUUUU                   @UU�kU��ZUUUUU                  PUU�kU��j�UUUU                  PUU�kU��j�VUUU                  TUU���:?��VUUU                  TUU�������VUUU           0      UUUꯦ�?��VUUUU   0       �      UU�ꬪ� ��VUUUU   �             @UU�����?���ZUUU               @UU��̪����jUU�                PUU�>���ϯ��kUUU                PUU�����Ͽ�jUUU             �  TUU��������kUUU             0 TUU��?�����UUU             �  UUUU��������VUUU                UUUU��?3��?̯ZUUU                UUU������3�jUUU               @UUU�������jUUU              @UUU��0���� kUUU          �   @UUU��?<���33kUUU          �  PUUU�������?���UUU          0  PUUU��?���?���UUU              PUU��������? �UUU�             PUU��� ��? �UUU              TUU��� ���̬UUU              TUU��� ��0̬UUU             TUU��� ��0̬VUU              TUU��� �?0 �VUU              TUU���?����� �VUU           �  UUU����3 �����VUUU           � UUU����3 ����VUUU           �  UUU���?��������ZUUU              UUU����� �?��jUUU              UUU�?�����?����UUU              UUU�3�����?���VUU              UUU�3�����?��3�ZUU              UUU�3?��  ?�3�ZUU              UUU�<��  ?�����ZUU             UU�� ���  ?�<��ZUU              UU�� ���  ?�<��ZUU              UU�� ���� ?�<��ZUU             0UU�� ����?�<��ZUU              UU�� ����?�<ϼZUU              UU�� ����?�<��ZUU              UU�� ����?�<��ZUU             UU��������������ZUU       ���������������������������������           �����������                       TUUUUUUUU                         UUUUUUU                         @UUUUU            @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            H�Z ��2�� �� �� �� �� �� �� �� ��� �� ���� �� �� ��� �� ����� �� �� ��� ��	���#�� �2�� �g �� ��� �������  3ة�n ��o �� 

m� 
��<�h ȹ<�i  �ޥ �Z  !��k ���l ��r ��t ��u  �۩�k ��r  �� -� Cǩ��q �"�p  �ǩ��q �"�p  �z�h` � ��? ��? �� � � ��������� � ��  �  ���<�?̫�<�� �� 3 ��� �?�����  � ��? ��? �� � � ��������� � ��  �  �3  �0  ?0   � ; ���   �0 ��� ��? ��  � ��? ��? �� � � ��������� � ��  �  �� ��� ���  ��  �0  �  3    �  �  �  ��  �� �3 �0 3 ������0�?  ��  ?0  ��  �? �? ��  �  ��  ��  00  �  �  �?  ��  �� �3 �0 3 ������0�?  ��  ?0  ��  �  �  00  �  �� 0�  � �33 ��? �� ��  �� �3 �0 3 ������0�?  ��  ?0 ��� ���0�?<��30��<���  ��  ����� ?�? ��  �� �3 �0 3 ������0�?  ��� ��� ���������� ��� ��� �� < < ���?����? � ��? ��? �� � � ��������� �?�� �� 3�� ��� � ������� 00< 0<0 ��� ����                                  �� �VU�V `UP�V U jU� ���  �*                                �    �  @ UU	 U�
 �� �
                         �   X  �Z  XU �ZU��U�UUUjUUU�ZUU hUY ���  ��  �� �* �  U(TUUUUUUUU UU UU         UU  UUUUU�UU���j�  �*  ���
   �
UU�UUU��U PUZ @U�  P�  PU PUUPUUUUUUUUU��U�������� �              �   
  V   Z�  i� i� i� i� j�  Z*  �
  *                ��
 jU)�U $h@�VUU��VU) ��
 ��                                       �� �* � P(PUUJUUUVUUUjUUU�VUU���� ���                ��  
   � PU UUUUU)UUU*UU�
U����� ��  �          ����W�W�W�W�էէ٧٧ڧڧ����?�?����W�W�W�W�էէ٧٧ڧڧ����?�?  ��  W�  W�  ��  ��  ��  ��  �?����W�W�W�W�էէ٧٧ڧڧ����?�?�����_�W�W��z��z��Wz��W~��U^��^���^�z�^�z�_�~�_�~�_��W���W���<��<�<<�������������<��<�<<�<��<�<<��?�<��<��?<���<��< �?<      <�  <� �� <�  <  <  <�  <<  �<  <<  <<  <�       �?�<��<��<�����<�?< �  � �� ��Q�`Ռ1 �\�*���  ������t��{'" � 0z@�  @       � �_5<p�;p���sհp���_��^U��W�5;W�5W}5�_U�0����0 � ? ?          � �_5 <p� p� �p��pի�_��^U��W�5 W57 W�7 \5 �� �� �?<�_���z�ð��<��� ��> ��: ��: �*2 �"2  0 �   � � �� ��      � �_= �z����?���ü�>ë�:<��: �*2 0"2 � 0 � �� ��  �                                 ����W�W�W�W�էէ٧٧ڧڧ����?�?����UU�U��ꩪ�ꩪ������UWUU����������������UU�U��ꩪ�ꩪ�ꩪ�� <� �p5 Ws5 \_ \W<�� ��� ��?�w��w������                         �? ?p����U_� �U5<�W��� ��?�w���w������                            ��          ܰ         ;p        ��         ���         _�9        ���        �oU        \�U        �B�        ��T�        p���        ���        p�=         pe�         \Y�         [Y�        [W�        [We=        [We��       l]eUU�      �]�UU�     �]�UUU>     �W]U�Z�     {�WU�j�    _}UUm��    �oUU[U�   �5�UU[U�7   �5�j�VU�7    � ��UU�7    < �UU�5      p�UU�9      p�UU�:      p�V�}      ��W�o      ��_��       �_l       �_l       �_�       �_�        �_�        �_�        �_�      ���W9�     |�_U9l�    WUU�:��-   ��������   �         ��         p�        ��       ��U�       \Օ�        i5        �Ue�        �_Z�        ��[�          \U         pU         pU         �i9         ��9         �U�         �U�         pUY        pUY=        pUV�        �UWU       ��UU�       �]UUU�      {]UUUU     {sUUU_=     |�UUժ� �   p}WU�V���  ��[U�UU��5   ?lU�UU]��    �U�UUu��    �V�UUu��     [�UU��     �UWU5 �     ��WU9 �      �WU �      �_U ;      �U ;      ��U 7       �W5 7       �_��:       ��U�       �W�       p\�       \\�        � ׀       ���5        �>|         ��                �         p?         �7         ��        ���        \��        _i�        ��V5     �> ��Z5     ��p)d5  �?  p\Je5 �U� �9�WZ UU=  7�W=�UUU� 7�W�WUUUU �  WUUUUUU �  \eUUUUU5 �  \YU�UUU5 �  \YUUW�_� �  �YUU]�����   _UU]]U��   p�U]WU�e9   �ZU_WUU�9   �W��WUU�   �U��WU��  �~� �UU�   �Z �UU9     _? �U�     |� �W�      �? �W9         �W         �W         ��        ���         ���         W�9        ��p        �|          W         ��          p5          �?         ��                                                                                                                                                                                                                                                                     � ��       �� _U�      ������    �����V    �@����<   ?����*�  ��U���(� ��PU��k  � � UU��k  T 0UU��f �> �R�V A�� O�o�S� U�����Z>��� ���������U���胫���U���C���CU������_���Ce������_���_�����������������>���������>  0�������j  <�������Z  <�?�?����7  �������?  ��ç� ���  �� �� ��� ��> �� ���� ��? ��  ��� 0� �� ���� �� �> �[������W? _��?��� �� ��?                                                                                                                                                                 �          �� �?      p���W�      ��K��    �@��T�    @�kT@�;   �@��V��   0@��U�B�  P	�kU�N�  �9T
@�:�  e:�
���? �C��#���� �P��Z���W�����Z�Z�V����UZ�Z�Z�L��@�n�j���L��U�n�*���<T�V�n�������Z�n�������Z��O���S�����C��������P���K����T��� �����U��� � ���� ����   ���U���  ������  ��?���?��  |������>  |� W����  p� \����  p� ����� �� |� �� ��  _�? �� ��?  ��? ��                                                                                                              ��         ��        �_�       ��_�       � ��       �Wi�      pU���      �*P?     ���zP�      ��Ao�       ���o       ��kU       ��Z�=       ��V��      ���n�      ��U�      ��U�<     ��T�V�     ��T�V    ���V    ��A�U    ��VT�E0    ��WE)@0    ��[E)@�    ��_Ai@@   ��oI�@�   ���I�E�   ���K�D�5    ��K�V�5    ��Z���U5    ��Z��U5    ��R��oU5    ��R���T5    ��T���j9    뿔����>    �o�����   ��[5 ���   ��U?�oU�    ������        �         �          �   �    ��      �>�:   0    3�:   �   ���:   �0   ���   ��   L���  ��   �_�[9      W�S�   <  ���C�   � ���@�   ����@�  0 ���:�C�?  �  �N�S�?    �:��R��   <   �����   �  �=���    �? �O���    ���S���      �U���     �WU���     �UU���     _U����    �WU�W��   ��U�_U��?   �W��SP��?  �WU� P��>  �U� P��;  pU�  @�O;  \�  <@�@;  �   <�>T;  ?   <�C�:       �� �:       �?P�:       �ի:       ���       ,��       ,>��       �:U�       ��_�       �?�      ��|�>      ����      ��\U�     ����W��     �������       �         �          �        ��        �>�:         3�:        ���:        ���        ��       L]�K9       �W��       ����       ���
�      ���J�      08�K�?      0N�W�?      0��V��      �����      �����      ������     ������     ��n���   ����[��   < ��W��   ���W�U�  ������V�  ��UU�>T�?  ��WUU�T�? ��Uk��U�>   �U�����;   p���C�O;   p�  @�@;   p?  P?T;   �3  .��:   �  ��@�:   �   �?U�:       �O�:       ����       ����       ����        ���:        ���        �_�        ���       ��_�       �{U�       ����        ���        �         �0         �2         ?�:         ���         ���        �j�        ��j�       �[��?       0U�.�       ���      �W�/�       ��+�       �_+�      ��T/�?      �8�_��      �8�[��      0�[��     0L���     0��V��     0��V��     0z�U��     0z���?     z��o�?     �m�W�>     ��m�[�>     ��]�P�>     �:_:P�>    ��>�>T��    ��>�T��    ����?�    �����    ����K�P�    ����T�    �������    �����T��    ��p�?���    ��p���:    �������    �������     ������      ����:      ����      ��>��      �z>�       ��U�        �^�        ��� � 0� 0�������z�k��Z���>����Z��k���z0����� 0     0�* �Ⱦ(�# �����<+8��:,8JU�,8Z �,� �� �bD �� ��X %�HU!����.�(0. �<�0� ��
 �2     �~������W��_��^{��^{��z{��z{�W{�^{y��_y��^{��~y��z���z{��z[��~�������W�-�_�/�^{��^{��z{��z��W{��^{������.�3�0   �~������W��_��^{�0^{�0z{���{������y�� {� 0�� 0� 0 � 0�� 0��                                ��j�Vj��iY�i��Z���j�YUjY��Y�Z��j��j�Vj��iY�i��Z���j�YUjY��Y�Z��j                                            3333��������UWUU����������������UU�U��ꩪ�ꩪ�ꩪ�ꩨ��*  ��*(�bUU�ZUU�ZUU�ZUU�VUU�VUU�VUU�VUU�VUU�VUU�ZUU��j������(UU	(UU	 UU
�TU�T��P� �R� �R�  B%  J)  J	  H	  h
     �  �    ��  �  ��  j�  V�  V�  ��  �*��  �  *�  V�  V�  V�  ��  �*  ��  �  ��  V�  V�  Z�  ��  ��    ��  �  ��  Z�  V�  V�  �*  �
��������[UU囙��[f��[����[������[������[�������������������  ��  W�  ��  ��  ��  ��  ��  ����  ��  [�  ��  [�  ��  ��  ��  ��  _�  �  ��  ��  ��  ��  ��    ��  ��  _�  o�  ��  ��  ��  ��                                  �  ?30�� ��  [ �V��P�Z����?����P�UO�C�O�S�C��S����>�S�??����O�S�S�S�W������?��  �?  �  �  C�  C�  C�  S�  �>���� � S� S� �� ��  �?  �  0  �  [�  [�  k�  ��  �:  ��? �� �V� �Z� ��� ���  ��  �??��� �* �V�`T	 U%|}%F��֪��֪��֪��V��V�z�X�^%X�W%`UU	�V� �*  �* �V�`T	X U%S�%�w�V�^�V�{�V�{�V�^�V�w�XW�%XUU%`UU	�V� �*  �* �V�`Uu	Xu}%X_s%VsÕ�pÝ�� ��  ��  �V �X�%X�)`UU	�V� �*                     �  � �����_��0_w� \w? �w �� 0� �3 ��<                        �  � �����_��0_w� \w? �w ��  �  �     �=  _��UUpu}6��s�W=|�gp�WUU�W�W�gU��W�W=W5�;�����  �   �   | �W� pUU�}]W�{6g=|�WpٗUU�g՗�WVU�|՗���\���?  �:  ��         �? �� �����p�����WUu�WUU�W�U�\uW��_U�pUU��W�� �? �� �? �� �����p�����WUu�WUU��_U� �U� pU��_U��W�� �?  �  �  �?                                                                  	         �   �      �   �                                            � 	                 � �       �                                         � 	                           �      �                                  � 	   �              
      
      
    �

     

     
      
     
   	   
      
     

     


  �                                                             �          �                       �                        �    �      �                                ��          ��           �                      �                            �        �                                            �          �                                                                      �      �      �                     �     �        �   �     �                   �        �           �                                 �    �                                    �     �     �   �     �                               �            �                 �              �       �      �             �                        � �    � �                                  �      �      �            �                       �                               �        �   �       �                                                                  ��         �                                                                     �       �                                                                                    �     �     �  �                                �     �     �                    �     �  �   �  �      �                                                                �                                                    �     �   �         �     �     �       �                   �     �   � �             �     � �   �   �     �                    �     �     � �       �     �                                �     �     � �       �     �                          �     � �   �   �                          �     �     �                 �      � �         �                        �                                 �       �          �                                �                �                                                                         �  �   �  �    �      �                  � �    � �           �        �    �       �  �      �           �      �            �      �         � �     �         �        ��                                      �     �                                           �    �                  �  �        �                        �   �     �          �         �    �       �          	   �                                                                      �      �      �  �      �      �                ��     �     �    �                                �                     �    �       �                �                �                   �      �                   �        �   � � � �      �     �     �  �    �     �     �     �  � � �      �     �     �  �    �     �     �     �  � � �      �     �     �  �    �     �     �     �  � � �      �     �     �  �    �     �     �     �  � � �      �     �     �  �    �      �                                               	        �   �              �     �   �             	  �              �                                  	       �                                �                      	   �   �                      �                                    � 	                                                         �    	     �                                                                                       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���ة��  ��� �� � ��� � �ύ& ��" � t ����� ��� �� � ������ ��� ��XL �H�Z� �� �Έ (z�h@H�Z�' )��d ��� w� w�� �� �# �$ �% (z�hX@                                                                                                                                                                                                                                                                                                                                                                                ���~  9�d�� �# � U�L �� U�LP�� U✬ �� �� �� �� �� ��� � �� ���� ��� �n�� �7�� �7�� �� �� �� �� L��  � �� [� �� Y� �� %� �� k� �� ǜj �� 

m� � �L���L#���LI���Le���L}���L����L����L����L���	�L��
�L;���LW���Lx���L����L��L�ĭ� �'0�� �#0Ll©�� ��� �� L�ĭ� �0Ll­� �ZLl©'�� �n�� ��� L�ĭ� �0Ll©�� �n�� ��� L�ĭ�Ll©�� �.�� �� L�ĭ� �'0�� �0Ll©�� ��� ��� L�ĭ� �'0�� �ZLl©�� ��� ��� L�ĭ� �&Ll©'�� ��� ��� L�ĭ�Ll©�� �.�� �� L�ĭ� ��� �10Ll©�� ��� �� L�ĭg �+��� �pLl©�� ��� ��� L�ĭ� �'Ll©�� ��� ��� L�ĭ� �'��Ll©�� �>�� � �� L�ĭ� �'Ll©�� �.�� � �� L�ĭg ���� �pLl©�� �n�� � �� L�ĭ� �'Ll©�� �n�� � �� L�ĭ� �'Ll� ��L<�L© U�L �� U�Li�H�Z� �  � �� �� �v �� �� ��  ��2�q ��p � 㭌 �)�
�� ��y ���w �w � �  ��� ��y ��LƩZ�q ��p � �[�q � �p  �ǩd�q ��p � �e�q � �p  ȩx�q ��p � 㩂�q ��p � �x�l ��k ��t ��u ��r  �ۭ  ��_ �l �x�?�v �� �z�hL������.�����.���>� �� �� Ί ��� Ό z�hLP� 9�d�� �# ���v z�hL�������В � �~  �۩��~ �l �x��x����l  ��L��Hڮ  ��  9�d�� �# � U⩀�v  ✂ �hL	� �Ɗ	� �Ɗ	� �Ɗ	� �Ɗ	� �Ɗ	� �Ɗ	 �Ɗ	� �������� �ة`��  �0��  ��h`��� dـ@����:��� -ـ1��� ـ(��� =݀��� dـ�� H�ɿ� �ހ��� `H�� � ��h ��h`H�� �� ���l �
�k  Y�h`H�� �� ���l �
�k  Y�h`H�Z�l ��w �x N� .x N� .x ��y �� �z ����� ���mv �� �k �� �������y �z �z ��x �� ������x �����?����y �y �� ������w �w Еz�h`H�� �s  p⭪ �s  p⭩ �s  p⭨ �s  p�s  p�h`H�� �s  p⭮ �s  p⭭ �s  p⭬ �s  p�s  p�h`H�� �
6m� �� �
008�
�� � �� �
0 8�
�� � �� �
08�
�� � �� �٭� ͯ 07��� �� �� �� �� �� �� ��� ͮ 0�孩 ͭ 0�᭨ ͬ 0�ݩ��q �"�p  �ǩ��q �"�p  �h`H�� 
i�r �� ���r ��t ��u �� �k �� �l  ��h`H�� i͗ �� �~  �ȩ��~ h`H�� ��� i��� �w ��� �� ��O�w ͚ �L�ɭ� i�w ��� �w ��w �W�� ��� i$��� i͘ �=�� iʹ �2�� �-�� ��&�� �w ��w i͚ 𼭗 �w ��w i͗ ��h`H�� �1�� �,�� �� �� ��  %ɭ� �� �̜� �� �� �Z�� �L�̭� �1�� �,�� �� �� ��  %ɭ� �� �̜� �� �� �Z�� �L�̭� �.�� �)�� �� �� ��  %ɭ� �� �̜� �� �Z�� �L�̭� �1�� �,�� �� �� ��  %ɭ� �� �̜� �� �� �Z�� �L�̭� �.�� �)�� �� �� ��  %ɭ� �� �̜� �� �Z�� �L�̭� �1�� �,�� �� �� ��  %ɭ� �� �̜� �� �� �Z�� �L�̭� �/�� �*�� �� �� ��  %ɭ� �L8� �̜� �� �Z�� �L�̭� �/�� �*�� �� �� ��  %ɭ� �Ll� �̜� ��Z�� �L�̭� �/��*��� ���  %ɭ� �L�� �̜�	�Z��L�̭�F��� ���  %ɭ� �L�������| ��}  %֜���d ��X  �� �֩
L�̭�F�� ��?��� �T��  %ɭ� �L�������| �T�}  %֜���d ��X  ��
L�̭�g�� ��`��� ���  %ɭ� �L�������| ��}  %֜���d ��X  �� �֩
L�̍�  <� =کc�� ��  
ɜ� �� h`H�� �k �� �l ��t ��u ��r  �۩���  � ܩ��d ��X  ��h`H�� �k �� �l ��t ��u ��r  �۩���  � � �~  �۩��~ ���d ��X  ��h`H�� �k �� �l ��t ��u ��r  �۩���  � �~  �۩��~ ���d ��X  ��h`H�� i͛ 0F�� iʹ 0;�� iͳ 00�� i͚ 0%�� i͚  x֭� 8��� � x֭� i�� h`H�Z�� ��q�� ��%��� �g �_�(��Y�� �g �Q� �M�#��&�#�$��L9���L����L����LD���LU���Ll��
�LD���L����L��z�h`�� �*�� ��g �� �L5έg �� �� �f i�� ��� L5έ� �L5έg �� �L5΍� �� �f i�� ��� L5έ� �*�� ��g �� �L5έg �� �� �f i�� ��� L5έ� �L5έg �� �L5΍� �� �f i�� ��� L5έ� �*�� ��g �� �L5έg �� �� �f i�� ��� L5έ� �L5έg �� �L5΍� �� �f i�� ��� L5Ύ�f ���L5έ� ���� ��� �\�� L5έ� �/���g ��L5έg � �� �f i�� ��� ��L5έ�L5έg � �L5΍��f i�����L5Ω�L5Ω��T�����L5�H�� � QЭ� � sЭ� � �Э� � �Э� � �Э� � �Э� �ԭ� � ѭ� � aѭ� �ѭ� \խ� ��h`Hڢ �� �� ���� �Ѣ �� �� �����h`Hڢ �� �� ���� �Ѣ �� �� �����h`Hڢ �� �� ���� (Ң �� �� �����h`Hڢ �� �� ���� (Ң �� �� �����h`Hڢ �� �� ���� &Ӣ �� �� �����h`Hڢ �� �� ���� &Ӣ �� �� �����h`Hڢ �� �� ���� �Ӣ �� �� �����h`Hڢ �� �� ���� �Ӣ �� �� �����h`Hڢ �� �� ����  Ԣ �� �� �����h`Hڢ ��� ����  Ԣ �� ������h`H�� ��	��� ����� ��r  x� �׭� � �� i
�q �� �p �p �p  +ܭ� �� �g 8� 

�w �n m� 8�w � ���(���  \� �׀ x֜� �� �2�� h`H�� ��	��� �!���� � �r  x� �׭� �g��y �� �t�2i�q �� �p �p �p �p ��z �p  +ܭ� ��z ��� �y �ǭ� �q ��w �� �p �p  +ܭ� ��q �w ��� �1�� i�p ��y ��w �� �q  +ܭ� ��q �w ��ι �y �ݭg 8� 

�w �n m� 8�w � �� �� ���(� \� �׀ x֜� �� �2�� h`H�� ��	��� �#���� �"�r  x� �׭� � �� i�q �� �p �p �p  +ܭ� �� �g 8� 

�w �n m� 8�w � ���(���  \� �׀ x֜� �� �2�� h`H�� ��	��� �*���� �)�r  x�� � �� �$���� �� ��
��� �
�w �L8�w �� ��  \� ��h`H�� ��	��� �,���� �+�r  x֭g 8� 

�w �n m� 8�w m� �� � �L���(�L�ԍ� �� i�q �z �z ���� mz �p  +ܭ� ��z ����� �8�� 8��q �z �z ���� mz �p  +ܭ� ��z ���� ��� �0� m� ��  \� �׀ x֜� �� �2�� h`H �֭��	���'�!��	���(���	���'����&�r �8���\��ȹ\�Ș8���2���� ����� ���  �֩@��  � ��h`H���	���.�!��	���/���	���.����-�r ��� ��T�� � �֩@��  � ��h`H �֭��	���1�!��	���2���	���1����0�r �������������m��� ���  �֩@��  � ��h`H 
� Uؠ  Uع��m| �� ȹ���m} 8���  �� #� 3��0� ��h`H�� �k �� �l ��t ��u  ��h`H� �~  \֩��~ h`H�� �k �� �l ��t �0�u  ��h`H� �~  �֩��~ h`Hڭ� �� �� �� ���� \֭� �� �� �� ���� \֭� �� �� �� ���� \֭� �� �� �� ���� \֭� �� �� �� ���� \֭� �� �� �� ���� \֭� �� �� �� ���� \֭� �� �� �� ���� \֭� �� �� �� ���� \֭�� ��� ���� \��h`H�� ��� i0��� i͛ 0<�� iʹ 01�� iͳ 0&�� ��� i��� i͚ 0Τ  Cǭ� �o0Τ  C�h`H�� �� i ͛ �+�� iʹ � �� i͚ ��� iͳ �
��� �ι h`H��t ��u �� �l �� �k �� �r  ��h`H�Z��y ��z �� ����� ��� �� � ����y �y ��t �y ��z �z ��z�h`H�� ��� ����� ��� �0��� ��  3�h`H�� ��� ������ ��� ���� �Μ  3�h`H�� ��� ������  3�h`H�� �� �� �ܭ� ��� �� �؀���  3�h`H�� �� � �ܭ� ��� � �� �؀���  3�h`H�� � d�h`HZ Uح� ������ �� �� ��� � Ξ �4Λ  �ܭ� ����� � Λ � Ξ � �ܭ� �� �ٜ� �� �� �� �
����  3� 7�zh`HZ�� �G Uة
�� ��� �� ��  �ܭ� �
� Ξ �� �� �߀�� ��� ��  3؜� zh`�  ���)���� =�`H�#�&��"�� 8�� �!�� �"�g ��#:i�#h`H�#��2 {ۭg 8�

�w �n m 8�w �!�!��$��# {ۀ U�h`H�#�Y�"i͛ �N�� i�"�C�!i͚ �8�� i�!�- {ۭ#�� ۀ�� (ۀ	�� Eۀ �!�"�# �� 3�h`H�� i�70�7��  Cǩ
��  <�h`H�� i
�70�7��  -ǩ
��  <�h`H��� �
��  <�h`H�#���r �!�k �"�l ��t ��u  ��h`H� �~  U۩��~ h`H�Z�r 
��� 轴�mv �� �t �y �u �z �l ����� ��� �k �0*�+&�m ���-~ �����������I����Q����� i�� �� i �� ��y �y и�t �y ��z �z Кz�h`� �~  �۩��~ `�ZH�q ����� ��� �p ���� hz�`H��w �� i�p �w �w ��� i8�w �q  +ܭ� ��w �� h`H��w �� �p �p �� i8�w �q �w �w � � +ܭ� ��w �� h`H��w ��y �z �� i�q �� mw �p  +ܭ� �	�z y �z y �w �w ڭz �� h`H��w ��y �z �� �q �q �� mw �p  +ܭ� �	�z y �z y �w �w ڭz �� h`H�� �a��� �� 
i�� �� �0!���  3ح� i�� �� i�� ��� �� ��  3ح� �� � �� i�� ��� � �^  T� #�h`H� �ɭ� ��N�j � 
ɭ� �p �p �p �p  ޭ� �!�p  ޭ� �� � �  ��� �� �� 
ɩ2�� �� �� �h`H�w �� mw �q  +ܭ� �
�w �w ���h`H� �ɭ� ��Q�j � 
ɭ� �p �p �p  ޭ� �,�p  ޭ� �!�p  ޭ� �Η Η Η  ��� �� ��	�� ��  
��h`H�� �!�� ͔ ��� �� �� 8��� �  -� �h`H�Z ��e �f �w � �e �� �	�e ��(�H�� ��	�� �<��8�g �3�h/�y )�$Ny Ny Ny Ny �y )�&Ny Ny �y )�% �̀ �h�0�r �n me �k �o mf �l  ����w �w �c��f i�f ɐ�L�ޭe i�e �f L�� �h������ ��� �g ��  ��z�h`Hڭ� � Iܭ� �q U�� ���� �g�� ��A Iܭ� �U�n ��j  �ޭn �H��n �g �g ͱ 0�� �h i	�h �i i �i �� ��� �' Iܭ� � U�� ���� � U� 3� ��h`Hڭ� �0 }ܭ� �L�� U�Κ ���� �l }ܭ� �a�n �00�g �09��n �g �g Ͳ ��� �� �h 8�	�h �i � �i ��n ��j  �ޜ� ��� �0 }ܭ� � U�Κ ����  U� 3� ��h`H�Z�r 
����� ��i �� ��y ��z �l ����� ���8�>�� �k �0�,��-~ ���� i�� �� i �� ��y �y �׭t �y ��z �z жz�h`H�Z�� �@�� �� ��� �� ������ ��� � �� ��z�h`H�Z��p �<�q � � �  � �� ���)��&  ����  �  ��� �ύ& ���  w� K� ����s  �ޜs  3ح� ��z�h`H�Z�� �@�� � � �m ��� ��������� ���z�h`H�Z�� ��� �� � ������ ���z�h`�Z�� � �	��������z�`Hڭ  �����h`H�� �  ����� �0�h`H�� �  �	�����	������ �
0�h`Hڪ���




�w ��)w �& �h`H�Z�� H�� H�� H�� H�s �.��%��a��$��d��&
��Z��� �Z�mv �� ��w �q ����� ��� �p ��-~ ��� �� i �� Ȳ�-~ ��� ��w ���p �p h�� h�� h�� h�� z�h`H�Z
��� �� � ���$��a��.��d�8�7�s  p�Ȁ�z�h`� � � �  �� �� � � � � � � � �* �W �` � ���X �d `H�Z� ���%�; � ��4 � �5 �  ��; �; �6 � �� ���%�H � ��A � �B �  z��H �H �C � $� ���X� ���� � �� � � �  K� ����- � ��& � �' �  ��� � � � ;��- �- �( � �� �� w�z�h`� �� ȱ� ȱ� ȱ� ȱ� )
��E� �E� � )0�" ȱ����X �d Ȍ � �  � �L#�!  �� �� � ��! ��Ȍ! � ���1 �2�4 ȱ2�5 ȱ2�6 ȱ2�7 ȱ2�8 )
��E�9 �E�: �8 )0�= ȱ2����X �d Ȍ1 �; �< �6 � �� � � �^ )����� �>  $�`�> �?�A ȱ?�B ȱ?�C ȱ?�D ȱ?�E )
��E�F �E�G �E )0�J ȱ?����X �d Ȍ> �H �I �C � Ш� � � �^ )��@З��� �1  �䀊�# �$�& ȱ$�' ȱ$�( ȱ$�) ȱ$�* )
��E�+ �E�, �* )0�0 ȱ$����X �d Ȍ# �- �. �( � Ч�/  -�� ��$ � ��/ ��Ȍ/ �# ���Z 
���\ ��] �\� ȱ\� `�Z 
��#�\ �#�] �\�$ ȱ\�% `H�Z� )?	@�K � I��-K �K �  ��� )@��J��K �K �" �8��" �� )0�" Ȍ  �����  � �  �K � z�h`H�Z�) )?	@�K �) I��-K �K �. �+��* )@��J��K �K �0 �8��0 ��* )0�0 Ȍ. �+����. �* �. �K � z�h`H�Z�7 )?	@�K �7 I��-K �K �< �9��8 )@��J��K �K �= �8��= ��8 )0�= Ȍ< �9����< �8 �< �K � z�h`H�Z�D )?	@�K �D I��-K �K �I �F��E )@��J��K �K �J �8��J ��E )0�J ȌI �F����I �E �I �K � z�h`� `� `H�Z�X ���%�Y ���X �` �Y )?
��e�b �e�c �a  $�z�h`�` �* �W `�a �b�S ȱb�M ȱb�N ȱb�T )
��E�P �E�Q �T )0�U Ȍa �O �R �S � m�d `�` �* �W `H�Z�` ���L�M �V �S I�V )��V �R �P��T )@��J��V �V �U �8��U ��T )0�U ȌR �P����R �T �R �S )�K �Y )����
�@����K �K �V �( �K �W ��* �W �O �O �N � $�z�h`H�Z�  �  -� �# ��! �/  ;� �� K� �� ���� z�h`H�Z� � �
� � ��_ �^ )?�_ �Q�� �K�_ 
��]�2 �a�? �]�3 �a�@ �1 �> � � � �^ )�����  $�^ ���  �� ��z�h` ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���<������ ��� ���.��.�� ��� ���T����.��T<�� ��� ��� ��� ��� ��� ��� ���     � ��� ��� ��� ��� ��� �<������ ��� ���.��.�� ��� ���T����.��}<��}��}�� ��� �����}��}��}�� ��� ���.<��}��}�� ���     � ��� ���.��T��T�� ��� ��� �<��.�� ��� ��� ��� ��� ���.�� ��� ��� ��� �<��.��.�� ��� ��� ��� ���T��T�� ��� ��� �<�� ��� �� �� ��� �� �� ��� �w�     � �� �� �<�� ��� �� �� ��� �� �� ��� ��� ��� �<��     ���\���<��\������<��\���� �<�������:�����:���<����\�����\���<��     � �� ��� ��� ��� ��� d��     �     � �
�� /d��     � /n��     � �
	�
�
	�
	�
��
�

		�
	�			�
�+�9�=�A�5�;�?�C����S�=�  ��              ]�`��������������9�Q��?�k�~���O   �      O   O   O   O   _   o      �   �      �Z    ����������,�2�PRESSaSTARTaBUTTON$ROUND$CONTINUE$END$SCORE$HIGHaSCORE$aaaPLEASEaSELECTaa$PAUSE$GAMEaOVER$"� �!�|�਍��U����Z�ǰ4����D�TG;GTG;GTG;GTG;GT
G	;GTG;GT         �		p��`����h����ȆΆԆچ�������9��v	�z���:��"�b�����:�z�:�z���⣺���:�"�b����:�z���z�����ȃȃ�H���Ȅ�H���ȅ�H���������ޞ�^���ޟ�^���ޠ�ޡ^����^��������������� �� �0�@�P�`�p����������������� �� �0�@�P�`�p��������������� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �<<<<�    ������    � �� �    ����    ������    �< � �    �0 �<<�    ���� � �     �<�<<�    �8<� �  ��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                          O� �c�