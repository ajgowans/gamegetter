>@BDFHJLNNPRTVXXXZZ Z"Z$Z&X(X*X,V-T.R.P.P.N-L-J,H+H)H'H%H#H!HHHHHFDDDBBBB B"B$B&B'@(>(>(>'<&<$<#<"<!< :888 6!6#6%6'6)6+6+6,4-2-0-.-.,,,*+(*()&)$("'"'"& & $ $ "    "$$(*,.02468:<>�>@BDFHJLNNPRTVXXXZZ Z"Z$Z&X(X*X,V-T.R.P.P.N-L,J+J*H)H(F'F%F$D#B"@!> < :!:"8"8#6$6%4'4(4*2+0+0,.-,-*,(,(+&*&)$("("'"' ' & % % # !  "$$(*,.02468:<>�>@BDFHJLNPRTTVVVVTTRPNLJHHFFFFFFDB@><<:866!6#6%6'6(6)8*:,<->-@-B-D-F-F-H-H-H,H,H+H+J+J+L+N+P+P*R*R*R)R'R&R%P$N$L$J$H$F$D$B$@$>$<$:$8$6$4$4%2%0&0'.(.*.+.,,,,-,-*-(-&-&,$,"+"* ) ( & % # " !    " """"""""$&(*,,.02468:<>�>@BDFHJLLNPRTVVVV V"V$T&T'R(R)P+N+N,L-J-H-F-D-B-@->-<,:+8+8*6(6&6$6"6 66688:<>@BDFHHHJJJ!J#H#H$F$D$B$@$>$<$:$8$6$4$2$0$0$0%0&0'0'.','*'('&'&'&&$&$%$#$!$&&&(**,.02468:<=>�>@BDFHJLNNPRRTVVVVVT R!P"P#N$L%J&J'H'F'D'D'B'B'B(B(B)B)@)>)<):)8)6(4'2&2%0$.",",!* * ( & & &$$$$&&(*,.02468::<<<<<<>@BDFHHJJLLLL J J!H!F!D!B!B!@!@!@ @ @@><:8642220000000022468:<>�>@BDDDFFFFFFHHHJLNPPRRRRRTTTVVV T!T#R%P&N&L%J$J"H HHHHFFFDB@><<< <"<$<&:':)8*6+4+2*0).(,',&,$,".!0 2246888::::8886420.,***** ( (!&!$!$!$ " """""""$$$$$$$$$$&&&(*,.022468:<>�>@BDFHHJLNNPRTTTVVVV V"T#R$P%N&L&J&H&F&D&D&D%B%B$B"B BBDDFHHHJJJ!J#J%J'J)H*F+D,B-@->->,<,<+<)<'<&<%<%<%>%>%>%>$>#>!>>><<::8664444 4!4"2"2#0#.#,#*#(#&#&#&$$$$%$&$'$($)&)&*&*(***,*,*,).).(.&.$.". ,,*(&$$$""""$$&(*,.02222468:<>�>@BDFHHHJJJJHHFDB@><:88866666688:<>@BDDFFFFFFHHJLNPP R!T"T#T%R'R)P)N*L+J+H+F+F+D+D+D*D*D)D)B)@)>)<):)8)6)6)6(4(4'4%4#4!4 6 68:<>@BBB D D!D#D$B$B%@%>%<%:%8%6%4%2%0%.%,$*#("(!& &&&(((*,.02468:<>�UUUUUUUUUUUUUUU TUUUUUUUUUUUUUUUUUUUUUUUUUUUUU TUUUUU @UUUUUUUUUUUUUUUUUUUUUUUUUUUUU@P�WUUUU   VUUUUUUUUUUUUUUUUUUUUUUUUUUU��PUUU  �VUUUUUUUUUUUUUUUUUUUUUUUUUUUP� PUU  �\UUUUUUUUUUUUUUUUUUUUUUUUUUUATvTTU  �^� PUUUUUUUUUU�ZUUUUUUUUUUUD�� �VPU�ξ<��UUUUUUUUU��jUUUUUUUUUUU �@UfjU���/��WUUUUUUU��	�UUUUUUUUUUU E�P������>0 �TTU P�ZVVUUUUUUUUUU ��t����</� <�S@@U   ��PZUUUUUUUUUU@�=��� 
0�0,� ?���
�  ��V�^UUUUUUUUUU��M�� �
 � ����> �/
0��c�T�_UUUUUUUUUP��C�� � 0 	����?�� �\ ��_UUUUUUUU TV7��=�(" �@�?�� ���  � T�_UUUUUUUUdTeUi> �� � ��? �� ���   ���_UUUUUUUUYUVe�? ��   ��� �� �?� � U�_UUUUUUUU &��C��/"(���������� �??0`fUe~UUUUUUUU e�������  ���������<"?��I�|UUUUUUUUY=dՙ� �� ��������(  jT �UUUUUUUU@EU_�ꪀ �� �?���������   XU�uUUUUUUU EYWe������������� ��� 0 �TU�WUUUUUUU@ieW�.�(��
��?��������   �	V�wUUUUUUPUUW�� ��� 0����������� �U�^UUUUUUPU�U/ *��+ 蠀������� � � ЦU�_UUUUUU�Z�Ճ ����*���������   ���E�_UUUUUUPU}� �(�*��#*�*+����? � EjV�_UUUUUU UU]?  �"* #
�������?    E�W�UUUUUU e�? � *�0� ������k�@? 0f�e�UUUUUU ju�� "�� "���
����� �
TyE}^UUUUUU eu�  ( 8��*��i����BP�A�UUUUUUD�U�  (��"����/���Z��
0  PU��UUUUUUDU�7   * �
����늪�fo*����PhU�WUUUUUTV�?  �*  (��(ﯣ������?� �V�AZE�[UUUUde�  ���?��������fj��� Ze�V�oUUUUe־ � ( ��>������گ�����j��U���_UUUE��^��     �?��������������jZ@�i���WUU                                                                                               ?                                       <                                                               �3                                    ���            ?                        �           3                       ��           <                        ��                                  �           3                       ��           ?                       �           3                       ��   �
      <           �           �   �!      ?           �6           ��  ���      ?           �           �  ���<     <           ��          ��  ���     ?           |#          �  ���   ��           �#
          ��  ��+   ��           o+          �  ���   ��           ��          ��  ��+   �<          �<
          � T���   �     �   ���          �� T��+   �� �   `  ���2          �� U���   �� �   `  ����         ��WP��+   �� ��*�j  �?��        ��������  �  �
�i 3?��?        ��ÿ����+� <   ?��e?�3/�0        ������������� ȫ��e��?��?        ������+����� ��(�U����;?�0�?      ����� ����� ?�3 ��OV2�������?��      �������+����� ������??���<�<��     ����?��:���3��� ���������#?��3�,/   ���0��ÿ�+?���<0��꿊�0��#?���ﳺ�  ���0�������<���
�������2?�����#�
 ����������������������������������������          �                                       �                                       0                                      0      
                               �                                     �?      
                               �                                     �     �*                              ���     ��                               �0     ��                              �<    � <                             ���   0���                             ���    ���?                             �<    ��0�                             �<    ��0�                             ���   ���0                             ���    ����                             ���    ����                          ���   ������        ?                  ���   � ���        ���                ���   �����      ��3�                ���   ����2      �����0              ���   ������     �������              ���   �
   �
     �������              ��   (����(     ����*��            �� ��< ��������   �?��  �0            ����< ��﫢�� � ��������0        �
�����>  �ﻢ?  �  猪����?        ���  
��>  ����  � �*���*�
        ��*�
��:�  �﫢  � �*���*�
       ��(�����
� ��������  ���������
       �( ����� �?�?       ������������       ��
�� ?3< ��������� ���
       �     ����*0���<� �?       ����?��������    ������������������������������;���  ����������������������������������������                                                                                                                                                                                                                       �                                   �                                      �	                                      �%                                      ��                                    W  �	                         �0     |	  `	                          �      ��  X                             �     W �                                  |	�%                        ��         ��c	                                   �k                                    l�      �       <                       =      ` �    :                     ���      �	 �    /                �     �on      & &    /                �    �_q	      ��	    /               �3     ��%      `o    �                    ����     ��    ��               �    p��\	     �9    ��               ��   \��p%     p�   �              ���  �����     ��   ï              0? �%�� �     �o ��̎              ���< `	�� �    ���	�����              �?��� `¯� � �  `��&��:�  ��       ����������� �� �𪚰�:� ��
*       ����   ���
 ��? ����/����(     �k���< ��¯������� ��
�Ͽ�����   �������<��ʿ��*�������������������
   ���0��������ꯪ����������������" � ����������������������������������������                                                                                               ?                                      ��                                    � �                                  � 3 �                                �  3 �                              �������?��                             ��30     �?                            ����?����?��                      �    ������������                      �   ������������                      �   ��� ��  ��                       0   �������<�=�                       0   �����������                       0   �����?�����2                       <   ���2�<(��;�2                       ,   �����<(��/�2                       ,   �����,��/�3                       ,   ���2��,��/�2                       ,   �����/��/�3                       ,   �����/��/�2                       �   �����/��/�2    �                 l� ����2��.��/�2    �                ,� �������/��/�2    �?    �           l� ������/��,�2    ��    ?0           � ������/��/�2   ��������          Ã ������/��/�2   ��    ��          ,ó �����,��#�2   �?������           ,������Ϗ�����>   ��33�3�          ,ó<��         �� �303333�           ���?�?������������� �?03333�        ������� � 0    ��0?03333��      �������?��?��3����?�����?��33���      ����������    �0   ���?0� ����*  ����������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�W��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU����WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���?�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU=0 ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU   �WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�     �UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU    ���UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�      ��WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU=   �  ��UUUUUUUUUUUUUUUUUUUUUUUUUUUUU�� � ���UUUUUUUUUUUUUUUUUUUUUUUUUUUUU= �  � �o�WUUUUUUUUUUUUUUUUUUUUUUUUUUU��� �3 �UUUUUUUUUUUUUUUUUUUUUUUUUUU= ? � ���WUUUUUUUUUUUUUUUUUUUUUUUUU������; ?���_UUUUUUUUUUUUUUUUUUUUUUUUU= (��?� ̰�~�UUUUUUUUUUUUUUUUUUUUUUUU�� ����
 <�Sz�_UUUUUUUUUUUUUUUUUUUUUU� �
>���0�0����UUUUUUUUUUUUUUUUUUUUUU=  ����̀2�< ����_UUUUUUUUUUUUUUUUUUUU� ������3�� �T���UUUUUUUUUUUUUUUUUUUU? �����������? ��?�_UUUUUUUUUUUUUUUUUU� ��/���������������UUUUUUUUUUUUUUUUU� �������������������_UUUUUUUUUUUUUUU� ���������� ���(P�P��_UUUUUUUUUUUUU� ����??  ��3  �?  �W����WUUUUUUUUUU������ ��  0�      ��U�T��_UUUUUUU��� ���?3?  �           ? 0��_���UUUUU�������?                  �  � 0��UUU�������������������������������������������������������������*���������������������������������������Z���������������������������������������Z���������������������������������������V���������������������������������������U��������������������������������������jU�������������������������������������jU�������������������������������������ZY�������������������������������������Za�������������������������������������V������������������������������������U�����������������������������������jU �jU��������������������������������jU PVU������������������������������ZU @UEA �����������������������������UU @T@@���������������������������XUU @ P A�������������������������U`UUUU@  U ���Z��������������������jUUUUUU   TD���V��������������������jUUUUUU   P��VU��������������������ZUUUUUU  @UAAUUU��������������������ZUUUUUU PP  TQUUU�����������j�������VUUUUUU  @ PUUUU�����������j�������UUUUUUUU     UUUUUU ����������V������jUUUUUUUU     PUUUUU����������U������ZUUUUUUUU     @UUUUU���������ZUU@�����VUUUUUUUU      UUUUU���������ZUUP��ZjUUUUUUUUU      TUUUU���������UUUU�VUUUUUUUUUUU      PUUUU  �������jUUUUTUUUUUUUUUUUUU     @UUUU  �������VUUUUUUUUUUUUUUUUUUU      UUU   �����jUUUUUUUUUUUUUUUUUUUU      TUU   �����UUUUUUUUUUUUUUUUUUUUUU       TU   ����ZUUUUUUUUUUUUUUUUUUUUUU       UU    ��jUUUUUUUUUUUUUUUUUUUUUUU        @   ��ZUUUUUUUUUUUUUUUUUUUUUUUU         P   �                                                                                                                  �                                       �                                       �                      ����            �                      (�
�*            �                     �
�
��           �                     �*�
��
          �                    ��
��*          h
                    ��
j�*          �
                 ���*��
Z�*          �                 �
�������          �                 ��
�����*
          �                  �*��*����*                         ��* *�������   TU                   ��� *��*
b���   @     �
            ����((�
b*�
   DD  @ �(            (���*�(�(b���   DDT�
  ��            (�����*�b�*�  DD �"@ ��         P  ���������b���   DDT��  ��         @ 
"�"���*b��
 TDD ��@ ��         P     *����b��  DDT��  �*        �PP �"����� b�"@UDD �*@T�
        �@  "
���� b�"@  DDT�
@E         �@  "
*��� b�"T PDD �@@!        ��*J  "
(��� b�" DDT� %XU      ����
  "
*��� b�"TUPUD �%HP        ��"
(����b�"  TDT� � !H      �������"
*����b�" DTD � �  HP        ���"
(����b�bEDDTD��  �*       �������"
*����
b�"  DT�(� ��"  �        ���
"
(����
b�"EDDT��� � *((     ������"
*����b�"  DT����  �**�"        ��� "
(����
b�"EDT�*���"�����      �����   "
*����b�"  ���*����*��
  ��������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ���           ��0�          �� �      ���������?       �<�          �3<�          ���                                                                                                                                                   �         ����������   �     �    �                           0 �            � �        �    0           0       �    0       �    0       �    0       �    0       �    �     � �    �     �    �    � �    �    � �    �    � �    �    � �    �    � �    �0    � �    ��   � 00    0 �   � �    0    �       0    �         �  �    0      ? 0    �     ��     � �             �?     ��<�<?        �<<���        �<<���     ��?�?<<����     �<<<��        �<<<��        ��<�<��                                                                                                                                                  �         ����������   �     �    �                           0 �            � �             0             0             0             0             0             0             �             �             �      �     �      �     �     �      �       0    �       �    �    �       �0    �       0�   0       0 <   0       0 �       0           �     < �         �<      � �    �       �?    �?����     � �<?�0      � �<?�     �����<�� ��?    � ��?��       � ��<��0      � �<��                                                                                                                                                �            ��������     �  �     0             �    �         �    0         �  ��         �             0 �        ���� �        �     �      ���     �     �       �     <        �                 �             �             �             �             �������     ��      0     <�      �     �      �    �       �    �       �  0  �       0  � �     ��   < 0  0        ��  ����                     ����< ?<�    ��<�<����3    ��<�<�����   ���<�<������  ��<�<��<��    ��<�<��<�3    ��������<�                                                                                                                                                �          ��������          �                �     �             �             0         �    0                       0             �  �           �  �    ����  �  0       0  �  0   �    �  �     �    �  �     �    �  �     �    �  �     �    0  �    ������  0    �       0  0  �         ����             �                   �             0        �                 �          ����                     ���?���     �0� �0      � � �     ���<���� ���   �0�� �       �0�� �0      ��?���                                                                                                                                                �           ��������       0  �    ?             �                          0  ������     �  0         �      ����  �           �           �           �    0       �  0  ����   0  ��                ��� �    �        <                         �       �      <            �        0  ��?         �  �            ���                                                                                     ����       ��<��<?       ��<��<?     ����<��<���     ��?�?�       ��<�<�       <�<�<                                                          �             <    ��     � �   0 �     �           �  0     0    �  �     �  � 0  �      ����  �        �    �             �             �     ��           0         �  �  �    �   � �   0 �    �    0 � �   ��    � � �   00    � � �  �    � � � �      �  0     0  0  ��     0  0    0     �           �                       �           �?     0  �           �  �             0            �              �                                                        �00����0      30��0      00�0�3   ���03��0��?��    �33�0�<      �33��0      ������0                                                                                                                                                 �           �����?         �  � �     ����     <             �    �             �             �          �       �?        �  0�    �   <        0   �  0 �  �      � 0  �    0  �� �  �    �  �� �  �    �  �� �  �    �  �� �  0  ����  �� �    0 �   �� � �   �   � � <    �    ���    �     �      �     �     0 0     0     ��                 �           0 <            ��                      <��?���     <�����<      ������<   ��?<������<��   �������<      <������<      <?0���<                                                                     ����             0         �    �         �    �         �    �         � �  0       �������      �  � �         0  �             �             �                                    �    �         �     ?        �     ���      �       �      �       ��?    �   ����  �   �   0     <           �               �                       ������                                    0      �       ����  <            �           ��?                                                                   ��                              � <                              �  �                            �?  �                            �?  �                            ?�   ?                            �?  �                            ��� �       <                  � �� �     ��                  �� � �     ��                 ��� � �     ��                 ����� �    <<�                 ? � �  �   �?�                � �? �  �   �3<                �  �? �  �   << <               �� �? � �   ? <               ��  ? � �  ?��<               ��  ? ���  �? �?<               ��   ��  �< ��?              ���   �� �  �?             �����  ��?  �  ��             �� ??  ��  �?  ��           ��� ��  ��   ��?  ���           ���  �  <��  � �  ���          ���  � 0��  �� �  ���         �� �  � 0�  �� � ���        �� � � �?  �� � � �?        �� � � �  � � � � �        �� �? �?     � � � �       � ���  ?    � � �? �         �? �� � �    � � �? �        ��� �� � �    � �  � ��       �� �3 �? �   �? ?   � ��       �? � �3  � �   ??�   ��?       � < �?  �<  �?����?  ��        �  <  ?  �   �� � �� ��        ��     �?  ��� ����        ���    �  �  � �?��?       �����    �  �  <� ����      �������      �  <�  ���       ���? � ?     �  ��?  �?       ����? �? �    �  � ?  ��       �� � �� �    �?  � �  �       < �  �  ��     ?� � �            <  � ��     ��� �            � �?�      ��? �          ��� ��      ��� �          0 �� ��      ���  �          ?� ��? �?       ��?  �?          ?0���?         �?    ?          ?  �? �          �/              �  �? �           ?               �   � �          �               �  � �          �               �  �?           �              �  �?           �              �?  �?            �              �? ��            ��              �� ��            �/              ����?             �               ���             �                ���                               ��                                �                                                     ��                             ��                           ���? �             �    (    �?�? �             �?    *   �?�����            ���   ��   �3�?�� �           ���* @U  ������           ��*�
TUU ��?�? ��
           ��BUiUU% �3����;           �( P�UU
 ����� �0?;           � U�U�
 ���?  0��           �@U�V�*�
��� /��          �@U��*�*��������          �PU�*���*����?��          �k�����������<��          ���� ������ ?<          ����  ?�����3?�<          �S	���* �<����?*��<��          �C	������<����/(�����          �O	�*U������ �?���         �O%�ZUQ����������?�        @N%�@U�ʣ���������        TN�l@UE��
��?�:������       @U�JAUU������*����?       TUU. XAh�����
��
����?       UU� XAU
��
�
���*����?      PUU� ZAU���� �*���������      UU��Z���
��*���������     PUU� �Z����
��*���������    TUU
 ��Z��������*��������    HUU�  ��Z�����������������    jUU* ���VA���*������> �����    jU� ���VA��*���*��� �����    �U*  ���V������«�� �����?    ��  Ȫ�V�����*���
 �����    �*   (��V�*���¯��  �����     �
   ���� �
������* �����     �
   ������(��"��� �j���      �*� �����������* ��V��       ** �����* ����
 �ZU��        � ���*T*���*��  �U�         �0���� �
"��
 �eY**        �򠪪�*���  ��� �Z��*         �򠪪����� j� �����
        ����P��* ��( ��*�
�        ��ʃ��*P����  �" �����
       ���
��
����� (������*        ���*��@���ʯ�  ��ꫪ�        ��<�.<�*@��*�[� �����
        ��?��<�
T��
���*����*         ?��������*�k����ꫂ        �?�����D)� ��j
 ���*(         ����������𫪪�����
        ������   ���* �����        � ��?���  ����� ���*          ����00* �����* ��ꪨ          ���� �
������
 ����
          ?��?�?3󫪪���  ��* (         ���<�<������� ����*�         ��? ��������� ����
"          ��<0�������* �����(          ?�� �������
 ���* �           ?�?�������  �ꣀ            >�? ��3���
 �տ�
            �� <��?��� Z���"             ����0�ü�* �����             ���<���� h���"              ������ �V�**               ��� ����
 `����               (?�?0��3? Z�*�
               ��?����������                �������h���
               ��� �?���V���                �?�?������*�                 ��?�������*�
                 �
?� �����*�                  
��?�������*                  ���?�������                   ���� ������                    ����������
                    �������?                     �������                     ��?����?                      �������                       �������                        ���?��?                        ���?��                        �����                         �����                         �����                           ��                           �                                            �                       �> �?           *       �� ?�          ��  �  ������         ��  T �;��?�         ��� U����0�<         � ^�WU� ,2�� ��?         ��U_�* ���?�??�         �� T_9���������         ��P���
�����        ����� �2�*�����        ���� �2�����?��        ����  ¨*��?�        ����� �
����
3��?        �U�ZU������>,���?        �W�TU������/*���?       @��nPU�������*����       T�+`PU)����� ����      @U�TPU
���� ������      PU�VP�*����������      U���VP������������     PU�������
��*�� ���     TU
��V��*������
 ���    @U� ��VP�����������?   @UU* ��V�*������* ���   XU� 
�������诪����    hU�  ����(����* ���    ��
  ��������������     ��   ��*������� �      �*� ����  ���
 ��*      ��(��*��  ��� ���
       �ȫ�*��
 ��* ���       �򨪪���� �� ����        ����*���� �* ��*
        �����
���
�� ��
         ���� ����  ��*        ��
�����
������        ���*�
�����*���"        ��*������*��+�        �?������
�
 ��
        ����*  𯪪 ���         ��� �
 ����* ���       ��� � ���� ��         ����� ����* �+�        ?3? �3�����
 ���         ��<������ �+�         ����3����
 ���          ���;������  �**          ����Ϡ��* �/�           � �?���� ��           ?���* ���           ������ �            ������: ���             ���?� ��"             ��?0�����*             <�?�����
             ������?���              ���?�����
              ��������              ���������*               �������                �??����+                 ??<����                 �?<����                 �������                  ������                  �����                  ����?                    ���                    �?�?                     ��                         �?                 ��     �          0�    ?<          0 ?@ ����        0�T ?3�?        0(�V)����<        0T�
���?0�        0U+*0�� �        0H�*��� ��       0�����?���       p�����?��?       u)n)*�*? ��?      @��R��������?      T��QU����(���     @UͨQ����
 ���     T��jQ��
������    @U5�j���������   TU�jP���������  �U� �j����*�.���   V 
Z���������   �  ���

�� ��   ( �����(
��
 �?    � ��*�"
��� ��    � ��
*"���* ��     �����*������     ��*�� �� �i      ��
��
 �
��     �
������� �*     ��
���
���8     �����*��* ��     ��?�  �� �"     ��� ���� �     �0�������* ��      �0�����
      ������� �
      � �󨪪
��*       �� ����*       ?� ��*���        ��0����**        ������* ��        ��� ���*         �������         ������ë�          �����*
          �??����            �� ���            ��0���            ��<�?             ����             �����              ��?�?               ���               � �                         �       �    ��           ?<         � ���?      �
�0<�      Je����03      ��
����      R������<�      �� ������    `������?�    eW����#��   P�HU������   U/`T��*(���  �� @����**��?  � h�j
��*��?  ��Z���*����?  �
�Z��������?   ��j��*��*��   ���*����
��    ���*(��� �   �
�

���
�   �����*��� �
   ?��*����*�*   �ÿ����*��    <��� ����   ��<������    �� ����*�+
    �? Ϫ���     ?����� /*     �<���
�     �?�ϯ� /"      �<�3�
�      �?�3� <�       ����?��       ��??��        ��3��+        ��3���         ����*          ����          �?��           ���             ?                           @ �     � T- ?�    Sբ��?<    �-���0    �V��? �    ����?��   P�~���?��  UF����0� `�@������ �F����� � �V�2���� �������� ������� �  ʿ*���
��  ������ �?  ?����
�  ��*��� �  ?����* �   ����� �   �����
�    ?���� �
    ����
�     ��?� �
     ??��      ����
      �����       ���
       ���/        �?�        ���         �?             ��    @��  ��?�  �?0�W  ���� P���W? �s���? 0p���? ������? ������?������������>  �����  y��?   W��    ���    ���     ��     ��     ��      <             �      ���� ����  ��� ����<���� ���?  ���  ��?   �*    �*    �        �����               �   �              ���0<�              �������             �������             �   ;�3             �����:�3             �����:�3             �����Ϋ�           ��� 3������       ���� ��Ϊ���?       �� ̬������       ������������       �������������   ��  �_UU������� ��� �_UU����� 0 ��� ������}U����0 �U ����������Z��3 ��U5 �������U9?���0<����: ��������:?�*��?���: ������:?��j ?���: ������������k�����? ���������  � ���> ���������?��������?�����������   o0  ����������������������     ���������������    ����������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �                  �                                   �                            �                              �                           �                               �                                  �
		##
		��������������̂ڃ����� �.�����čf����Ƒh�
������,�:�H�V�d�ދ�����:�:�:�����@��8�F�T�b�p�~�����<�J�X�Ҏt����p�p�J�p�n�|���������Њr��������L��������������Ά܇�����"�0�>�����$�2�Ԓv�3���̈́ۅ�����!�/�=�K�Y�����?�M���J�b���
�"�z�������z���������ʠ�:�
����2�2�j�J�b�
�"�R�R�J�b�:�z�r�j���Ҟʞ ����
�"���ʠB�:��r�*�����ʡ⡒���������:�2�*����
���z�r�J�b�������z������ʤҤ����ҡҡʡ⡺�����:�R�J�B�:�2�����z�J�¢��r�򢪤
��        %%#!		��R�J�
�
�
�*�j�������j�j���ʞʞꞪ�ʠ
�
���z�:�z�Z�Z��
�J�J�J�j�*�J�J�J�����ʞ�������
�ʠʠ*�Z�:�z�:�����ڡʡ���������*�2����"����r���R�Z�����j�r�������ʤ⤚���ڡ�ҡ⡲����2�b�R�B�2�B�����j�z�����z�򢺤
�"� %#"!
	 �J�b�*��:�J���������z��������Ʝ��
�R��"�r�B�j�J�J�
�"�j�R�z���R�Z�b�r���ʞ�� ���"�ʠ�Z�b�2���*�����ʡҡ���������:�B�B����z���j�R�R�¢��j�j���¤�ʤڤ����ҡҡڡ⡪�����B�R�R�:�B�*�������b�����r��¤�� %$"! 
	��Z�J��"��"�r�����r��������Ҡڠ*�:���:�2�z�Z�J��
�Z�b�R�b�2�j�r������Ҟ �� �����*�2���r�:�����ҡʡ���������
�
�
���
�J�J�j�*�J�����j���������ڤڤ����ʡʡʡꡪ�ʣʣʣ*�*�J�
�
�*�j���J�J���ڢ��������              %#"!
	 �J�R����"�j�������������ҠҠB�"���2�B���Z�b�
��R�R�Z�b�*�z�����ҞҞ�� ������*�*�򠂟B�����ʡ⡪�����ʣ��"�2����
�z���j�2�b���Ң�����¤�ڤʤ�����ҡ��
�ңڣ��:�B�J�:�B�*�r���J���ڢ⢲�����
�                      %$"! 
	 �J�b�*��:�Z���������z�r��������Ҡ
�R��"�r�B�j�J�J�
�"�j�R�z���Z�R�b�j�����ʞ��  ��ʠ�Z�b�2���*�����ʡڡ������������"������2�J���Z�J�¢������z�2�r��⤊���ҡ�ڡ򡪣��ң�:�*�:��
�B�������r�¢Ң:�r�2�"�"�      %%"" 	�R�J�2��B�R�����������j�����Ʝ��
�R��"�r�B�j�J�J�
�"�j�R�z���R�Z�b�r���ʞ�� ���"�ʠ�Z�b�2���*�����ʡ��������:�B�*�:����b�J�r�:�B�������B��b��Ҥ������"�2�������B�*�2�"�
�2�z���J�J�*�*��2�"�"�� $#!!  �J�R���B�*�r�������R�Z�J�������b�z�������������Z�J�
��R�Z���j�2�Z�b�J�������z�b�R�����r�j��"� �B�����ʡҡ���������:�B�B����z���j�R�R�������R�2�z�ڤʤ����ҡҡڡ⡪�����B�R�R�:�B�*�����j�R�*�*��r�:��
�              %$"! 	 �ʡ⡪�����ڣ��"�*����
�j�����2�R���Ң�����¤�ʤڤ�����ҡ���ڣң��:�2�J�*�B�B�r���J���ڢ⢲����
��J�Z��"��2�j�z�����z�j�z���ʞ�ڠʠB�2��������b�R�
��R�b�Z�r�*�:�R�b�������r��� �
���B�R���򟲡����           � �%%"" 	 �ҡʡ����£ң�"�
�:��������j�2�b���Ң�����¤�ʤʤ�����ҡ��
�ңڣ��:�B�J�:�B�*�r���J���ڢ⢲����
�
�J�z�*�2�b�r���������j�r��ʞ򞺠 
�
�j�j�r��b�R�
�:�j�r�����z���j�z��������������ʠʠ��������������                � � �$#!!  �ʡҡ����£����"�
�ңڣʣ:�"�����2�*�"�b���*��ڤʤ����ҡڡ�ꡲ�ڣ�ʣ��
����ң"�:���b���B�j�¤�
�J�R����"�j�������������ҠҠ*��j�j�ҟ���J�J�
��R�R�Z�b�*�z�����ҞҞ�� �����Ҡ������򟪡����     � �%$"! 	 �J�Z����"�z��������������ʠҠ:����:�B�r�Z�Z�
��R�R�Z�b�:�j�r���ʞʞ������
����Ҡ*�*�����2�����ʡڡ������£����ڣ��:�:�j�b�Z�2�:���B��:�ʤҤ����ʡڡʡ���£��£�*�2�����*�z�z����B�*��*���
��  %%#" 	 ���ꡪ�ңңң��
�"�ڣ���J�Z�B�:��*�B����*��z�ʤʤ��������ңңʣ��:�*�
���z�B���:�B��2�:�
�
�   %%"" 	
	 ���ڣ���Z�Z���j�*�R�Z���¢¢��Z�2�*���2���:�ڤڤ�����"�*�2���B�*�j�����b�����¢����B�2��:���ڤڤ  %%"!	 �ʡʡ��������ҡڡڡڡ��������*�"��j�����*��z�ʤʤ����ҡҡҡҡ��������ڡ����ڣң�b�R�*�R�2�B��2�:�
�
��       %%$" 
	ʡڡ����������*�2�B��
�
�r�j�r�J�R�����j�j���¤�ڤڤ����ҡҡڡ⡺����B�J�J�2�*�2�����z�R�����z������J�Z�
��
�B�r���r���Z�j�r�������ڠ������j�j���J�R�
��J�Z�J���2�B�2�B�������z�z�������r�z�������z�����         �  �� � ���%%#" 	 ��j�j�*�R�R�R���������Z�z�j�ʞڞ��������r�z���r���J�J�*�*�j�������R�R�J�b���������������r�r�����j���������         �    � �����������%%"" 
		 �j�r�Z�b�j�r�ڞڞ�Ɦ�Ҡڠ"�B�B��ڠ������r���z���Z�Z�*�2������������� ��������B��r�j���r���z�Z�Z�                  � �����%%"!	 �J�J�����R�Z�Z�Z��:�:�������������r�����r���J�J�
�
�R�R�R�R�����Z�z�z�Z�R�j��Ҟ��Ҡ��j���������%%#! 	 �     � ����z�
�R����*�l����������h�0 � �� 0 0 � � 0  ��?�  �00� ? ? ? ���   PPP      �����?<    << �? <��?��?�� �:��� �:����:����:�����?< �? <<    <�����?         ��? 0<0��:��:<0 0��?     �?00�?  �����   �   �0  �<  ��� ��������?����������<���0 ��  ��  ��   �����������   �   �  �  <� ����������������������<��� ��?  �  �   �����������   �0  �<  �������?���������������<���0 ��  ��  ��  ��   �����������   �  �  <������������������������<��� ���  ���  ���  �   ���������������������������*                     ���������������������""                    ""                    ""                    ""                    ""                 0  ""                 0  "" ��<<?���        03""����<0��       ��""���< ��       033""����<��       00"" ���<���       0 "" ��<<��       0� ""��� < ��        � ""��� <0��        0"" �� <?���         ""                  ""                  3""                   3""                   3""�3?               ""�0<               ""�0�              ""�0               ""�0              ""�                  ""�   ?               ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    ""                    "" ��<���           ""  ����           ""  ���0           ""  ��?�           ""  ��<�           ""  ������<           ""  ������0           ""  � ����           "" �� ����           ""                    ""                    ""                    "���������������������"                     ���������������������*      �  �?�����
  �  �*�
�* �� �����������?�����������/�
���?  ��      �  �?�����  �  �*�
�*�*���*������������ ����������*�
���*  ���* �������   <    ���* ��
����<������������ ������?�����?�����?�? ���* �������   <    ���* ��
����<������뫾��������� <�����?�����?�? ����
 �� ����*   <  �
��* �*��� ��+<�?������> ��>��������������������� ����
 �� ����*   <  �
��* �*��� ��+<�?������������< ����������������� ������������ <�< �����*0�? �?�����:�����?�����������?����?  ������ (  �*��.��(�*�������3������� ��� ���� < �(?�<�����<�� ��03��<��    �    � �  ? �  Ͽ�  ���  ���?���>??������?��������?  �    ��    ��  � �  �� �  ���  ����?��������?�������?������  ���� ��* ������ ������ ��:���
��: �� ��� ��: ������  ������� �� ��: �� ��� ��:  ����� �� ��  �� �� ��: ��  �� ��: ��  �:  �� ��  �� ��  �: �� �:  �  ��  �:  �� ��   � �� �  �  �:  �  ��  �:   � ��  �  �   �  �  �:  �   �  �:  �   ;   �  �   �  �   ;  �  >      �   >   �  �   �  �                :       �       �   �  �  �  �  �:  �:   �  ;   �   �   �  �  �  �   ;     <   <   �   �   �  �      �  0 :   � �  :  � 0�   0   : �  0 �  : � � �      : 0   � � : 0 � � �   �  :    � 0 :  �� � 0 �  0  :  �  �  :  �0 �  0    :�  0  �  :�  � �      :0    ��  :0  � ��    �   :    �0  :  ��  �0  �   3   :  �   �  :  �3  �  >      �   >   �  �   �  �                    :       �   �       :  :  �0  �0  ��  3   �   �   :  :  �  �  �3  /   <   >   �   �   �  �  �   ��: ������ ��:��������� ��� ��: ��� �� ��:��� ����� ��� ��: ��� �� ��: �� �����  �� ��:  �� �� ��: �� �� ��  ��  �:  �� ��  �: �� �� ��  ��  �:  ��  �  �: ��  � ��  ��  �:  ��  �  �:  �  � ��   �  �:   �  �  �:  �  �  �   �   ;   �  �   ;  �  �  �   �   <   �      <  �     �   �   �       �       �       �       �  �:  �:  �  �  �  �  �    �   ;   ;  �  �  �  �  �    �   <   <        �  �  �   �  ��  �  �0  ��  � ��0  �  � 0 �  �  ��  �  �0 ���  � 0 � � � 0 � � �  �  �� ��  � � �  � 0 � � �  � 0 � ��  �  �  � � �  � 0 � � � �� 0 �  �  0�  �  � � �  � 0�� � �  0�  ��  �  0�  �  � ���  �  ��   �  0�  ��  �  0�  ê  �   �   �  ��   �  0�  ��  ̪  0�   �   �   �   �  �W   _  �  ��       �       �       �       �   �  ��  ��  0�  0�  �  �  ê   �   �   �  ��  ��  0�  0�  ̪   �   <   �   �   _  �W  �W  �V�0<<<<<<<<<<<<<<<<<<<<<<0�����������������<< < < < <��< < < < < <0�?�<< < < < < �  < < < <<<� ���<<<�?      �?< < < < < � < < < < < <<<��80<0< < < < �<<<<<<<<<<<<�� < < < < < < < < < < < < < �<<<<<<<<<<<<�<<<<<<<<<<<<��<<<<<<<<<<<<�? < < < <<�  �///////////�/  �������/  �/// /�// //�/  �/// /�/ ///�/  ������/�  �// / �/ ///�/  �//// �/////�/  �/// /����  �/////�/////�/  �/////�/ ///�/��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?                    �    �              ��  �00��00���33030�3�����������������      �      ��?���<��<��<��<��<��<��<�����<��<���?<���      �      �      ��������?��� ����������������� ������� ���������<����� ������� �<�?�<�<�<�<��� � ������������?       �       �       ���?������0�� ��0��� ������������<��� ��0��       �       �       ���������?H�Z��� � ������ ��������  s���r� �������������� � ��� s������� ���� s���D� ��L�� �� �������� � � ���i��  s��� �� ���8���  s���� ��L�����  ���d� � ��z�h`�
����� 车��  ��`H� � s����h`H�� � ��h`���� ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                                     0    �   � � �<� � 03 0 ���  �                        �  �              0  �  0�� ��"      �       ( �( 0     � 000 �  �          �( ( �  ��  ��  �0  �� �  0  3�  ��  � �0 �� �� � 3 � � 0< �< <0 ?0                     �                        � �     �� ?    \����   ��:���  ���:��  �����  �����?  ������?  �� ����?  �? �?��    �:��     ���?     ��      [00      [��0      ���0      l��0      ���      ���      ���?      ��:�      ��:�     ���     ��0     ��0     ��0     ��:0     ��:0     ��:0     ���0     ���0     ��:3     ��:�     ��:     ��:3     ��:3     ��:3     ��03     ��0     ��0     ��0     �0     ��     ��?<3    ����?                                                        �     � �     �  � �  �  ���  �  ���?  � ��? �: � ? |�� �<? ��� �?���>� �����;�������������  ����?�:  �Z�0 �   [��0      �z�0      l��0      ���      ���      ���?      ��:�      ��:�     ���     ��0     ��0     ��0     ��:0     ��:0     ��:0     ���0     ���0     ��:3     ��:�     ��:     ��:3     ��:3     ��:3     ��03     ��0     ��0     ��0     �0     ��     ��?<3    ����? ���� 0 ��  0�  0�  ��? ��  0� 0� ?0��30<�0��8���������:2���:���>��>���>���>���>���>���:���:�������� �� �� �� ��: ��: ��: ��: ��: ��: ��: ��: ��: ��: ��: ��: ��: ��: ��? ��� ��   0�   0�   ��?��� <0�� 0� � 0� � 0<�� 0�� �8�#�믫����������:���������>���������� ��� ��  ��  ��  ��  ��  ��  ��  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��:  ��?  ���   ��  �� 0� �0��0 3 ���? <�? �?�� ?�� �<� ��������<��� ��� ��� ��� ��� 0�� 0?� � � � 3 � 3    ��     ��    0�    �0    �0    0     0�?��  ��? �  �? 0< � ? ���� �  ?� �  � ���  �����    ���    ���    ���    ���    ���    0��    0?�    �    �    �    3    � 3  �       �   �   ?      ��<��     �         � P  <  �  �        ?�� ��  ���: ���: ���: ���: ���: ���� �� p��� p��� �� 0��� ?����3����0����0����0��:�?��:  ��:  ��:  ��:  ��>  ��  ��  ��  �  �  �� ����  �   ��  �<  �   ��  ���  �<� � �  ��: �� ���������������:�V���Vz���z� �^z9   �   ��  ��?  ���  �3� � � � �: � �: �?; �
�:����:����:�����Z���Z�������n��   �    �?   �0   �3<   �3<   �0   ��3   �   ���  �?� ��< � � ����  ����  ��3 ���3 ���3 ���� 0�� 03�  03?  �  �  �  0  0�     �    �?   �0   �3<   �3<   �0   ��3   �   ��   �? � �� � � � � ��� 3 ���� ������ ���30 ���� 0�� 03�  03?  �  �  �  0  0�     �   0   0   ��   0  ��? ��
< ���3 ���� ����𪪪:����� ���� ��[� ��[� ��[� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ���� ��� �� �� �� �� �� �� �:� �:� �:� �:�  �:�  �:�  ��  ��  �� ��   �    0    0    ��    0   �?<  ��0< �������>������ ����� �����  ����  ��[�  ��[�  ��[�  ����  ����  ����  ����  ����  ����  ����  ����  ����  ����  ���  ��  ��  ��  ��  ��  ��  ��  �:�  �:�  �:�  �:�   �:�   �:�   ��   ��   ��  �� ��  �� 0� �0 �0 0  0�? ��?  �? � ? � ��� �0�������������0������� ��� <�� 0?� � � � 3 � 3   �   �?  �0  �3<  �3<  �0  ��3  �  ��  �?  ��  � �  ��� ���� ���� 0��� ��� ���� 3����0��00?�� �� �  �  3  � 3 ��� �? � ���?   ���? � ����?  ����� �: ����   ���� �: �����𪪪�� �� ����  ����ê� �:��������>����ê��� �����ê��:��j�:��j�ꬩ������� �����ê��9k�V�:��V�ꬩg���eU�  ��eU����g9[�UYꫥ��֬�g�s�e�?  p�e�?��e�e5[f]Y֫UUU�lY�UUs�U   p�U �eUUe5WVsU�WUUU�\UUUUsUU�  pUU��UUUU5WU�U�WUUU�\UUUUsUUU  pUUU�UUUU5WU�U�\UUU5\UUUUsUUU  pUUU�UUUU5WU�U��_U�\UUUUsUUU  pUUU�UUUU5WU�U� pU5 \UUUUsUU�  pUU��UUUU5WU}U� pU5 \U�UUsUU   pUU �U�UU5\UUU� \U5 \UWUsUU�?  pUU�?�U5WU5\UUU5 \U5 \UWUsUUU� pUUU��U5WU5\UUU pU5 \UWU�UUUU �UUUU�U5\U5\UU� pU5 \U\U�UUUU �UUUU�UpU5\UU5  �W pUp� _UUU  _UUUW�U\U�   � ���? ����  �����  ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ���ة��  ��� � �� � �	� �ύ& d� t ���d���� � �������� �XL �H�Z�����+���ə�i������Y���i��d����i��d�d�إ� ���� ��� �
� ��
��	�����������������������Ƒ(z�h@H�Z�' )������ �� ���# �$ �% (z�hX@                                                                                                                                                                                                                                                                             ��n�� �#  o���� q��� � � � 0� �©�� � ��  ��� I� /� � d�  l� � �� c� ʭH����`�D�� �#��i 9� ��� �<��
��"ȍ �"�i@� ���-� �� ��ȍ �  ��� ���`� ���
��IÍ �I�i@� �YÍ�`Í�gÍ �nÍ ��� ��� I�� �ʀ�����<� � �����  l�����  uÜ� � ��D�
�O����� � 9�O`�]�h�o�sv�w8xU\G5* 
	"&-/�
� ����@��"� �í �& I� ��� � �8����`�
��IÍ �I�i@� ��)� ���  ��`�����1�N��� ������#��H� � � �O�� � ��$� ��
 ��	���A�@�B�C� �$ �. ��	���(� �(� �2� �2� �(� ��  ��! ��" ��# �
�=�>�?�- �7�8�P�Q�R�9�:�;��� �� �� �� �� �� �<�6�� �I��� �w ��	���3�4�5�� �� �� �� �� �E��F��G ��`�
���ɍ ��ɍ � ����� � ��� i�� �� �  .�Ȁܭ� 8��� �� 8��� `ڢ �B���B��C�B�����`������ ��!���"`���;�� �h�� �h�� �� �� ����#�� �<��(��������� j�)����!�� �<��(�������U� j���`�� �.� �F��$��(��� � � ��)� ���  �`H�Z� �8�� �	�	���	�,8� ����� �������� m� � i � �� �� ��������� ����#� i0� � i � ���m	���z�h`�(8�� �.� �F��$��(��� � � ��)� ���  ��`H�Z� �8�� �	��	�����	� �8� �i���� �� ������M-����-����0� m� � i � �8��� �� ��������� ����3� i0� � i � � �������m	�L=�z�h`� ��� ���
��"ȍ �"�i@� ���-� �� ��`�B @�GFE�JuR/M�OZ�� �0� �� � 8�d
�� iȍ � i � �
�����FJJ�
8��+� �8��+���1� ���1����1ȱ�,���)���* '�z`�+� �,��*��)��
���ȍ ��ȍ  5�`j�t�~���ک� �0� �� � 8�d
�� iȍ � i � �
�����IJJ�
8��/� �8��/���2� ���2����2ȱi�0���-���. K��`�?�-�/� �0��-��.��
���ɍ 轔ɍ  5�`���������;��� �;��  �����"� ��:�0� �:��:�
�� �:��? �`�Z�
���ɍ ��ɍ �z�`*� ��J���>�ـ	� �é �� � m� ���)��*��+��, '��-��.��/��0 K� �� �� �� T� Jŭ� � �� �� � &� � �� �� �խ � �ީ� � � � �� �� � 2� �� �� _ɩ
� �  	������� ��� ؜ !� Bԩ�� cӭ� ��� �� ��H���LS˭<ɪ� ~̀g����] u�����Lkʭ� ��� /� {حM��$��U������������ ����<���	 �� 	�LS�LR�` Jũ�� �� �� � c� q�<� ��� �H�� �˩���  ��� ���<� ���� �˩���  ���x� ���� �I`H�I�� � )�Ih`�
���̍ 轻̍ ���� ���`�� �H��	������̍ 轻̍  ��` o�� �� �� ����  ���� � �ܩ�������� �F������ ��̍ 轻̍  ���"���$� �� u������� ��� Bԩ�� `� cӭM��$��$ J���������#г I� � ��`�~���Ʃ�Ⱥ�0����� L:��0���	���N�0������<�	0�����	�*�����

��N�� ȹN�� �7 }z�8�� �
��N�� ȹN�� �7 }z�� �id� ��`H��� �� �� )���"�"��h`�D�� �J�� 9�x� � �� � ��`���  l��=�����/��� �D� 9��/��� �D� 9�x��� �D� 9�<ɪ�� 9�"��  �b� w뭂  �b� w뭁  쩆��� � 9�<ɪ�
�d� w��=�
�� � ��=�� π�� Ѐ�� Rр ,Ҁ
��� |�` �D��O�� � �� 9� I� I�� �4�� 9� I� I�� �H�� 9�S��� � 9� �O�� �n��!����
��̍ 轻̍  ��  ����L©F�����  �� }ϩ
� ��  bϭ  ��0� � }�� }ϩ
� � �� bϭ�����ȩ���`�C��� �
��2�� ��`������/0���F���� � ��`�����Z�� ��ύ ���i@� � �� �� ��`�x
���ҍ ��ҍ  ��`�� �]������  ��` �ϩ��� �� ѩ� �x� �  ��L�Э � �Э������� �Щ� ���$� �� ѩ� ѩI��� 6ѩ� ��� У 6ѭ����� 6ѩ� �� ѩ� ѩx� L!�`�-����������C��� � �ϭ�����
��
�����C��� �i ��`��������� �
���� �C�� ��`�� �������
 ��`���� �� �� � �ѩP� �� �  ��H� � �ѭ������� �ѩP� � �� �ѭ������� �ѩ� ��`�����C��� � ��`�����T��� � ��`�� �C������ ��`�� �]������  ��`���� �� �� �ҩ� �2� �  ��H� � �ҭ������� �ҩ� � �� �ҭ������� �ҩ2� ��`�,�������� �
���� �C�� ��`������� �
���� �C���� ��`M���������?� ���>�p������m�¶^�����ָ޹F�H���: �� �� )ܭ͎ � ֭͏ � ׭�� ���8�"��" �߀�h`�
 �	�:�; �ɢ �
 � �� ��� ��$ � ��
  ����	��� �� B�`� 8�@��$ 8�A�2��0.� �0�� !i��� 08�����0	� �Ӏ���w `�
�
�	8���	�w ���i
��7 � ������������}z��m �}���m �}���m �`� �w ���L�8�d�01�����m � �w 8�d�+�0� �0� թL���0���	��m � ��E�0�����m � ��-�	0�����m � �	��m 8�� �����

��N�� ȹN�� � ��0�(	�w � ����	�LD�`�w 8�d�!$� ��@� ��@��A��@�- �9 �ڀk� �3�������C �3�� �m �G����C �3�� �m �1�������^ �!0ͩ� �m �����^ �!0ͩ� �m `�, �C��# �B0���<`��=� �$ �A�0�
� �@�0�=��	���=` �թ#� �/��D�=�
�� �`�� ���L׭���'�$��� �0Ύ Ύ ��� ��Ύ ���� ��&8�� � ���7 8�� � ������>�8���7 8�� �����
��8���7 � � ������� �� 0S�,O�
�	8���	��
��	؍ �	؍  �����#�$���0���0
���� �  0�`�� ���Lح���'�$��� �0Ώ Ώ ��� ��Ώ ���� ��&8�� � ���R i� � ������>�8���R i� �����
��8���R i� ������� �� 0S�,O�
�	8���	��
��	؍ �	؍  �����#�$���0���
���� �  0�`������6�� �s�
��N�� ȹN�� �� ������� �� �/�$�$�$�$� �� �� ���� �� ��� �� ���`  �@���@��A�@�- �9 �ڭ$�X�8��)�8�@���@�- �9 �ڀ�A�@�- �9 �ڀ�8 ڭ� ��Ύ ���� �� ��Ώ ���� � �. �. ݼ��� �� ��$ �� �. �:�;�
���ٍ 轼ٍ ����. �. ��� �� ��$ �� �. ��	�ڭ- �0_8��- �� �  �ɍ���"�>���>��� ��� � �����<�'� � 9��� 
��� ���� ^� �`��������������	"
	%	#
	%&
	.!	8#
�P�ݖ��)�P� ��� �:�; �ɀ�$ � �:�; �ɀ�P�Q�ݞ���Q� ��� ��% � ��Q�R�ݦ���R� ��� ���& � ��R`


(���9�
�� �9��9��� �9`�#
����� 轀�� ��m!�!m�� 0Z� �"��#
��� ���� ȹ�� ��聍 ȹ聍 �
��� ȱ� ������ � 5� ����7 �#
����� 车�� ���m!m�R �+N� �"��#
��� ��Z�� ȹZ�� ��4�� ȹ4�� �
��� ȱ� ���� 5�`� � �"���7 � 0i���� j��R �, �� �"��,8����� j���`ڮ�ˁ)�� 8�� �m��ˁ)�ɀ������M� �^��!m�0�8���� � � j�#
����� 车�� ��m!mi�,� �,8� �� � j�����L*ܜ�`�� �� �
�����
��� ����
������� ����N�� �N��  ��`�� ���M����F�� �B�6��8���L���M�E�N
���ލ 轘ލ �� �J����K ��L ޭ����M���D�X �08���L���M�F�N
���ލ 轘ލ �� �J����K �� 0�K���D�= ����L���M�G�N
���ލ 轘ލ �� �J����K �� 0�`�N���j�L��M��N
���ލ 轘ލ �J� �K� ��N� ���E�/���E�&����G�����G�����F���F���N`��ɭ���#�8��6�
�Lz�����9�3� ��4�
�5� �L��LD߭5�0*��j�4�0��_�3��L�߭5��
�4��L�߭3��#�3�3�6���$�
l�3���3�3�]�4�	��3�4�N�5�3�4�C�3�0�3�3�4�4� �
��3�4�#�5� �i�	�4��3�5���4�3�5�,�5��4�������4������ �3�4�5�"� ����D�5 ��4 ��3 ��`�� �!��D��  �b� w뭂  �c� w뭁  �`�- �0��  �����V��� �M�����������������H��� �����
��m�� ȹm��  ��`(�x�ȕ�� � �
�$� ���� `�  	����2�  	����s��6��$�
��$�6�w�0��$�l�$�g�6�$���$�V�#)�
�7���$�7�?�7�:��$�1�$�$�)����$�$���6��$�0�0��$��$ �`����� 0��� � &�'�����0��������� ���� �  	����(�� ���(�����������4�  	����(�� ����������(������� � �� �� ���� A��� �� �� `�� �� L������?�$��	4������ �ۭ�����0��
����� �G�$�0��<���� �� � �)������0��������� `H�Z������ ��(��������0������0��؀ 9�z�h`�  	����� �6�$�#+i�$��$�0
�$��6��
�6�
�$�� 0�`� �6�$�#i�$`�����#�8���G����#�8���3�� �#���"�
��#�i����#�i�`H�Z�����!L��L���0���K���0����<�6������+���$�0 �������6��
���0� 
�z�h`����
�#�i������#����	�#�i�`H�Z���#����Z�����K������<�6����0���+���$�0 ���0�����6��
��� ��z�h`�����#�i������#�����#�i�`H�Z�����%��`���0����N���0�����<�6������+���$�0 �������6��
���0� ^�z�h`�����#�i���3���#���"�
��#�i����#�i�`H�Z���)����`������N�������<�6����0���+���$�0 ���0�����6����� �z�h`���0�1��#���2��0��#�i�����#�i�����#�i�`H�Z� ��
� ��)� ��� �-���
�
�����
� ������z�h`H�Z��	� ��
�� ��)� ��� ��-�����(�� i(� � i � ��
�
����Ŝ
� ����Ф�	�z�h`H�Z� �	��
�� ��)� ��� �������(�� i(� � i � ��
�
����Ɯ
� ����Х�	� z�h`H�Z� �	��
�� ��)� ��� ���Q����(�� i(� � i � ��
�
����Ɯ
� ����Х�	� z�h`� �� �+�'�,�(�)�%�*�& ��`�� �� �/�'�0�(�-�%�.�& ��`� �� ��'�H�(�	�%��& ��`H�Z�'��(��
�� ��)� ��� ��-�����(��� i(� � i � �
�
�%���Ŝ
�'����&Фz�h`�� �0� �
��]� �]�i�� � �����+��@��� i@� � i � � i@� � i � � ��`�   �������� � � �
���� ���i�� � � ����(���� i(� � i � � i(� � i � � ��#��`��~^>/�#�)H�Z�+� �,��)��*�� � ��  ��z�h`H�/� �0��-��.��� ��  ��h`�� �H��	���� ��  ��`H�Z�P� �� ���� ��z�h`H�Z����  �� (� ,�� �� �� ��  o��� �4�� �D 9��)��&  I� /�  	��� I� /� �� �� ����� �� ��  ���� �4�� ��D 9��������z�h`H�Z�  	���  �� /� _� ���Hz�h`H�Z� �@� � � � ����� ���z�h`H�  ����h`H�Z
���� 轭� � ��$� �a��b��c��d��e�8�7� w�Ȁ�z�h`H�Z� ���O� �D
��)� �)� �D� ������������� ��a��$��b��%��c��&��d��'�e��(
��� ȱ�  ��� � � z�h`H�Z)� w�z�h`H�Z�)�JJJJ� w�)� w�z�h`-��v���������Ʀ֦�����&�6�F�V�f�v���������Ƨ֧�����&�6�F�V�f�v���������ƨ֨���J�h�����¥����:�X�H�




�
��)
�& �h`PAUSE$PRESSaSTART$aTIMEaa$aRANKINGbaa$TRYaaAGAIN$FIRSTaRACE$SECONDaRACE$THIRDaRACE$FOUTHaRACE$FIFTHaRACE$SIXTHaRACE$SEVENTHaRACE$EIGHTHaRACE$CONGRATULATION$DISQUALIFIED$adabadabad$DRAWINGaBYaBANYONG$MUSICaBYaXIAOLIWAI$PROGRAMMINGaBY$XIECHENGWEN$eBONaTREASURE$�������������������+�7�F�S�^�q����  0@P`p��������  0@P`p��������  0@P`p������������������������������������������ 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P����@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^______� �� �� ��  (� ,�� � � � � � � � �* �� �� � ���� �� `�� ���%�� � (��� � �� �  ^�� �� ͸ � �� ���%�� � ,��� � �� �  ���� �� �� � n� ���X�� ����� � (��� � �� �  �� ����� � ,��� � �� �  ��� �� ͜ � ��� �� ͪ � ��� ��� <� ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��&��� �&��� �� )0�� ȭ� �	������� Ȍ� �� �� �� � �Lm�  X�� ��� � ��� ��Ȍ� �� ���� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��&��� �&��� �� )0�� ȱ������ Ȍ� �� �� �� � �� �� � �� )������ ��  n�`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��&��� �&��� �� )0�� ȱ������ Ȍ� �� �� �� � Ы� �� � �� )��@К���� ��  ������ ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��&��� �&��� �� )0�� ȭ� �	������� Ȍ� �� �� �� � Х��  v�� ��� � ��� ��Ȍ� �� ���� 
������ ����� �ݍ� ȱݍ� `�� 
������ ����� �ݍ� ȱݍ� `H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����΢ �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����ΰ �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� ����� )@��J��� �� �� �8��� ��� )0�� Ȍ� �����ξ �� �� �� � z�h`H�Z�� )?	@�� �� I��-� �� �� �Ȫ�� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� � z�h`� `� `�� ����  <�`H�Z�� ���%�� ���� �� �� )?
������ ����� ��  y�z�h`�� �* �� `�� ��� ȱ�� ȱ�� ȱ�� )
��&��� �&��� �� )0�� Ȍ� �� �� �� � o��� `H�Z�� ���Lh��� �� �� I�� )��� �� �Ҫ�� )@��J��� �� �� �8��� ��� )0�� Ȍ� ������� �� �� �� )�� �� )����
�@����� �� �� �( �� �� ��* �� �� �� �� � y�z�h`H�Z�  X�  v� �� ��� ��  �� �� �� �� <����� z�h`H�Z�� � �
�� � ��� �� )?�� �Q�� �K�� 
����� ���� ���� ���� �� �� � �� �� �� )������  n�� ����  �� <�z�h`�6���� ���F� �� ��  o����� �� �1���� �� ����� � ��� � �����  �������  ��� �� ` ����� ���� ���� ����� ���� ���� �`��� ���� ��� _���� ����� ���� ���� ����� ���� ���� ����� ���� ���� �����     � ���� ���� ���� 0��� ���� ��� ���� ���� ���� ����� ���� ��� q��� �0��� ���� ���� ���� ���� ���� ���� ����� ���� ����     � �0��� ��� ���� q��� ��� ���� ���� ���� ���� ���� ���� ���� ���� ɐ��� ���� ���� ���� ���� ����(���P��� ���� �0��� �0��� �0��� �`��� �0��� ���� ���� ���� �H��� �0��� ���� ���� ���� `���     � ���� ���� ���� ���� ���� ���� ���� ���� ��� ���� q��� ��� d���� �H��� ���� ���� ���� ���� ���� ����� ���� ���� ���� ���� ���� �����     ��0��B�0���0��B�0���0��B�0���0��B�0���0��B@0���0��B�0���0��B�0���0��B�0���0��B�0��     � � ��� ���� ���� � ��� � ��� �@��� � ��� � ���� ���(���(��� � ��� ��� ɀ��� � ��� ���� ����  ��� � ��� d���� d ��� K��� K��� ? ��� C ���     � 2���� d ��� d��� d��� d ��� K ��� dT��� d ��� q ���  ��� ��� q���  ��� � ��� � ��� �`���  ��� ��� q���  ��� � ��� d ��� �`���     �� ��J! ��
� ���! ��
� ��J! ��
� ���! ��
     � �?� �
7� �
7� �?� 7� �7� �(?� �?� �
7� �
7� �?� 7� �7� �(?� �(?� �(7� �(?� �(7� 7� �7� �7� �7� �P?�     ����
���
���� �����(����
���
���� �����(�\(��(��(��(� �!����!���(��(�     � ��     � ��     � _(��     � _(��     � �
�� /d��     � �
�� �
�� 
�� ?
�� �
�� ?
��}
�� 
��     � �
�� �
�� 
�� ?
�� �
�� ?
��}
�� 
��     �     �     � 1<	 0<� /<� .<� -<� ,<� +<� *<�     � *�	     ���;�^�e�p�w���������������� 8�d�<    & � �� � �_ �O �o ��     &�����_�O�o�   ��   �
�/�   o<   �_v�Ovq�v   p�< p�< p�< p�< p�< p�<     & �� �O �o �� �� � ��    (�(�    ����_ �O�o�    $ �     $ �    
	 �
		

		
 �
	�
�



	�
�
	
	 �
	
	
	�

		�
	���������
�g���u�S�  ��  g��  ��  ��  Y�  ����1���������g�������.�>�H�|���������                                                                                                                                                                                                G� ���