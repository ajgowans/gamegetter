           �?             �        �?      ��    ��     �?      �:        ��      ��   ���    ��     ���       ���     ��;   ���    ���   ����       ���      �~   �z�    ���   ���V�      �z�      �W   �ZU   �z�   ���U�      �ZU     �U5   �^�    �ZU �j�U�      �^�      �U    _�    �^�  ��Z�W�       W� <    �U    {=     _�  ��U9�       ��= �    ��   ��    �{= ��ZU         ����   �:    ��    �� ��V�          ��p5   \��    l�   �� �oU�          �Z_  �W��    \�   pm� �V�:          �V�U  pU���  W�   \k� �U�          �VU�   \ժ�_ �U�   \Z� |��?         ��ZU5   \��zU p��   �Z��W���        ���_   \��Z� \��    �V�WW�W=        ����   \���  |U�    �VUU�WU}�        ���     \��   �_U   �^U� \U�W       ��?     \��    ��W   ���  �WU]       ���     \��    ��   �    �Uu5       ����?   p��    ���   ��     _��       ���U�   ��    ��    ��     �շ      l�~UU  ���    ��   ���      W��      l��jU  ���    �_   �ת7      \��     lU��U  ��W   �U    W��      ���     [U��   g�U   �U    W�f     ��      [� ��  ���U   �W   �U��     ��      [� �5  pfW5   �W   �U�f      �      [5 � ���\5  ��W   pU�             �V5 � �f> p5  ��W   _� l             �U � �� p  ��U  �U5 �             lU � �?  \  ���   �U g           ��[U �� �  \  �p�   ��  �            ��V�  ��  _  �p5   �? ��            �n�   � �  �   ?|   � �?            ��?      � ��   �   � ��            �          ��  ��   � ��           �           ��>  ��   � �           ;            ��   �:       �                       ��   �?                                    �?          �       � �VUU�VUU        ���         �     ���ZUUUZUU       𿪪        ��     ���jUUUiUU       \���      ����   ����U�UUU�UU       [eU�     ���j�:  ���z�?U�V��VU      �Z�U�     ���Z�:  ���Z�?U�ZU�UZU      �jU�     ���Zu;  ���Zu?U�jU]WiU      ��U��     ���U}�< ���U}� UU�UUU�U      ��zU3     ��Z��?  ��Z��? UU�V��V      ���_     ��U�    ��U�   UU�ZUUUZ      ����     �jU    �jU   UU�j��Wi      ��:       �V�    �V�   UUU�UUW�      ��?       kU�    U�   ����V�U�      �����    [��5    _��5   ����Z��U      ��zUU=   �W�~�   �W��   UUU�jUUU      ��^UU�   pU�oU  pU�oU  UUUU�U�_      ��^��U  p�Z�U  p�Z�U  UUUU�VUU      [ծ��Z  ��o�V  ��o�V  UUUU�Zu�     �VU� o5 <  �U[    �U[  UUUU�j�}     �V�   ������kU[  ��kU[  UUUUU�U_     �U5   �o�:�V�l  �V�l  UUUUU�VU    �U    ��_U?l  �_U?l  UUUUU�Z�   ; lU     � ��� l  ��� l  UUUUU�jU  ���[�      < �  �   �  �   UUUUUU�U  �zUU5        �  �  �  �  UUUUUU�V  ����        �   �>  �   �>  UUUUUU�Z  �               ��      ��  UUUUUU�j  <                �?      �?                        ��                     ��     ���   ���    �� 0  0         ���      ��?   ���    ��� 0          ��?      ��   ���    ���  �          ���      �   ��    ��� 0|3�         ��      �W   �_U   �� �[ݕ�         �_U     �U5   �_�    �_U�UVf=          _�      �U    _�    �_�  geY�          W� <    �U    {=     _� �            ��= �    ��   ��    �{= ��            ����   �:    ��    �� ��*           ��p5   \��    l�   �� � �
          �Z_  �W��    \�   pm� � ��         �V�U  pU���  W�   \k� 8  �         �VU�   \ժ�_ �U�   \Z� 9   �*       ��ZU5   \��zU p��   �Z��    �      ���_   \��Z� \��    �V�    �      ����   \���  |U�    �VUU:    �9      ��     \��   �_U   �^U�8    �9      ��?     \��    ��W   ��� �    ��      ���     \��    ��   ��  �     �      ����?   p��    ���   ��  �
   �     ���U�   ���    ��    ��  ��  �     l�UU  ���    ��   ���  ����  h     l��jU  ���    �_   ���7  ���* h     lU��U  ��W   �U    W��   � �
�9     [U��   g�U   �U    W�f  �  ���9     [� ��  ���U   �W   �U��  �   ��     [� �5  pfW5   �W   �U�f  8    ��     [5 � ���\5  ��W   pU�  8     ?    �V5 � �f> p5  ��W   _� l ���?��      �U � �� p  ��U  �U5 � \]}�UW     lU � �?  \  ���   �U g ��w���   ��[U �� �  \  �p�   ��  �  \_}���   ��V�  ��  _  �p5   �? ��  ��s���   �n�   � �  �   ?|   � �?  W�p�UW   ��?      � ��   �   � ��  �0�?��    �          ��  ��   � ��           �           ��>  ��   � �           ;            ��   �:       �                       ��   �?                                    ��    �WUUUUUUUUUUUUZUUUUUUUUUUU       ��   ]^�������UUUUUiUUUUUU�����     ����   ]^�ffffffUUUUU�UUUUUUfffff     \���   Wy�������UUUUU�VUUUUU�����     [eU�   WyujfffffW�UUUUZUUUUUfffff    �Z�U�   UUթ�������WUUUiUUUUU�����    �jU��   ����fffffuUUUUU�UUUUUfffff    ��U��   ���������UUUUUU�VUUUU�����    ��zU3   wUUujffffUUUUUUUZUUUUfffff    ���_    �UUթ����UUUUUUUiUUUU�����    ����    uWUU�ffffUUUUUUU�UUUUfffff    ��:      �]UU����������
UU�VUUU�����    ��?      UwUUujfff�����
�������fffff    �����   U�UUթ���UUUUU������������    ��UU=   UuWUU�fffUUUUUUUU�UUUfffff    ��_UU�   U�]UU����UUUUUUUU�VUU�����    ��_��U  UUwUUujffUUUUUUUUUZUUfffff    [կ��Z  UU�UUթ��UUUUUUUUUiUU�����   �VU� o5 <UUuWUU�ffUU�_�UUUU�UUfffff   �V�   ����UU�]UU���UUU�UUUUU�VU�����   �U5   �o�:������zjfUUU]_UUUUUZUfffff  �U    �������꩙UUUu�UUUUUiU����� ; lU     � UUUU��U�f      UUUUU�Ufffff���[�      < UUUUu�W��      UUUUU�V������zUU5        UUUUu�Wuj      UUUUUUZfffff����        UUUUUUUթ      UUUUUUi������           UUUUUUUU�      UUUUUU������<            UUUUUUUU]             UUUUU             UUUUUUUU�             �����                                                                                                                                                                                                        � ݆ `� ݆ `� ݆ `� ݆ `� ݆ �� ݆ `� ݆ �� ݆ `� ݆ `� ݆ `� ݆ �� ݆ �����> T > @  > O > @  > � > W 	> � > @  > Q > O B P C G B Y > ; %< U < @  < M < @  < � < Z < � < @  < X < P B ] C ? !B _ < V 
> Q > @  > Y > @  > � > T > � > @  > Q > O B M C O B _ > V 
< Y < @  < S < @  < �  < Z < � < @  < J < Y B E C D B ] > F 7 Z 7 @  7 @  7 [ 7 � 7 @  7 � 7 V 
7 P 7 @  7 _ 7 @  7 [ 6 [ 5 [ 5 @  5 ^ 5 @  5 � 5 [ 5 � 
5 @  5 \ 5 @  5 O 4 N 5 R 4 J 7 T 7 @  7 [ 7 @  7 �  7 Z 7 � 7 @  7 H 7 @  7 W 	7 @  7 T 7 L 5 ] 5 @  5 \ 5 @  5 � 5 ^ 5 � 5 @  5 Y 5 J < X < @  < s M����B N C N J @ �J F zJ I H � ,G G yH C }J K uB K C \ J L tJ K uL O J KB J C T J L tJ = �J G H G O qH ] cJ H xB M C > "H V jH i WG V 
C� �> V 
@ Q C ^ bC q O@ 5 +F � E S C C }C Y @ S C I w> ^ @ _ C < �C F zE W 	C [> Y @ H C ; �C G y@ 2 .F � E N C N rC O @ E C O q> ^ @ T C 8 �C F zE S C� �                                                                                                                                                                                                                                                                                                                              �?   �   �                 UUUU        ��   \  \          �      UUUU        ��  \  \          �     UUUU       ���  \  \          h     UUUU       �Z� �_ �_ �?�  ��� �9     UUUU      ��V� �^��_ ��� ���� ��     UUUU     ���V���^��_���� ���� �    UUUU    𪪪~5��[��[���\���\�h    UUUU    ����� �zV�V�z�\��\�9    UUUU   ��j�  �������ZU_�_U_��    UUUU   𪪪�   ��� ��� �^�p�_�p� �   UUUU   ����W   o�  o�  _�p _�p� h   UUUU   ׫�?W   [=  [=  {=\ {=\� �9   ����  �U��\  �V �V ���W���W� ��   ����  pU�5p  �V �V �VUU�VUU�  �  iUUU  _U�W��5  �U �U �UU� �UU� �  h  �UUU �U� |��5  ��: ��: �V� �V� �  ��  �VUU<_U _5 �  ��: ��: �Z:  �Z:  �  ��  UZUU�U� �U �  ��: ��: ��:  ��:  �   �  WiUU�� |�  \ ��: ��: ��:  ��:  �   �  ]�UU�?  �  \5 ��: ��: ��:  ��:  �   �  U�VU� ��  �� �� �� ��  ��  ��: �  �UZU� ���   � �� �� ��  ��  ��� �  uUiU�  �?   ��� �� ��  ��    ��  �U�U         ? �� �� ��  ��    ��  ��V        �� �� �� ��  ��     :�  UUUZ        ���� �� ��  ��     ��  UUUi       ����� �� ��  ��     ��             �_��� �� ��  ��     ��            ��W��U �U �U  �U      �           ���V�pU pU pU  pU      �          𪪪~5�U5 �U5 �U5  �U5      �         ����� �V5 �V5 �V5  �V5      �        ���j�   [�  [�  [�   [�      �:        �����    [�  [�  [�   [�      ��        ����W   g�  g�  g�   g�      �       ���?W  �Y5 �Y5 �Y5  �Y5      ��      �U��\  �Y5 �Y5 �Y5  �Y5      ��      pU�5p  pV pV pV  pV               _U�W��5  �V �V �V  �V              �U� |��5  ��  ��  ��   ��              <_U _5 �  �5  �5  �5   �5              �U� �U �  �  �  �   �              �� |�  \ �  �  �   �              �?  �  \5 ��  ��  ��   ��              � ��  �� �� �� ��  ��             � ���   � �� �� ��  ��             �  �?   �                             ����������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������������������������������������������������ffffffffffffffffffffffffffffffffffffffff����������������������������������������ffffffffffffffffffffffffffffffffffffffff����������������������������������������ffffffffffffffffffffffffffffffffffffffff����������������������������������������ffffffffffffffffffffffffffffffffffffffff����������������������������������������ffffffffffffffffffffffffffffffffffffffff����������������������������������������ffffffffffffffffffffffffffffffffffffffff��������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��������������������������������������������������������������������������������UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU������������������������������������������������������������������������������������������������������������������������H�w�j�Ņkhdd �� kͩ  ۥd����i`d>d?dIdJdKdAdXdY��EH�q���h�_�E��H�����h�m��BH����hH��� �h ��H�����h�m�E��H�q���h�_��<H�$���hH�(�� �h ��d=H���L���MhdPH���N���OhdQH���R���ShdVH���T���UhdW� � ��*��+ �� ��H�ͅ&�ƅ'h�(�  �H���&��'h�h� ��H���&��'h�`� �ȢT �� o� �� ��H����h !�H�$���h !�H����h�E��
H�$���h 	�H�$���h�E��
H����h 	� �� W� � �͢,�P��*��+ �֢4�XH�҅&�ƅ'h  �d5 wʰ_�4�XH�څ&�ƅ'h  � wʰI�4�XH��&�ƅ'h  �xH�#��΅ hX�^�"d#d$d%dA��5�
�6��8��7��]��:��;d9�� ۢ<�x�� �� � ���dL�d!dCdD o� �� �ѥ]�"�]�,�P��*��+ �֢4�XH��&�ƅ'h ԥX� �(�P��*��+ ��H��&�ƅ'h�0�X ԥY� �$�P�	�*��+ ��H��&�ƅ'h�,�X � :�H�Ce>�>�De?�?h %� ��H����h�E��
H�$���h 	� ��H�$���h�E��
H����h 	� �ѭ  I�ɀ� ʭ  I������i` �� ͥX� �(��$ �Ӣ@��#�i�d��8� �ҥX�;�$�,HH�����h�E��H�����h��B��7��8h:�X�L�L,��Y�:�Y�L�L,�� 8�^�!���&8�r�'��)L,��)�Xd\�$�[�#�Z�(��[ �Ӣ@��Z �� ��L,�H���$��%h�E��H���$��%h�"�Y��;��<L,�d\�$�[�#�Z�$H� ���h ��H�����hH�����h � �� ��`�B��L߷� �L���8� �ʥ7J�8�L��:�8�L�� �ʥ7�8H����h !� �� 9�H� ��!�hH�L��M�hH�P�� �h�E��H�R��S�hH�V�� �h gХG����EH� ��!�hH�N��O�hH�Q�� �h�E��H�T��U�hH�W�� �h gХG�(����BH�����h�E��kH����h�]�F��`�A�\dA�7���R�G�#��BH�����h�E��8H�ٍ��h`��BH�����h�E��H�č��hd8�(�6 0�`dA�8�:�8���7J�8H����h !� ���F��ة �BH�w���h�E���H�����h`�8:�8Ю�7�8H����hL!�H��C� �Dh�8�70HeC�C� eD�Dhm � � m!�!`�<��L��� �Lt��:� �ʥ;�:� �Ls�:�:�Ls� �ʥ;�:H�$���h !� ɹH�&��'�hH�R��S�hH�V�� �h�E��H�L��M�hH�P�� �h gХG����EH�&��'�hH�T��U�hH�W�� �h�E��H�N��O�hH�Q�� �h gХG�(����<H��$��%h�E��kH���$��%h�]�F��W�=�Sd=�;���I�G�#��<H�ٍ$��%h�E��/H�����h`��<H�č$��%h�E��H���$��%h`d=�:�	:�:���;�:H�$���h !� ɹ�F��ک �<H���$��%h�E���H�w�$��%h`H�$���hL!ϩ8�;0m&�&� m'�'`H���j�Ņkhdd �� kͩ  ۥd����i`d>d?dIdJdKdAH����hH����h�[H�6�� �h �Ω�B� � ��*��+ �� ��H�Ņ&�ƅ'h�(�  �H�*�&�Ʌ'h�h�  �H������h�p� P�H�,�&�Ʌ'h�`�  �H������h�p� PҢT ��xH�#��΅ hXdA��5�P�6��8� �7��^d!dCdD �� � �� �� U�H�Ce>�>�De?�?h i�H����h 	� ˭  I�ɀ� ʭ  I������i` �� �̥A�)� 8�Z�!��� ۢ<�x�� �� � ���dL�LǺ�7��6�8dAH�����hH����h !� �� � �� ��H����h 	� /�d�Z8�^�H��� �h �Ӆ
em�� m��P8�8JJJJ�8d]dBd!dCdD �� � �� ��H����h������������������������������H���h������C�]����8� eC����C�Ce�� e�����e�H���h���H���h���H���h���������������H����h��H���h����B�H�Ce>�>�De?�?h i�H����h 	Х]���H�$���h 	Э  I�ɀ� ʭ  I������i` �� ���]�]0c�d��H�[���h�"�g�J�H��8���]��BH�v���hH� �&�!�'h�m&�&� m'�'�"i�(�b�) 0�LŻ� 8�^� �!��!�L/�H� ��!�hH����hH�e��e�hH�e��e�hH�e��e�h�JJe�� e��^8�0��08�^��18�
e�� e�H��_��`h�(� P� ��H�_�a�`�bha&bH�_ea�a�`eb�bhH�����hH�����h �� �� ��`�8� �ʥ7J�8�L�:�8�L� �ʥ7�8H����h !ϩڮ � �8� � �!�!�!�!��B�0 9�H��C� �Dh�8�70HeC�C� eD�Dhm � � m!�!�F���B�H�w���hdB`@ p�^v\�v]�v]�v]�v]�v]�v]�v]v]"v]6v]Jv]^v]rv]�v]�v]�v]�v]�v]�v]�v]��
 �a: �_��_�_$�_A�_^�^~�m��� ��V�����r�� ����������8�������� k�y �������� {���,��������������������������������µ�������������������������������     0       0       0       0       �     �       �       �       �   =    <     �       �       �       �   =  �    �    ��     ��     �   =  ��   ��     ��     �#     �  T=_���    �#     �#     �     �  �?����   �#     �     �     �  ����   �     �     �      �    �  \�;�  ��    ��    ��    ��  ��w���  �����   ����+   ����   ���� �?�����  ����   ����   ����   ���� T=_w���  ���   ���   ���   ���#  = ���  ��    ��    ��    ��   =   ?   ��    ��    ��    ��   =       ��#    ��    ��#    ��          ���    ��#    ���    ��            ���    ����    ���    ���            ���    ���    ���    ���          ������������           ���?            WUUUUUUUUUUU         �������                              ���������                             ���������                           𪪪�������                           �����������?                         𪪪���������                        �������������?                       ���������������             0         ���������������            �         ������WUU������?            �        ������UUUUU������          �       �����WUUUUUU�����         �       ����UUUUUUU�����         ��       �����UUUUUUUUU�����         ��       ����~UUUUUUUUU�����        �        ����WUUUUUUUUUU����       ��/       ����UUUUUUUUUUU����       �����     ���^UUUUUUUUUUUժ��?       ����     ����WUUUU��UUUUU����       ���     ����UUUU����UUUU����      ��/      ���zUUUկ����_UUU����      ���      ���^UUU�������UUUժ��      ���      ���WUUի������_UUU���?      ��    ����UUU��������zUUU����      ���     ���zUUU���������WUU����      ���     ���zUUժ��������^UU����     ��0     ���^UU����������zUUժ��     ��      ���WUU�����������UUU���     ��      ���WUU�����������WUU���  ������������ ���UUժ���_Uկ���^UU���?  ������������ ��zUU����~UUU����zUU���?  ���������������zUU����WUUUU���zUU����  ���������������zUU����UUUUU����UU����  ���������������^UU���^UUUUUժ��WUժ��  ���������������^UU���WUUUUUU���WUժ�� ���������������WUժ��UUUUUUU���^UU��� ���������������WUժ�zUUUUUUU���^UU��� ���������������WU���zUUUUUUU���zUU��� ���������������UU���^UUU�WUUժ�zUU��� ���������������UU���WUU���UUU��zUU��� ���������������UU���WUU���WUU���UU��� ���������������UU���UUժ��^UU���UU��� ���������������UU���UU����zUU���UU���? ��������������zUU���UU�����UU���UU���? ��������������zUU��zUU�����WU���WU���? ��������������zUU��zUU����WU���WU���? ��������������zUU��zUժ� ��^U���WU���? ��������������zUU��zUժ: ��^U���WU���? ������������
��zUU��zUժ: ��^U���WU���? ����  ��  ��zUU��zUժ: ��^U���WU���? �� ��  ��0 ��zUU��zUժ� ��^U���WU���? �� ��  ��; ��zUU��zUU����WU���WU���? �  �  �~� ��zUU��zUU�����WU���WU���?       �WW��zUU���UU�����UU���UU���?       �U�� ���UU���UU����zUU���UU���?       �U}5 ���UU���UUժ��^UU���UU���       ��W ���UU���WUU���WUU���UU��� �  �  �_U ���UU���WUU���UUU��zUU��� ����  U�  ���UU���^UUU�WUUժ�zUU��� ����  _U=  ���WU���zUUUUUUU���zUU��� �  � �^�  ���WUժ�zUUUUUUU���^UU���      �^�  ���WUժ��UUUUUUU���^UU���      ���  ���^UU���WUUUUUU���WUժ��      ���  ���^UU���^UUUUUժ��WUժ��       ���  ���zUU����UUUUU����UU����  �  � ���  ���zUU����WUUUU���zUU����  �� ��  ��    ��zUU����~UUU����zUU���?  �� �� ���    ���UUժ���_Uկ���^UU���?  ���� ���    ���WUU�����������WUU���       ���   ���WUU�����������UUU���       ���   ���^UU����������zUUժ��       ���   ���zUUժ��������^UU����       �^�   ���zUUU���������WUU����    WU;�  _�   ����UUU��������zUUU����   �U�:\  Wy    ���WUUի������_UUU���?   �U�:W5  W]    ���^UUU�������UUUժ��   �U�:W5 �U_    ���zUUUկ����_UUU����   pU�W5 �UW    ����UUUU����UUUU����   pU�\ \�\    ����WUUUU��UUUUU����    pU�� W5\5     ���^UUUUUUUUUUUժ��?    \U�P�Up5     ����UUUUUUUUUUU����    \U��p� p5     ����WUUUUUUUUUU����    \U�m|= p5     ����~UUUUUUUUU�����    WU� m� p5     �����UUUUUUUUU�����     WU� �� p5     �����UUUUUUU�����>     WU; �� �     p�����WUUUUUU�����:     WU� P� �     pժ����UUUUU������:     WU�   �  �;     pU������WUU������W;     WU�      ��     \U���������������U�     \U�     ��    \U������������^U�     \U�     ��    \U믪�����������_U�     \U�            WU�𪪪���������_U�    pU�            WU; �����������?pU�    pU�            W�: 𪪪�������pU�    pU�           �U�:  ���������? pU�    �UU;           �U�  ���������  �U�    �UU;           �U�   �������   �U�                   pU�     ���?    �UU;                         ���� ������?��?��             �?      UUUU ���������?��        ��   ��  ��  UUUU ���������?��    �  �� ��� �� UUUU ? �����  ?�   ��:  �� ���  �� UUUU ? �����  ?�   ���  �W �^7  �_ UUUU ? �����  ?�   �~5  {�  �Z�  �� UUUU ����������   ��  ku �_�  �� UUUU �����������   �V7 �U l]5  �U UUUU �����������   �W5 �u�  [u  �W UUUU  �����?�  ?�   [W l�5  _�   � UUUU  ���� �  ?�  �V] t�  w� �W�  UUUU  ���� �  ?�  �W=  �� �ծ �U�  ���� ������ ��??�  �]�  W� p�� pU�  ���� ������ ��??�  p�� �կ \�� \��  UUUU ����� ��??�  \�� @ժ \�� \��  UUUU                 T�� p�� \�� \��  UUUU?������� ?    W�� p�� p�� |��  UUUU?��������?�?    W�: �� ��  ���  UUUU?����������?    ߪ: ��5 ��z ��:  UUUU?��� ����?    �� ��5 �� ��;  UUUU?��� ����?    �� ���5 ��� ���  UUUU?��� ����??    �� ���� ��� ��j UUUU?���������??   ���: ���� �� ��j UUUU?����������?   ���: ���? ��� ��� UUUU?���������?   ��� ��^ p�^ �׺  UUUU?�� ������?   �W}5 p�W p�W �U�  ����?�� ������?�� �U]� pUW p�W �U_ ������� ������?�� pU]� pUW p5W �UW UUUU������������?�� pUs� �UW \5\ �UW UUUU���������?��?�� \�pU�UW \5\ p�W UUUU�?������� ?�� \5�U���  \5W p�\5 UUUU                \5�Up��  \W \5\5 UUUU                W�U\�5  \W \p5 UUUU                W W\u  W��  \p� UUUU               ��  WW}  W��  W�� UUUU               �5  WW�  W��  W�� UUUU               p5  \׿  W?  � �� UUUU               p  \��  W��  �  7 UUUU               �  ���:  ��� � � UUUU               �  �:��?  �� ���UUUU               �  ���   �� ���UUUU               �  ��     �     ��UUUU               H���j�Ņkhdd �� k�dXd_d`�  ۥd����i`xH����΅ hX� � ��*��+ ��H�*�&�Ʌ'h�x�  �H������h��� D�H�,�&�Ʌ'h�p�  �H������h��� D�H���&���'h�0�  Ԣ(��X @ӢH�	�� ��H�_��`�h�H� :� �ɢd �� ��)�J ��)�GdK ��)?i3�0 ��)?i[�1��B��8�0�] k� ���q� �j �ע �"��*��+ �֢�*�� �ץK��� �K��H�G��eJ��>�2 
ע�2�{��$8�J��<�2 
ע,�2�eK �׭  I������i`�  I���0�Le����8d8��8���8����B)�B����B)��B�B�B�8i�7�0�1�B���e7ɚ�������B���8�7�1���B	�B�1��B���8�7�+���+��B���e7ɚ������0�1�x ���]� �F��*��+ �֢�R�]JJJ �ҥ]�� ۢQ�E�� �� �� ���dL'��  I�ɀ� � �� ��L�� k� ���q� �j ��d^� �<��*��+ �֢�DH���&�ƅ'h Ԣ�L�@ 
� �� �̭  I�)0�dA�^�Z��^�^��L�^ �� �� ��L����/�r�K k� ���q� �j �ע�s�K �� �� ���K�/�ܥ^�Z�/ �͠ ZZ k� ���q� �j ��z�[�y �� ��hi������L7��G�
�0ieJ��0i8�J�4��L7�ɒ�L7��0��^8�-0
e1��-8�^
��18�i�2��L7�ɒ�L7��1�ʈ��z �� �� 0ݥ08�4�0����_8��0�18�2�1����a8��1H�ԅ���h�0e�� e��1��0e�� e���L7��(�HH ��he_�_� e`�`h�d� �3�C��*��+ �֢C�KH���&���'h  �H�_��`�h�H� :� �� �ͥX�X��L�H�_��`�h&H��a��bh&H�ea�a�eb�bhH�����hH�����h �� ��`BULLSEYE! /5 �n�3�1 �שo�9�� �שp����L��H���j�Ņkhdd �� kͩ  ۥd����i`d>d?dIdJdKdAH����hH�����h�[H��� �h �Ω�B� � ��*��+ �� ��H�Ņ&�ƅ'h�(�  �H�*�&�Ʌ'h�h�  �H������h�p� P�H�,�&�Ʌ'h�`�  �H������h�p� PҢT ��xH�#��΅ hXdA��5�P�6��8��^d!dCdD �� � �� ��H����h !�H����h 	Э  I�ɀ� ʭ  I������i` �� �� �� �� �� �ͥA�)� 8�M�!� �� ۢ<�x�� �� � ���dLʝL��dAH�����hH����h !� �� � �� ��H����h 	� /�dA��5�P�6��] �� � �� ��H����h 	�  �H�>8� �?�!h���7��C i̩e>�>� e?�? ���]ж�6�8 �ʥ7�L�H����h !�H�$���hH������hH� ��!�h�e�� e��X �Ω��)�Z8�^)�m$�$� m%�%�
�]�8�7�X��Xd!dCdD �� � �� ��H����h 	ХG�H�$���h 	�H�&��'�hH�8�>���?�h��Ѭ(����8� JJJJiˠ� �� �� �̭(�~�L��H�$���h������������������������Ce�� e�������]��,���
ee�~���~�dG�8�0� �����GH���h���H���h���H�Ce>�>�De?�?h ^̭  I�ɀ� ʭ  I������i`�X�L&��]�L�����$8��$�%� �%��m$�$� m%�%�]L� B� �� �� �� �� �� �� �� �ͭ&8�_�&�'� �'�L�H�&��'�hH�e��e�hH�e��e�hH�e��e�h�^8�!��!8�^��"8�e�� e��P8�8e�� e�H��_��`h�(� P�H�_�a�`�bhFbfaH�_ea�a�`eb�bhH�����hH�����h �� �� ��`_ p�� ��O�����?����                                               





                                     










                                 














                              

















                            



















                          





















                        























                      

























                     




















                   

















                  















                 














                












              













             












            












            










           










          










         










        










        









       









      









      








     









     








    








    








(((((   








((((((((   







((((((((((  








(((((((((((  








(((((((((((((  







(((((((((((((( 








((((((((((((((( 







(((((((((((((((( 







(((((((((((((((((








(((((((((((((((((







(((((((((((((((222







(((((((((((((222222







((((((((((((2222222







((((((((((((22222222







(((((((((((222222222






((((((((((2222222222






((((((((((222222222dd






((((((((((22222222ddd






(((((((((222222222ddd






(((((((((22222222dddd






(((((((((22222222dddd� � ��xH����΅ hXd8d5�� ��*��+ �֢D� ��dFdG�GI�G k�H�+�&���'h�8��
H�:�&���'h��  � �ɥ8��� �����L���X��*��+ ��H�&�>�'�?h�8e>�>� e?�?d/H�I����h�d��-��.�(ZڲH�>��/�B�G�h E׀h 
��/���hi
�z�.�Әi
��-�Ģ8�,��*��+ �֢D�8 ԥ8����H�*Z 
�z���	


iD��@�* 
ע�6Z ��z�x �ɥFdF���F��"�� �ԥ5ɀ�L&��@��8�8���L�d8L��8��+ �ɥ5��������q�:��	��	�� ��[�5���B8��3i(�.���Bi�(��8�(���	�B:�'���$�B�(�� �BH�I����he�� e���>d5 ��Lf�� L�ENTER INITIALS CHOOSE COUNTRY ABCDEFGHIJKLMNOPQRSTUVWXYZ .-[0123456789�i��` �͢,� ��*��+ �֢D� �ɢ� �ɢ�� �ɢ�V��*��+ ��H�j�&�k�'h�&��&��'�b  �H���&���'h� �j  �H�*�&��'h�X�j  �H���&���'h� �x  � T��X�x  ԥi�	����� �ע�(��*��+ �֢,�8H���&���'h�i�-H�|�&���'h�,�0�i��H���&���'h� �4ژ��4  ���<  Ԣ�i��� ۭ  I�ɀ��� L�YOU HAVE QUALIFIED YOU ARE DISQUALIFIED GAME OVER SCORE: TOTAL: � �H��L� �MhH�:�N��OhH�`�R� �ShH���T�0�Uh� � ��*��+ ��H�s�&�ǅ'h�$�  ԩ�]�]�:�]�	�  I�ɀ�? k�H�L�� �h ��H�N�� �h ��H�R�� �h ��H�T�� �h �� c� �̀�� L۩�/H�H�&��'h�(Z�(Z �z�&�&��'i��Z����ZH ��hz�� ��z�P �hi��/��`��������i�ɬ�� ��)?8�����H���h�����L�Ԣ��Ɲ)���H�a��b�hH�)���h #�H�a��b�h T�H�&��'�hH���h���*���3�e3d3�:��0�3����H���h����`�e:
�&
e&H�0�&��'he&�&� e'�'`H�H���h�7�ZH����h�e�� e� T����&��)������&��'���h8���e�� e��г`H���h�h��H����h�e�� e������ ��H�&��'h�&��&���� �ɩe�� e��� T�H�&��'h�&��&����L�� ��;  X�4   �@1   ��N/< 7 ��?/P;YAAA AAA AAA AAA     DBZ  50000 ACB 32000 SML 24000 PDS 16000 PSB 08000 TTS 04000 ���  � �ȍ# � �� � � �L�ͩ � ��V�*�IӅ*�*�	d�xH�܅�΅ hX`xH����΅ hX���.��/�dH �ͥ.�:�.�H���� �h �ץ/�8��/�_H���� �h ��h:�� ȳd!��.�_�/�H �ͥ.�i�.�<H���� �h �ץ/�8��/�<H���� �h �� �ͥ!���	� �  �h:ж 
��F �����`�܍ � �� � �� � �O� � `�v� � � � � �2� � �O� � `��	@� � d!�!������� � `�΂7 ^ 2C ; U7 - 39 - 9 - 3E > R9 ( 8; - ; - 3? ( hB ) 7G + 5; ( ; ) ; , ���; - > 4 ,; ? Q7 7 )= * @ 9 '= < T9 1 /? ) B ; %? B ;  ? " B & 
G 6 �� ݆ �� ݆ �� ݆ `� ݆ �� ݆ �� ݆ `� ݆ �� ݆ �� ݆ `� ݆ `� ݆ 0� ݆ 0� ݆ 0����; r ; : = Q o> | > ? 6 � 5� ����G k I ? J l C ? O Q oN T lMY �� ݆ �� ݆ @� ݆ �� ݆ @� ݆ �� ݆ ��݆ ��� ݆ `� ݆ `� ݆ `� ݆ `� ݆ �� ݆ `� ݆ �� ݆ `� ݆ `� ݆ `� ݆ �� ݆ �����> T > @  > O > @  > � > W 	> � > @  > Q > O B P C G B Y > ; %< U < @  < M < @  < � < Z < � < @  < X < P B ] C ? !B _ < V 
> Q > @  > Y > @  > � > T > � > @  > Q > O B M C O B _ > V 
< Y < @  < S < @  < �  < Z < � < @  < J < Y B E C D B ] > F 7 Z 7 @  7 @  7 [ 7 � 7 @  7 � 7 V 
7 P 7 @  7 _ 7 @  7 [ 6 [ 5 [ 5 @  5 ^ 5 @  5 � 5 [ 5 � 
5 @  5 \ 5 @  5 O 4 N 5 R 4 J 7 T 7 @  7 [ 7 @  7 �  7 Z 7 � 7 @  7 H 7 @  7 W 	7 @  7 T 7 L 5 ] 5 @  5 \ 5 @  5 � 5 ^ 5 � 5 @  5 Y 5 J < X < @  < s M���*  B � (��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� �   �  �          �? ?         �   �� 0  �  ��      ��? ��            l5� 0  �    ��  ��?   ���    ��?�   [�� <  �      ��?     ��  �����     [�� <  �               ?         �   [�� <  �                              k�� 77  �6 ��       ��?                �:� 77  �8 ������������?              �� 77  �:              0 ��������� 0    � 77  �9              �0       0     � 77  �5               �       ��     ��5� ���      ��                       ��5� ���      ? ?                      ��5� ���     �  �                     ��5� ���    �   �         �         ��5� ���   �     �       � �         ��5� ���  ��      ��     �  ?        ��5� ��� ��       �� 0  �   �  0    �p5Wp�e�         �   <     �       �p5Wp�U<            �           �p5Wp�V              �      � �     �p5Wp�X               �      �     �p5Wp�X                              �p5Wp�`      3                       �p5Wp�`     ��                      �\5W���                 �          �\5W���    � �          �         �\5W,�	    0            0 0         �\5W,�%       <          �        �\5W�Օ   �    �        �           �\5Wl�V   ?     ?       <   �        �\=_\�X  �     �                 �Wp5W�`5  �      �?     �            �� �5���5 �?       �     <     �       �7\7'\6 �       �  �            �_=<_=8 �        �?   �     �      ��_�<�_�8                  ��     ���0���0    �?         �      ?      ۳V�3�V�3    ��            �?         ��Z�3�Z�3    ��            \�        ��U�3�U�3    ��:            WU        ��j�3�j�3    ��:            WU5        ����0���9    ��?            \�5        ����<���9    ���           ��?        ��?<[�9    \���          ���       �7�7W�_5    \�ת>          \���      �� �5W�U5    ��U��         \�ת>      �Wp5W�Z5     �U��         ��U��     �\=_\�`     pի�:          �U��     �\5W���   � |ծ��          pի�:     �\5W,�    W�W����        � |ծ��     �\5W,�
  �WU���        W�W����     �\5W,�%   �U���      �WU���     �\5W�Օ   ��?  ��       �U���    �\5Wl�U   �� ���       ��?  ��    �p5Wp�U  ��  ��        �� ���    �p5Wp�V  � � �W�       ��  ��     �p5Wp�X  0 < pU�       � �  �     �p5Wp�X  0 ��_U�?       0 <  \�     �p5Wp�X  0 ��W���       0 ���W�?     �p5Wp�`  � W�<      0 ���U��     �p5Wp�`  ��? W_?� �    � �U�<    ��5� ���  � �� \�?�� <    ��? p�?� �  ��5� ���   ��\=  �  � �� \�<�� <  ��5� ��� �  0�p=�<     ��\=  � ��5� ��� 0  <0?��0�  0 �  0�\5�<   ��5� ��� 0  <0���0� 0 0  <0?p�0�  0 ��5� ���   ���   � 0  <0���0� 0 ��5� ���   ��o�  < �   ���   � � 77  �5  � ������    ���� < � � 77  �5  �  �< ���   � ?�����  � 77  �5  �  ������   �  <����  � 77  �5  0  ��?�<   �  W����  � 77  �5     �?     0  �= 3  � <  �    � 0��?   �        33   � <  �    �      �    � 0�3   � � <  � 0   0    0   0    �      � � 0  � 0   0    0   0 0   0    0   0 � 0  � �       �    0   0    0   0 � �   �    �      � �       �    ۪������ � <      � <    �      � ��_�W�ouu  �       �   � <      � <  ���	���9   �� ���      �       �  �d���P  �� �׫        �� ���    �Tdp6@  � � p��       ��  ��     ��l�9  0 < \��       � � ���     ��P�y��  0 ����?       0 < p}�     �+:o>�WW  0 ���_��       0 ���_�?     �UUUUUU    � �]�<      0 ���_��     ��?�    ��?  _5� �    � pW�<    �����   � ��  \=�� <    ��? �U=� �  ��0�    �� W  �  � �� �U?�� <  ���  �  0� W�<     ��p�  � ���  0  <0? W0�  0 �  0�p5�<   ��� �  0  <0� W0� 0 0  <0?\�0�  0 �?����    ��W  � 0  <0�\�0� 0 � � �    ��\ < �   ��W�   � �������   � /\333�    ��W�  < � �UUUUUU   �  �����   � _�����  ����?�   �  ������   �  �? ���  ������   0  ̪?�<   �  ������  ������      ���    0  ë�? 3  �0�?�     � 0W�   �     W 33   �����     �  �   �    � �13   � �����  0   0    0   0    �      � ��?�  0   0    0   0 0   0    0   0 � � �  �       �    0   0    0   0 �������    �      � �       �    �?        � <      � <    �      � �7         �       �   � <      � <  �?                        �       �  �  �������                �� ���    � �_UUuUUU�               ��  ��     � |�������U              � �  ��     � WjUUuUUUj5 UUUUUUUUU    0 < ��     ���U�����j�� ���?�?�    0 ���W�?     �pY�UUuUU�ZY� �������    0 ���U��     �p�V�����_�e� �� ����    � pU�<    �\f�������Wf�?��?���    ��? \�?� �  ۜe�������~��������   � �� W=<�� <  לY�������z���������    ��W  � �٪��������?�?�?�  �  0��U�<   ۜY�������z� � � �  0  <0���0�  0 לe�������~����������  0  <0���0� 0 �\f�������Wf   UUUUUU    ����   � �p�V�����_�e   ?���    ����  < � �pY�UUUUU�ZY   �����   � �U�333�  ���U�����j��    �����   �  o< ���  � WjUUUUUUj5    <����   �  ������  � |�������U    ����   0  ��?�<  � �_UUUUUU�     �����         �   �  �������     ?���     � 0��   � �                � �     �      � �               ������  0   0    0   0 �������������������?    0   0    0   0 �UUUUUUUUUUUUUUUUUU    �       �    �UU��_��W�W����_UU      �      � �UU�U}U_�W_�W�U}UUU     � <      � <  �UU}UUU_�U}�U}U_UUU      �       �  �UU��U}����WU_UUU                    �UUUU�U}�U}}U_�WUUU                     UUU_}U��W_}U_�WUUU                     UUU�_U��W__�W�UUUU                     UUUUUUUUUUUUUUUUUU                     ����������������������������������������                                      ��                                      ? �                                    �   �                                  �     � ������������������������������ �       �WUUUUUUUUUUUUUUUUUUUUUUUUUUUU��         \UUUUU���_�U�UU__��U}U}UUUUU5          \UUUUU�UUU�U__U__�U�U_U_UUUUU5         pUUUUU�WUU�W_�U__}UUU_U_UUUUU    ��   pUUUUU���U�W}�W__��W���WUUUUU   � �  �UUUUUU_UU�W}U___UU_�W�WUUUUU  �   � �UUUUUUUUU_�U�___�W�U�UUUUUU �     � WUUUUU}UUU_�UU__��U�U�UUUUU� �       ��WUUUUUUUUUUUUUUUUUUUUUUUUUU��          ���������������������������?      H���j�Ņkhdd �é  ۥd����i` k�xH����΅ hX� � ��*��+ ��H���&��'h�h� ��H���&��'h�`� ��H�˅&�ƅ'h�(�  � �ɢX ��d>d?��JdId8d7dBdGH�_�� �h�H�J����hH����h ��H�_�� �h�WH�J����hH�$���h ��H����h !� 뜩�H����h 7�H�$���h !ϩ�H�$���h 7� �� �� �͢,�x��*��+ �֢4��H�҅&�ƅ'h  �d5 wʰ)�4��H�څ&�ƅ'h  � wʰ�4��H��&�ƅ'h  Ԁ� ۢ<�x�� �� � ���dL�xH�#��΅ hX�P�"d#d$d%��]dXdYd5d!��;�h���; k� m�H�$���h !ϥ8��7�N�8���8�D�8�Cm � � m!�!�Ce>�>� e?�?�JeC�J���8��J�IeC�I���8��I 뜩�H����h 7���H�$���h 7��;m&�&� m'�' ���  I�ɀ� ʭ  I������i`�]�"�]�,�x��*��+ �֢4��H��&�ƅ'h ԥX�"�(��% @Ӣ8��$ �ӢP��#�JJe �ҥX�:�L6��XH��&�ƅ'h��Y�':�`�YH��&�ƅ'h�$�d�	�*��+ �֢,�l Ԁ3� 8�߭!��	 �۩�X��&8�߭'����Y�$�[�#�Z�%�\ �� ��L���Y�,H� ��P�h ��Fbfa�\�H�����hH�����h � �� ��`�X���C`�B��  I��0�@H����h !ϥF�>dB�:�  I��0�"H����h !ϥF� ��B�7������GI�G��7�:�7dC�7��C���
�C����C`�IiHH��  �עO� h �ע�� h �ש�/�Ji�ZZZ��  ��z�M�  ��z���  ��hi��/��`���������������������H�8�>���?�h�/��+��8���Z�i%�� ��zhi���Z ��hi(���L��`H�����hH����h���������J����H�8�>���?�h�����8�������� ��H����h�e�� e���`x  t ,_  �  w  �  � 3 � K � � ��  	  
    �Y�        �J�H���j�Ņkh �â � ��*��+ �� ��H�M�&���'h�(�  �H�˅&�ƅ'h�(�  �H���&��'h�h� ��H���&��'h�`� ��H�Q�&���'h���
H�V�&���'h�P�  �xH�#��΅ hXH���>��?hH�[����h� H����hH�����h ��H�m����h�H�$���hH�����h �Ωc�"d#d$d%dXdYdId^dC�x�c��7d8dGdA��5�
�6�hi�; k� 3�H����h !�H�$���h !� �� � �� � ��H����hH�$���h�"�(��H�$���hH����h �H����h � �� f��7i�@�8�&�8�7Je@�@H����hH�$���h�� Q��@H����hH�$���h �ڦ>�>�8�>�>�?d?�?�?��@eI� ��8� �I�7Ji��c8��c0�����c�7��:�7�P8�6JJJJec�c�x���x�c�;iH�$���hH����h ��(H����hH�$���h�� ���d���� Q�H� ��!�h�8�2��� �H����h �����8��8� @ӥX�"�(��% @Ӣ8��$ �ӢP��#�JJe �ҭ  I�ɀ� ʭ  I������i`�X�:�Lա�XH��&�ƅ'h��Y�':�`�YH��&�ƅ'h�$�0�	�*��+ �֢,�8 Ԁ3� 8��!��	 �۩�X��&8��'����Y�%�\�$�[�#�Z �� ��Lx��Y�=H� ��Z�h ��FbfaH�����hH�����h�����\��� Ȁ 0� �� ��`��e�� e����e�� e����8���� ��e�� e���������ڦ��8���d���H����h�8�2��� �H����h ��H����h�8���� ��e�� e���������8�2��� � ��H�8�����h�"������e���8�0���������H���h����` 0ݩ ` ֣�  I��H����hH�$���h�����ȱ���H�8�����h�)��1��9��)���	���6 ���1��� ģ�������ǰ� ������ ���
���
������:� �`�  I�����`�c����7���
�`�7:���7`��������������������� ���d�8���^�d �Ӆ�e��d8��H����h��3�8�2��� �H����h ��H����hdd�8����� ��
H����hddH����h�8�(�����
H����hH����hH�>��?�h�8�2��� � ��H����h�8�(�����H�e��e�hH����h�8����� ��H�e��e�hH�8�����h�.����I�E����Hi��Z�3 ��zhi 	����'i������ɠ��Zڥ3 ��hzi ɠ���3�`H�Z ��hi��hiL�ԥ^)�i�3� �^)�eI� ��8� � �̩(8���^JJJ�.�8�.�.�.�#0!��3�i� ��8� HZ ��hi�h�.��`�҅3�P8�^��IL�̩�-�H��0�d�-��^

�d �Ӆ�e��^J���8�e�� � ��h
�-�Ţ ���L�ԩ�l�� ��H�>��?�h�8�2��� �H����h ��H��� �h �Ӆ�O8��� 
����ik�ȹ��i���L��H�>��?�h�8�2��� �H����h ��H������h������������4�H�8�����h�����ϲ�C�dG����G�	�"�8��G�^eC� �����^`\]1 $%0: $%1: '  +  /  3  7  �[�;  ?  C  G  K  �m��X�X�XXX��� ��  L��� >��
		
	
 !"#$%&'(())
)	(('&%$#"! ����������������������������������������������������������������?<<<300030003000                           ?<<<300030003000                           ?<<<300030003000                                                                                                           																















    				



    !!!!""""####$$$$%%%%&&&&''''(((())))****++++,,,,----....////0000111122223333444455556666777788889999::::;;;;<<<<====>>>>????  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|��������������������������������  $(,048<@DHLPTX\`dhlptx|����������������������������������������i����!� 	� \ 'q 2!"4VDEh��h�ۻ��������������������������쇾�Ez�Fu  Q                            #42#VeVf��w����˽���������������˪��ۘ�������������������������������������������������������������̻��������˻�̻�����������ffvUDC332                          "#324D3DUUUVfgffwwgxwwwx�ww�ww��wwwwwwwwvgwfgvffffgvgwwwwwwx����������������������������˻�������������wwffeUUTDD3333""""""""""""#333DDDDUUVffwwwx���������������������������������������������������������������˻�������������������wwwwwvfffffffUUUUUUUUUUUUUUTEUUTDDDDDDDDDDDDDDDDDEUUUUUUUUUUUUUUUUUUUUUUUUUeVfffffffffffffffffffgwwwwwwwwwwwwwx��������������������������������������������������������������������������������������������������������wwwwwwwwwwwwwwwwwwwwwwwwwwwwwwww�������������������������������������������������������������������������������������������������������������g�@�KV�������o���  �   `    ���(���������������@�0���P���������             �PJm�~���������������������ٶ�
p\_��I�P                       ?o�������������������o�u� b        # @(� @          8��������������������������W�B�a       ��<P�R����)"�?��Tf����������������������&�@              $ %Sl������̞��)�50F��X��������������������o�d��Q                @�n��������������������{猃z��4sWRfGA aEf����W�h���v�6Tc�8TFr$&eVTVGC�k���������������������eW2 0            E8GU>���������������z��G��X6=U4q6G�S�xF������G��5K�1b Q3B#5F�$�3xuh�W�EGu�������ܬ��������������ʗ�cU       4!��e�����x���ݚ���������}ּ��ic{e~�3f�uId�X�x�y{v~ۅz�gxw�y����W���ggGde#Ev%dGSTFggtifkhf����������������ۻ���8CfT3$1tTSTGBx%TJe�eewsw�V�xdytxY��������������������tFC3   10SWf����̻�쬺�ʌ����ewFg4r$"%2V2eGdh��z����̽�������ܺ����wVvT%TDER2D32UcU6cxww��y��������w�j��g�w��v������̬����������˪�v�44#       !DdXx�������������껩�v�WwfvdvFvVwgwy��y�j���xvvFwDfWuwV�v�x������̫�˻����G�WeT5DVDFefV�v�����۫�ܼ�ܺ�����xwvfVfwgewffwhvw�f�wx������g�wvh�x���������v�wehdVVeF�Wxv�y��˹���������ۛ��efD3       35Txx��������������ʺ���eeEcED5ETFvfvy����������xx�fuWUeUFfWfWww�y������ܽ��̺������gugeUFeFTTFffxw�x�����˼˻�����wuUUDD3B"""4CUUvx��������������̺���xeUUDB4"31#3DDTVUWvVwvgx��������������˻������x�wudUTDTDDUEfwhh�x���������������xxwgwgfgWgww���������������������������x�x��wfwfUVTTETEDUVffy���������̻�̻�����wvuVdUDDUUCUVVgx��������������y�wvwufefVeffgww�������������������wwfvgfffVfvfVfvww�wx���������������wvwwgwvwwwwxw�w�����������whvfEVUVeeVfwww���������˼������ufUTCDC3DDDDVff����������̻��������wffTeVEEUUUffw�����������������wwvffVeUeUUVUWgxx�����������������wvfeEDUDDDTUEUfvwx������̼�̼�����wfeTD332"#333DEffx�������������̻�����fUTD4333C4DEUVfgw�����������������wwwwvfffffgwww����������������wwwfffUUUUUUVVfffwx�����������������������wwfffffffffffffgwwwx����������������������w��Uy���1 $h�����ʆS   5i�����S!#Ex���˻���fffwx���������wfwww��x�������ww��wx�������w�������wwwwx���������������x�x��������w��w����������x������������w�������ww������������x�����������ww�������������wwww��������x����������x��������������������wwwx��������������������������������������������������������� rw�r��љv� �8+j�UUա�O  ��둙����O���H�'��af��r���w'""��"�""rw�www""'"""""""ww""w'""""""rw""r""""wwww'""""""""""""""r'"'""""""""w"rw""""""""""'"""""r""""""w"""""""ww""""""""""""'""""""""""rww"""r"""""""""wwww"""""""r'""""""""""'""""""""""rr""""""""www'""""""""""""""""""""""""""""""""""""""""""""""""""""""""" ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������xآ����
 �� ղ �d� �۩�
 ��H�I����hH� ���h�� ��������������
 �� �X��
 �͢�~��������������B����G�����r��������l� �g��fd
 ��xH����΅ hX���A��6 �ͩ �dI���0dK���J�� ��*��+ ��d1d8��7dCdG�����H�/���h���Ƒ����e�� e����d5H�����h �͉�
H�-���h�jH����hdd ��H� �>� �?h k� �ũ��0�" �ץ0����� �0���3�I�0 �� :˥I:)�I �˥J8��Jɠ��ɸ�����J�K��K��dKH����h !�H����h 	Х5��1��:��E�@�A��Oɀ�Li�d5 �� ^� �̭ ����LJ�L��1��8��1�8�٥1�!��i�1�8�ʥ8�=���� ��L���8�8�����LXǩ�l�f�������l�f:���f���g���� ��g:��gL���  �dh�f���f�l� �� ǥgH���ǅh��HH�&��ǅh��:H�0��ǅh��,H�:��ǅh��H�D��ǅh��H�N��ǅh��� F�L��dh�l� �� �H���ǅh F�H�&��ǅh F�H�0��ǅh F�H�:��ǅh F�H�D��ǅh F�H�N��ǅh Fåh�h�ЦL����e�f��H�ZH����h�e:e�� e���>dadbdi �� �ͩ�
 �� � q��i��H����h�e:e�� e��� t��ez���h:Г`l  �͢� ��*��+ �֢��� �ע,�2��*��+ �֢D�> �ɢ�> �ɢ��> �ɢ�d��*��+ ��H�j�&�k�'h�&��&��'�p  ԥf������� �׭  I����ɀ���Z �ͭ  I�������L�ͺ�蚩�i`��&��*��+ �֥gH�l�&�Ņ'h�PH�w�&�Ņ'h��BH���&�Ņ'h��4H���&�Ņ'h��&H���&�Ņ'h��H���&�Ņ'h��
H���&�Ņ'h�&�&��'��2 ԥfH���&�Ņ'h��4H���&�Ņ'h��&H�ą&�Ņ'h��H�υ&�Ņ'h��
H�څ&�Ņ'h�&�&��'��= Ԣ4�HH��&�Ņ'h Ԣ0�SH��&�Ņ'h ԩ�H�$�1i2��> 
עt�1i2��< 
�`,FULL GAME 4HURDLES ,LONG JUMP 4ARCHERY 0SHOT PUT 8ROWING 4CYCLING 01 PLAYER ,2 PLAYERS ,3 PLAYERS ,4 PLAYERS 4LINK-UP SIGN-ON HI-SCORE �C��C`H��� �h�G�
H����h�7� �� �7���T�H��Ch�'d���e�� e��� �ץ7���C�GI�G`��8����7d�H�e��e�h ��`d�H�e��e�h�� �ץ78���8����7d���e�� e� ��`00000 ;=& UP 00.00 0:00.0  READY  GET SET   GO!   YOU WON! YOU LOST! �  ۩�
 �ͩ�e�f� 4��e����dl`� �
 ��L �� �
 ��L๩�
 ��L ���
 ��L����
 ��L ���
 ��Lh��  ۩�
 �� �� �� �� ��L��HIGH SCORES ��
 ��H�>����h�h�&H�K����h��H�X����h��
H�e����h�������`�������H�8�_��`h����i�������H�8�_��`h���`�H���h��_��K`�����[��
���Z����i�\�J�����[��
�:��Z�4�2�Z�H���h��[��<���+��* ��H���&�ȅ'h�H�L �`WORLD RECORD! d�\��<��[e��Z�H�8�����h�
H��a��bh`H�&��'�hH�,�&�Ʌ'h��H�&��'�hH�*�&�Ʌ'h��ZH  �h�zhe������Z ��zhi��.�Z 
�zhi�����L��# $% ��x��*��+ �֢��H���&�ƅ'h Ԣ ���@ 
� �� �̥A�dA�^�Z��^�^����^ �� �� ��L^�`dH�d���	�ک+ 
����+ 
�`���eZ�Z� @�hi�zH�&�ƅ'h  � ���hi�L �H��&��'h�e:

e&�&� e'�'` �ɲi�L�� �ɲi�L�ץeH����h:e�� e�`H��� �hxH�܅�΅ hX��`��*��+ �֢�l��H�p�&�ʅ'h �ע8��  Ԣ
 ������  I�ɀ��xH���� hX`PAUSED �d �ͥ5���
��蚩�i`�5)0����`8`�6����%������#����-����7��	��F��� �7`�9�9�
�d9 ���2����=��;�h��;``����� �Ԣ���c�!����� �Ԣ>�������` �Ԣ>���P8�6JJJ��.�Z�� ��zhi��.��`���p��-� HZ� ����i�zh�-��`� �Zک��$ ����i �z���`� �Zک��L ����i �z���`���p�
�-� HZ� ����i�zh�-��`�i�d� L�שj�p� L�צJ�KH�ʅ���h� �&H�ԅ���h��H�م���h��
H�ą���h�z��������������� ��hi���`�`�Ji����-�KH�ZH�@���he�� e�� ��z��i����8���h�
��� �-��`�C�� �̀�C� z̥I8�)�I`d�7�!�8�7��J8�)�J(��K�
��� �K`���3� �I �̠@�Ii)xi����-�Z�3 ��z��i ����8����-��X`H�����hH� ��F�h��.H� ���hH� ��F�h��H� ���hH� ��O�h�x� ����������X`x�H����h� �������H����h�0e�� e�����X`H� ���h���0H����h� �������H����h�0e�� e����`�d �����`����`�





	�& `ڢ�)Hi8

&&&�����`� � �@�� �� ��������`H�Z�' J� έ$ �	J��%  �z�h@���# `d�`l xH�!�#�"���$� �#�$�<���%� �$�  )����A�5��� ���������+�  )0I0�� �5��  )0I0� ��5�6���8��6��6�P���O�6�6�$ ����# Z��y ?�斥�� ��zhX@xH�!�  I���A��6��5�A��6�dA��xH�$ ����# hX@�������������������������� �`� �F������������������������������H���h���@I�ڦ��8���d����e�� e��������e�H���h���H���h���H���h�����"��F����������H����h��H���h���`����������������H�8�>���?�h�����&�����i��
���ɠ��������L��`dG�������H�8�����h���
�����G`H�L��M�h�iH�P�� �h %�H��L��MhH�N��O�h�iH�Q�� �h %�H��N��Oh`H�R��S�h�yH�V�� �h %�H��R��ShH�T��U�h�yH�W�� �h %�H��T��Uh`������H���h��H�8�>���?�h�2���������i���'������������� �`���ɠ��k���i��� ��`H�����h�.H������h�"H�����h�H�H����h�
H�j����hH����h���������^����H�8�>���?�h�����&�����i��
���ɠ�������� ��H����h�e�� e���`��H� ���hH����h �� ��H�d�� �h �� �ө.����H�
�� �h �� �ӥ �ө �H� �&��'hL �dd�H� ���hH�d�� �h �ө�H�
�� �h �� �ө �H� �&��'hL �d�dH� ���hH�d�� �h �� ��H�
�� �h �� �ө�� �ө �H� �&��'hLԩ��d�dH� ���hH�d�� �h �� ��H�
�� �h �� �ө�� �ө �H� �&��'hL �d�dH� ���hH�d�� �h �� �ө�H�
�� �h �� �ӥ �ө �H� �&��'h�M� �����i0������`� H����hH�8�����h���H����h`��H�dH�&�&��'� ��Z 
�zhi���`����d�&&&&��&e��e��JJe�� e��)�`d�&&&��&&e��e��JJe�� e�`������i������`d� ����������L�֘8� �� � <ԩ e���e��d�&&e�� e��Ke���e�����H� ����h��H� ����h��
H�J���h���������8������iJJ�*����eL�օ+e8���	��+8��+�� }�H�e��e�h�+�L��ɠ��L�֥*�,H����hH����hd)��(��H��4���(�)� �� �� �(�)� �)�&�(�)� �� �(�)� �)��(�)� �(�)� �)�(� 2(�����)� 2)�����,�L��H����h�(e�� e�H����h�0e�� e��+�L��`��H�dH�+�-�*�.�� �֘i��� �֘i��-���ZH�.�/hH �֊i�hiH �֊i�h�/��i ��z�`�ZH <ԥH)�� e���e��� e��@e�h ��z�`d��e��e� <ԥH)�� e���e��� e��@e�d4L��d��e��e� <ԥH)�� e���e��� e��@e����4�TH <ԩ e��@e�h�: <ԩ e��@e�d4�,���	�H�i��h����`H <ԩ e���e�hd4d�H����h&&H�e��e�h�Ke���e�����H� ����h��H� ����h��
H�J���h��������������iJJ�*�����+�� }�H�e��e�h�*�,H����hH����hd)�E4�(��Z��4���(�)� �� �� �(�)� �)�&�(�)� �� �(�)� �)��(�)� �(�)� �)�(�����)��
�(��������,�L��H����h�(e�� e�H����h�0e�� e��+�Lt�`���`�چz�
�{�5�%��A�{�|}�9�{i�� Y��.�z�5�%��%�{�����z��0�{�|+�|��})�ڠ> �ۀҀg)�����
I

��@�  �ڀOH�z��	���hu�����I

�ڹ>ܝ ��ܝ �{i|� f�ڦz��)� ڊ�{�����	@�� �z�� 	@� ��0LF�`H� �n fۡ �m f�hem�m��n)�uFnfmFnfmFnfm�z��)�u���n�m`R�R�S���cڋڤ���۽�`�z
i|�� �z�� Lfۦz�5�I�%���t�� � ���� ���� ���( `��)����t��� �ۜ �( d�`�{i|�ڦz��)� ڊ�{����`�{�|�|��}�z�� `�{i|�� H fۡ � fۡ  f۪���h`hL�ۥ�8�


e{��{��ܙ| ��ܙ} �zt�`���u��� �ۜ �( �* �u�L��


�� ��ܙ| ���������t�����t�t���d�d��u��`� � ����`� ��`
�m��em�m�i �n��m��m��m�n` m�lm H�Z� �n�mm	 � ��m� ȱm� ȱm� ��� z�h`dy�y��`x �۩��X` �ۜ � � � `� � � � `��* ��* ���( ���) d����`���`��d��( `��JJJJ��yJJJJ)} ����	��( ` @��v
�F�F��o/�R"�ʢ|X7�����zdP=+����Ǽ������}voic]XSNJFB>:741.+)&$"                                       Ֆ���  ��    *�z�ʴ  &�N�v�  ��  ��  /�-�    0I��I�I����� P ( � (�		 ��ݠL�ۢݠ	�L�۩�ݠL��� ����� �  ( (( (((T 4T5T5T5  4 4 4 4 �� �K
 �� X
X
<|
H|
0r
<r
 b
b
Hr
�H o. l P  Q  R  S  T  U  V  W  % @%
\o |o % @%
\S |S % @%
 R @R % @%
\7 |7 % @%
 6 @6\& |&
\o |o\& |&
\S |S\& |&
 R @R\& |&
\7 |7\& |&
 6 @6 (  )8(| $( )44) F( E)8F(|E$( n4T)T 4n$�n t) pnTcXmTE * (*,/L/</`/ d�< @�0t&TM �4hc \ h 22      @  @  @  `  � � \ D L T LDLTLTu+ v*v*,v*@v*D*cdu<d�<                 (     0 H ` H       0  `  � �   @ @  @ 0@ @@ P@ `@ p@ 0 (  �0  P H� 0� �@ @ �h $ tP0 ��   `�      X  `  h  p  x  �  �  X ` h p x � x �  � � � (� 8� H� P Q R S T U  pp X�   Xp  Yp  Zp  [p  \p  ]p  ^p
  _p	  `p  ap  bp  cp  dp  ep  fp  gp  Xp  Xp  Xp  Xp  Xp  Xp  Xp  Xp  Xp	  Xp
  Xp  Xp  Xp  Xp  Xp  hp  hp  hp  hp  hp  hp  hp  hp  hp	  hp
  hp  hp  hp  hp  hp  hp  ip  jp  kp  lp  mp  np
  op	  pp  qp  rp  sp  tp  up  vp  wp  xp  xp  xp  xp  xp  xp  xp  xp  xp	  xp
  xp  xp  xp  xp  xp  xp  yp  zp  {p  |p  }p  ~p
  p	  �p  �p  �p  �p  �p  �p  �p  �p  x� P8 0P 8P @P XP X8 `8 h8 p� hP 88 (P 08 P � p8 x8 �8 �8 �8 �8 �  �  � ( HP  P PP � @8 `P  0 0 0 0  0 (0 00 80 @0 H0 P0 X0 `0 h0 p0 x0 �0 �0 �0 �0  8 8 8 8  8 (8 H8 � �c P�O P ���Q P �w�R�S�S�S TP��w�R	�S�TP ��w�Q	 TT P ��w�e �f  f  e  e  f  f  e  e  f  f  e �e �e �e e e ���P  �w�R����S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S�S S S S S S S �[�[[[[[[[[�p�[  e�e  �v�P
 Q  P O� ���  �  � � �  ��� �  ���d V�U V ���W V ���X�Y�Y�Y ZV����X	�Y�ZV ����W	 ZZ V ����g �h  h  g  g  h  h  g  g  h  h  g �g �g �g g g ���V
 W  V U� �-������������ƪ������%UU�������������������������    ZUUUU����������������?UUUUUUUUUUUUUU�?�nUUUU��QUU��UUUUUUUU�}w__�]�u��u} <<<�������TUU��_UUUUUUUU�WwwWw�����uw]W <<���������������__�W���]w___�]����u]]�����������������_�W���uwWWw�]���uw]u� <<�������������W}}_�W���_Wwu��u��u]_� <<��������������_�W���UUUUUUUUUUUUUU� ��e  ������  ��_�W���������������      �e  ���UU�  �W}}_�W�U�UUUUUUUUUUUU����e  ���UU�  �W}}������}��}���]��}u�	<<<<�e  ��zUU���W}}����������]��]�]�ݫ&<<<?�e  ��zUU��_UUUUUUUU�����}��_u}}ݫ��?�?�e  ��zUU�  UUUUUUUU�����]�]W]]���: <�<�e  ��^UU�����������?}]�}��WW���u� <<�e  ��^UU�����������UUUUUUUUUUUU�������������������������������������      �J���ww���ꫪ���ꫪ  Uի�����UUUU  ���S�J�
���]UUի����ꫪ  Uի�����UUUU0VUU	J�P�ww���ꫪ���ꫪ  Uի�����UUUU�ZUU%�PH!���]UUի����ꫪ  Uի�����UUUU������
AA��ww����WUUUUի�  U�    �UUUU�fUU� @ ���]UU�WUUUUի�  U�    �UUUU��f}��WUUUU�ww����WUUUUի�  U�    �UUUU  f}��WUUUU�WUUUU�WUUUUի�  U�    �UUUU  f}ߗ @ �������WUUUUի�  U�    �UUUU  f}ߗ�
AA��WUUUU�WUUUUի�  U�WUUUU�UUUU< f}ߗ�PH!ꫪ���ꫪ���ꫪ  U�WUUUU�UUUU� f}ߗJ�P�WUUUUի����ꫪ  U�WUUUUժ���<f}��S�J�
ū����ꫪ���ꫪ  U�WUUUUժ��� f}���J���WUUUUի����ꫪ  U�WUUUU�ZUUUlUU�������������������������������iUUU  �����������������������������������UUU      ������    ���  ��������    ��VUU  ���������    ���  ����������   �UZUU  VUU	������    ���  ��������3�� �UiUU  ZUU%    � � ���  ����������*��U�UU  ���� �  � �
 ���  ��������3����U�VU  fUU� �
 � �* ���  �ꫪ����3���UUZU  f�� � � �* ���  �ꫪ������� �UUiU  ���� �
 � �* ���  �ꫪ������ �UU�U  ��}� �  � �
 ���  �ꫪ���� �>�UU�V  f�}�    � � ���  �ꫪ���� ��<�      f}}�    �    ���  ��WUUUU� ����      f_}�������    ���  ��WUUUU� ���      ����������    ���  ��WUUUU�  <�      ����������    ���  ��WUUUU�    �      lUU�������������������������������      ����                                        �����?�?�<<� <<<< <<<������?<<<<<<<<< < <<<<� <<< ??�<<<<<<<<<<<�<<<<< <<< < < <<� <�< �?�?<<<<<<<<< ��?�< <<��<?�?� <� < �<�?<<�<<���<<<<< <<< < <<<<� <�< <<?<<< �?<< <�<<<<<<<<< < <<<<�<<<< <<<<<< <<<<<�<<����?< �<<��<<�?<<<�< �<<<��                                        <<<<<<<<<�?    �<<� � ���? �?�<<<<<<<<< <    <<�?<����<< �< < <<<<<�<<      <�?0 ��� <���< <<<<�<���     �� ���  < <�<<<<�?���     ��    ���� <�? <<<<<�??<<�< ��   �     ���� << <<<<��<<<��?�< �       � ��?� ��                                   @   ������������������������  PT�
  VUU	VUU	VUU	VUU	VUU	VUU	VUU	VUU	  U��  ZUU%ZUU%ZUU%ZUU%ZUU%ZUU%ZUU%ZUU% @EUU� �������������������������������� PEUU�
 fUU�fUU�fUU�fUU�fUU�fUU�fUU�fUU�UUUUUUUU����W������f�������f��f����ן������������������������������������������������f�}���}��W}��W}�f�}���}���}��}�����J���Jf}���}��}��}�f�}�f}���}��}���UUI�UUIf}���}���}���}�f}}���}�f�}��}��nUU�nUU�f�}�f�}�f�}���}�f}}���}�f�}��}��n�Wen�We����f�����������f_��������������nuYenuYe���f������f��f_��f�������ןn`en`elUU�lUU�lUU�lUU�lUU�lUU�lUU�lUU�n`en`e��������������������������������n�en�e� 0�                      0����n�en�e� <�   �              � ����n�en�e� �   �  33�0??0����n�en�e���
   �U  33333�� � ����n�en�e�� �
   ���?333?�3�<� 0����n�en�e�< �*   ��  ?3?333�0  ����n�en�e�      �  33<?3?3??  0����n�en�e�      �                  ������������                            ����UUUUUUUU  ����?��?�� �����?�� � �������j���� � <����0 � � �� <�  ����nnnf~�n� pUu�\WWWU�U� �U�U�uUupU5 ����[[Zj~�[� 0�0� ���� ����0000�0 �������i�}�i p�u�\WU�\�5�  \�5�u�up? ����fffn^�f� 0�0 ��0   ���0�0�0  �������j�i�� 0�0   �0   � �0 0 �  ����nnnf~�n� �κ�������:   �Ϊ���� � �������i�i�e �κ����?�:   ������ � �������i�k�e p�up5�\� �5�  \�5�u�u	��5 ����������� �����:�� ���  ��:�κ���: UUUUUUUUUUUU pUuUu5�\� �U�  \�5�u�uUuU5 UUUU�������j �����:�� �:  ��:�κ��� UUUU~�����nf  ����?��� ��  ��?�����?� ����~��[j                            �����}ff�f�i                            UUUU^�����fn                            UUUU�if�f��j <3<? ���0����   � 0 ����~�����nf 333����<3 �0�  ? 0 � UUUU�iffvf�i ?33������ �0� ��03��UUUU�k���i 3330�� ����0�  �0 � ���������� <3? � �0� 0�0�   � 0 UUUUUU}�~UU                            UUUUU�  �WU                            ����U}  �~U               0           UUUU�    �     <<��� �����3��0�0   UUUU^    ��     �� 0�03�  �0303   UUUU�������     <<<00 �����  ��0��    ����~��fzg��     ���  �03�  �000�    UUUUmwfݙ�]v     ��<< ��03�  0�3�    UUUU�fj�����                            UUUU ��fzg�                             ������������                            UUUUUUU�UUU� <��� <� 33?������ UUUU  �  � 33333��30�� 3333�� 303UUUU�������� 3?��0<� 3333�����0UUUU�������� 33333�30�0 3333�0003����UUUUUUUU 333��� <0 �0?���3� ������������                            ����UUUUUUUU                            �   ��������                            p�              ������� �0?<     �	���������     �������0 ���03     �&�UUUUUUUU     �������0 �0     �>�UUUUUUUU     ��� ����0 030     ��UUUUUUUU      � ����0 ����0     �  U�_��UU�                            ��_�wuUW��                  ��00?������ W5pf�U003����������0 Ws���5WUUUU� e`Ypf00��00�00�0�03 �������UUUUUU?TPY�Y003�0��?�0�0��3 W����5|UUUUUU9?�@U �U033�0 � 0�0�03 �������_UUUUU��  ��<3��� ������0�7ps���|UUUUUU9��<�� �                  ��?3�jUUUU��>�<;�                        W������ �����5������������������������  ������ ���W{ժ�_UUUU�UUUUUUUUUUUUUUUU     ��  ����{���{UUUU�UUUUUUUUUUUUUUUU     ��  ����_W��+    �                          ���W���+    � �    � �              f���﷖+    � 0033?� ���            V��U�e�V+    � 00333� 303           Z��e�W�Z+    � 00333�����0           U��U�[�Z+    � 00333003 ��������  ����j+    � 00333003 RUUUUUU�  ���ګ���+    � 00�0?�3�        �  ���ׯ �+    � �    � �          �  �拏�ʨ�+    �                      �  �U���������ު���������������      �  �U����ꯪ����������������������������  �u����������������������������������  ��U����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � ���