                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                PUUU�UeUYY�ePUUUUUeUPVUU�UUePUUUUUYUPdeVA���eY�UPYY�e�UVP�e�YY�UPUf�e�YVPUeYAVYU�UYYPU�Ue�eUPVUUUUUUPVUYUUU�              "                                                                 UUAUU             @TUUUAU        eUUUPUYeAVV             @TU�UAZ        eYUYPU�UAUU             @��UVA�        U�eUPf�UAeY             @TUUeAV        YUUUPUYeAUU             @��eVAY        ��Ue�UUf�fY             @TYUUAe        Ue�UPY�UAUU             @&��YZAV        YUYUPUe�AiV             @TUUUAU        UUUU�U                                                                                UUUUBVUUd�eUAUUUUUUUAUVUTUUUPUUUUUUUYe�YA���TVUVAVVV�ee�AYef��VePV��YeUU�U�eAfeUdY�eA��ee��YAe�UdeYZPeefUVUfUeUUAUUeTUUUAYVUUUUUAUUUTUUUPUUUeUYUU���������������������������������������W�                                    _�_�                                    _�W�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�_�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    �W�                                    _�_�                                    _�W�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    �W�                                    _�_�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    _�W�                                    _�W�                                    �W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�W�                                    _�_�                                    �W�                                    _�W�                                    _�W�                                    _�W�������                        ������_�W}UUUUU�                        _UUUUU}�W_UUUUU�                        _UUUUU���     �                        ?     ����������                        �������߿�������                        󪪪����_UUUUUU�                        �UUUUUU�WUUUUU��                        �WUUUUUժ�������                        �������UUUUUU��                        #WUUUUUU      ��                        #      UUUUUU5�                        �\UUUUUUUUUUUU=�                        �|UUUUUUUUUUUU�                        �pUUUUUUUUUUUU��                        �rUUUUUU                                                                                                                                                                                                          �
  ���
�
�
����      8     888        �     ���  >>      �     ���  >>      �   �������>>      �   �������?>      �   �������?>      �   � ���  >      �   �� ���* >      �    ��� � >      �    ��� �>      �   ������>      �   ������>      �   ������>      �   � �
��  >      ��* ��
(������
      �   8� ��    8      �#  ����  >  �      �#  � 
�?  >  �    ���꣪�� �����>����    �������� �����?����    ������� �� ���?����                                                                                                                                                                          ����� *������
���
��* 
 
�� �#��8 �#8 �  8�� �#��8 �#8 �*�*8�⨊����( �#8���/��8
�������� �#8����8(� �����"�#8 ���8�� ���� *�#8 �  �8��� ����(�#8�
�  �8�� ����( �#8 8�  �8�
� ����� �#8�:�  �8�+� ������#8�?�  �8��� �����
�#8 ���8��� ����8+�#8 � �*8��� ����8,�*8�*�* 8�� � ��8  8 � 
 :�� � ��8 
 : પ��>�� ����:���>��������� ���?������       ��                           ��                    ���  ��?                    ��� ���� ��  �            ����? ������ �?     ����?  ����? ������ �?     �����  ����? ��������?     ����� ���� ��������? ��? ����� ���� ��������? ��� ����� ���   ����������������� ��?   ������>������?�����  ��   ������>������>����?  ��   ����  ��������>  �?   ��   ����  ���� ����>  �?   ��   ���?  ���� ���  �?   ��   ����  ���? ���  �?   ��   ���� ��� ��    �?   ��   ����? ��� ��    �?   ��   ����� ��� ���    �?   ��?   �����  �� ���   �?   ���   �����  �� ����   �?   ���� �����  ��  ���  �?   ���� �����  ��  ���  �?   ����? �� ��  ��   ��?  �?   ����? �� ��  ��   ��?  �?   ����? �? ��  �� ���?  �?    ���        �� �
��?  �?    ���        ��  ����?  �?                �?  ����?  �                    ����  �                    ����                        ����                          ��                                                                                                                                  �?                          ���                         ���?                         ����           ��  ���    ����� ���      �� ����    ����� ��� ��  �� ����    ����� ��� �� ��?  ���    ��������? �� ��?  ���    ��������� ��? ��?  ��3    ���������� ��? ��?  ��    ������ꃪ���? ��?          ������� ����? ��?          ����� �� ����? ��?          ����? �� ����? ��?          ����? �� ����? ��?          ����� �� ����? ��?          ������ꃪ���? ��?          ��?���������? ��?          �����������? ��?          �����������? ��?          �����������? ��?          ��?���������? ��?          ������������? ����         ���� �������? ����?         ��� ������������?         ��� ������������?              �� �����ꫪ��?              �� ����������              �� ����������              �> �� ����                        ����        ����> 8��8��8��8��8��8��8��8��8��8��8��8 8��>��   �� �� �� �� �� ��0�� �� �� �� �� �� �� ����, ��������> :�*8��8?�8 �8�+8�8�?��? �?��;�:+ 8��>������> 8��8��8 �8�8��80 8��8�8 �8��8��8 8��>��    |  �  � �5 �5 p p�\s\s�p�=WU5�= p p p p �����: 8��:��� ����: 8��8��8 �8��8��8��8 8��:������> 8��:��� � ����> :��8��8��8��8��8+ :��>�������� ������� � �� �0 �8 , ,  ��������� � ��_U=��5' 6' 6' 6' 6��5\U����5' 6' 6' 6' 6��5_U=���� <��0# 2# 2# 2# 2��2 2��2 �2 �2 �2��2��2��<< ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �
�.8�<�<��*�
�������+�*�*��(����/�
�������� .�/��(����* *�<�<8<���� < (�*�*�*�� �(𸺠*�*�*� �*��<𸰠*����(� .�����
�*<0�*������*�*��<���� �.�
��?��<�����<�<��?��<�����<����?�?����< < �����?��?<�<�<�<��?�����< �?�?< ��������< �?�?< < < ��� <�<������?<�<�<�����<�<�<��?�?�����?�?�?�?   <��<�<��?��<?<�<�< < < < < < �?�?<�����������<�<�<���������<�<�<��?��<�<�<�<����?�?��<�<����?< < �?��<�<�<�<��?���?��<�<��?�<<<���?<�?������?�?�?������<�<�<�<�<�<����?<�<�<�<�<����?�<�<�<�|�|�|��?�<�<��<���<<�<�<<<<<<�?�������� ��?������                  ���:�:�:��      ���    ����? � ?����� �  �������?����� �  �������?����� �  �����?�� � �  �����??�� � �  ���� ??�� � �  ���� ??����� �  ����� ??����� �  ����� ??����� �  ���?��??�� � �  �����??�� � �  ��?��?��� � �  ��?� ?��� � �  ��?� ?����������?���� ?�?��������?���� ? ��������?                   ���?�����?  ���������?  ��?�������?  ???����    ???����    ????���    ????����  ????����  ????����  ???����    ???����    ???����  ��????���  ��????����?��????����?��????����?��                                                          UUU�)��	�	�����	�	�)����������UUU�!""����������!""���������UUUթ���������������������������UUU�UUU�UUU�UUU�UUU�UUU���������UUU�  �  �  �  �  ���������UUUթ*�����)  �����*����������UUUՁ"��
*𡨢��
*��"���������UUU�  ��*��
(��*��  ���������  ��*�������UUUթ���)(������� �������������UUUUU�iUUUU�i�����i�����iUUUU镪����������      UUUUUUU�U�������i�������i�������iUUUUUU镪��������������             @   P  T  UU @UUPUUT�WT�_U�UU�~UU�UU�_UT�WPUU T      @   P  T  UU @UUPUUT�UT�ZU�UUU�UUU�YUU�ZUTUUPUU T      @   P  T  UU @UUPeUT�ZTiiUieUUiiUU�ZUUiUUTiUPUU T      @   P  T  UU @UUP�VT�VT�VU�VUU�VUUUUUU�VUT�VPUU T      @   P  T  UU @UUPUUTUUTeeUi�UUj�VUi�UUeeUTUUPUU T      @   P  T  UU @UUPUUTUUTVUUZ�VUj�VUZ�VUVUVTUUPUU T      @   P  T  UU @UUPYeTUUT�VU��UU�VUUUUUUYeUTUUPUU T   ��?�������?���?���������?�_W             W _P� � � � � � � � � � � � � � �P�W�������                        ������_�W}UUUUU�                        _UUUUU}�W_UUUUU�                        _UUUUU���     �                        ?     ����������                        �������߿�������                        󪪪����_UUUUUU�                        �UUUUUU�WUUUUU��                        �WUUUUUժ�������                        �������UUUUUU��                        #WUUUUUU      ��                        #      UUUUUU5�                        �\UUUUUUUUUUUU=�                        �|UUUUUUUUUUUU�                        �pUUUUUUUUUUUU��                        �rUUUUUUW���                                ��_�W}U�                                _U}�W_U�                                _U��� �                                ? ������                                ���߿���                                ��_UU�                                �UU�WU��                                �WUժ���                                ���UU��                                #WUU  ��                                #  UU5�                                �\UUUU=�                                �|UUUU�                                �pUUUU��                                �rUU �
  �*  �# ��� ���� *P
(U(hU(`U��`U��`U���U�  �*  
< ��  �*  ��  Ȏ  �����
� ��@�(PU((TU)�VU	�VU	�ZU	 ZU ��  <�  ?� ��  �� �:
 ��
 ��:��*��8��@	�?T	�BU�RU V�  V�  �
 @< P� ��  �� �:
 ��
 ��:�������8��.	��C	��P�>T 
�  J�  �
 � �P �*  ��  �� �����j��V���������*���
���
������ ��  �� @�@� �*  ��  �� �����j
�V�*���*������������������� ��  �j �P�@ � ��
 ��
 ��* ��* ���,��*`��*`��
���� V�  Z�  ��  �@� � ��
 ��
 ��* ��* ���,��*`�*`�
�U��U� V�  Z�  �j  <P�@�   �  �? �  ��������

�

��� �� �2 3�0 �?0 �0      �� ���  �0 ��� 0

0

������0

0
� ��0 �� �� �  �    �/  �0  0���0�0(3|,(����2+(8+(� ��2 ��2 �i? �� ? �          �/  �0  0���0�0(3|,(����2+(8+(� ��2 ��2 �i? <�  <  �  � �� �� ��0 0
� 0

������0

0

���  �0 ��� ��        �0 �?0 3�0 �2 ������

�

������ � �  �?� �   �    3  �=�(00(80���0����,(� /(� ��� ��� �i� ��� �        �    3  �=�(00(80���0����,(� /(� ��� ��� �i� 0�< < �        � � �� ��  <  �  �.  �+  �+ �����  �; ���                � � �� ��� �� �� �� �� ��  ��  �+  ��  �0 � 0                   0  �� �� < �?�� �"� ��  �                         �   � ���<D01�O�3 0 ?�>�< 0  �   <                  
�  ((     �  0  0  �?  �  	�  �  _�  �?  ?�                0�0 �3 ��  �  1  0    �,  >2  0     �                 ? ���0<� �� 3 ??��0' ��  0                             ���00<�L���  <�� �  �  <                 
$
$$,
,,,,,,",4
444444"4<
<<
D   $$$
,,,,,
44444
<<<<<
DDDDDLLL   $$$$,,,44
444444"4<
<<<<<<
DDDDDD   
$
,,,",4
444<<
<<<<"<DD
DDDDDLL
LL   $
$$$$$$,,,4
444444<<D
DDDDDD   
$$$$$,,44444<<"<DDDDDL"LTTTTT
\\\   $$
$$$$,,
,,,,,,44
4444"4<<<"<D"D   

$
$$$$$$,
,,,,,,4
4444444<
<<3<3<<<<"<
DDDDDLTL   $
$$$"$3,3,3
,3,3,3,,,,",
44444"4<<<<"<3D3D3
D3D3D3DLLLLTT
TTTT   $$$$$
,,,,,,4
444444<
<<<<<<D
DDDDDDL
LLLLLLT
TTTTTT   

$$$,
,,,,,,",4
444444"4<<
<<<<<<"<DD
DDDDDD"DLL
LLLLLL"L0 ,1&   
$$$,,,,",44444"4<
<<<<<
DDDD   ,,
,,,",44
444"4<<
<<<"<3D3D3D3D
DDDD3D3D3D3 D3"D3$DLL
LLLLLL"L   
""$
$$$$$$"$
,,,,,,",4444"4<
<<<"<DDD"D   
"
"$
$$$"$,
,,,",44
444444"4<<
<<<<<<"<DD
DDDDDD"D   
$
,,,",44
4<<
<<<<"<DD
DDDDD3"D3$DLL
LLL   
3
3$$
$$$3$$$,,
,,,3,,,44
444343434343 43"43$4<<
<<<0 $1&   
"
"$$
$$$$$$"$,
,,,,,,",,44
444444"4<
<<<<<<
DDDDDLLLT   
"
"$$
$$$$$$"$,,
,,,,,,",44
444444"4<<
<<<<<<DD
DDDD3"D3$DLL
LLLTT
T\\   
"
"$$
$3$3$$$3$3$$"$,,
,,,,,,",44
434344434344"4<<
<<<<<<"<   

$
$$$$$$,
,,,,,444
<<<<<
DDDDDLLLTT\"\   
"
$$$3,,,,3,344343<<3<3DDDD3D3L
LLLLL3L3T3
T3T3T3T3T3T3T3T3T3T   $$
$$$$$$"$,,
,,,,,,",44
444444"4<<
<<<<<<"<DD
DDDDDD"DLL
LLLLLL"L   
$
$$,
,,,,44
44444<<
<<<<<<DD
DDDDDD"DLL
LLLLLL"L0 $1&d   
"$$"$,
,,,,,",,4
44444"4<<"<
DD"D   
$
$3$3$$$$,,,,4
44343444<<<<D
DDDDDD   

$$$,,,444<<<DDLL
LLLLLL"LTT
TTTTTT"T   ,,44444<<
<<<<<<DD
DDDD"DLLL"LT   
"
"$
$$$$"$,,
,,,,,",44
444444"4<<
<<<<<<"<   ""$"$3,3,,
,,3,3,,,,3",3$,44"4<<"<DD"D3L3LL3"L3$LTT"T\"\                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ��� ��ة��  ��� � � � � � � �ύ& ��" � t ����
 �� �� � �
���� ��� ��XL �H��1 �/ � ��/  ��(�h@H�' )��. � ��. �0 � ��0 �' �# �$ �% hX@                                                                                                                                                                                                                                                                                                                                                                             <� �� E� �� �ƭ$ ���� �� �� �� �ʩ�Z  �� X� �� �̮U �{�[ �x�  �ӭ[ �\  �� �� ҩ  ��] ���K� ��  �� ��Z �0 ��L	��Z ��a � ��� �� �� �� �ۢ �(� ���� �] L1­^ ���>� ��  �� ��� �h� � �˩ �� �( ��� �� 8� ����L	�L+� �ͭ_ ���L	� �����! �ԭ` ���� �` � � ��� �LI� �����	 � �� �L]©
�' �# `H�Z��	 �� �� ��� � � � � �  �ĩ���  �� �r� � 8�� �ҩ� ��� � 8�� � � � �  �ĩ� ��	 ����  �� 8�� � � � ��	 �� � �ĩ���  �� �D� �L�� � � � �� � � ��	 �  �ĩ ��  �� i� � �  �ĩ���  �� � ��	 � �ĩ ��  �� 8�� � � �ĩ���  �� �� �L� ��<� �� ��z�h`H�Z
���� 轷� z�h` ��� �*� � �
���� 轾�	�)�� �D� ��	 ����  ��ύ& �� �x� �	 �˩� �* �d� �+ ��  �ө�a �-�W  _� H� �ީ$� �x� � � ��  ��� �$ L�ŭ ������$ L��� �* � ��+ � �* `� �L"Ů ���  �ӭ 
���� 轒� L"Ů ��� Leũ ��  �� ��` �Ʃ�Z  �� � �  ��d�[ �\ �.�b � �  �ӭ( � ��� �b �W  _� H� �� 3� wӢ ��� �( ��� �b �W  _� H� �� 3� �Ҝ  �ѭ ���l�  ��e ������ ���  �ѭ )� �I�( � ��� �b �W  _� H� �� 3� wӭ JJ���� �( ��� �b �W  _� H� �� 3� ��LƢ ��� ��`�6 �7 �8 � �^ �] �` �_ ��a ��b �V `�9 �: �; �< �= �> �? �@ �A � �]�B �H �N ����$�B �H �N `�  ��! �� � � ����! ���`�Z ��� �P� � �˩� �\� � �˩�$ �	� �P� � �ˮ  ���0 %̩c� � �  C�� � � �\��P� �ϭ i� �����0 %̩c� � �  C�� � � �P��\� ��� 8�� ��� � �� 9�L��L6ǭ �P�� ���z�`H�Z� ��  �� ��� �P� �
 �˩� �\� � �ˢ �P ���z�h` �ͭb ��L��b �/�W �( � �) �  _� Hҩ ��  �� 3� �ө.�W �( � �) �  _� Hҩ���  �� �ҭ( i�* � �) 8��+ � ��a �,�W  _� Hҩ���  ��`� ��  ���L�����L6ɭ( ���.�W �( � �) �  _� Hҩ ��  �� wө,�W  _� Hҭ* � �+ �  ���( �( �( � �) � �.�W  _� Hҩ���  �� 3� �ҩ,�W  _� H��* �* �* � �+ �  �� �L�����L�ȭ( i�&�L�ȩ.�W �( � �) �  _� Hҩ ��  �� wө,�W  _� Hҭ* � �+ �  ���( �( �( � �) � �.�W  _� Hҩ���  �� 3� �ҩ,�W  _� H��* �* �* � �+ �  �� �L��`H�Z �� ���)��&  "ʩ� �n� � �ˢ� �� ���  ��� 9� mʩύ&  �� ��z�h`H�Z� �" ��# ��$ �j�s�i� ��i � � ��"��0���" i�" �# i �# �$ ��z�h`H�Z� �" ��# ��$ �j�s�i� ��i � � �"���0���" i�" �# i �# �$ ��z�h`H�Z ��� �(� �  �˩� �P� � �˩� �\� � �˩� �h� � �˩ �U �	� �P� � �ˮ  ���= %� � �c� � �  C�� � � �h0�P� � �U �ĭ i� �U �����@ %� � �c� � �  C�� � � �P��h� ��U L	˭ 8�� �U L	�� � �� 9�L��L	�z�h`H�Z
����" 轉�# � �"�$�$�c��b��]�8�7�  C̢� � �ʀ�Ȁ�z�h`H�Z
����" 轉�# � �"�$��c��b��]�8�7�  C�Ȁ�z�h`H�1 �  ����1 � 0�h`H�  ����h`xH�Z� �c��$��b��%��]��&����� ���� ��$ � �s�� ��� � ��� Ȳ�� ��$ ��� � z�hX`H�Z�  �� �� �ͩ��� �  �� �ө2� � ����� �Ӡ � �� ��0� g� �ө+� � ���� Ҡ  .ҭW � �Z _� H� ���0�� �2 �2 �2 � �3  3� Ӏ0�1�� �4 �4 �4 � �5  3� Ӏ�3� 3� vҀ 3� ��L�̩.�W  _� Hҩ� �( ��� �) ����  �� 3� �ҩ,�W  _� Hҭ( i�* � �) 8��+ �  ��z�h`Hک� �� �c�  C� C� C̩� �� �b� �V �� C�ʀ��h`�( � �) � �  �����_ L����	 9� ��L�� �����L�����H 3� �% �% � �&  �����|�+ Ɉ��* �( �( 8�* �L�� ���( �(  X� �L�����I 3� mb �% � �&  �����/�+ Ɉ��* 8�b �b �( 0
�( �L�� ���( �(  X� �` HэX �@0L��
���� 
���
l 
��LX� m� YЭV ���V  �ͩ�LX� m� YЭ[ �\  �ѩ�LX� m� YЭa ��9�,�W  _� Hҭ* � �+ �  �ީ-�W  _� Hҭ* � �+ �  �ީ�a ��LX� m� YЩ7�W � � ���  _� H� �����  �� ���LX� m� YЩ6�W � � ���  _� H� �����  �� g��LX� m� YЩ�b �) � �( � J� 3� i�% L�ϭ i�%  H��2��/�W  _� Hҩ���  ��LЭ 8��( � �) � �/�W  _� Hҩ���  �� �ҩ�LX� �� �� �� �Щ LX� �� �� �� �Щ LXЩ LX� m� X٩��] LX�`�s �s ��c

��c �W �c � �c � �X �W ��s �� 3� ��s L\� _� H� �ޭ )� ��  Oӭs 

�� �c �c �c �c `�� �� ��LG�

��t �W �t � �t � � 3�% 8� � L���0� L�Э& 8� � L���0� L�� _� H� �� 3� Oӭ� 

�� �t �t �t �t `�Z�&  �Ӭ% � z�`H�Z�( � �) � �+mb �W  H� _� �� 3�b �� ��L�� ��z�h`H�Z�( � �) � �+mb �W  H� _� �� 3�b �� ��L�� w�z�h`�Z�. � �� ���z�`�Z�/ � �� ���z�`�Z�0 � �� ���z�`H�\ �. h`H�	�/ h`H�<�0 h`HڭZ 
����" ���# �h`Hڱ"�W  _�ȱ"� ȱ"� ��h`HڭW 
����	 轷� �h`HڭW 
��5� �5� �h`H�Z�  �Ӭ �W � z�h`H�Z�  �Ӭ � � z�h`H�Z�  �Ӭ �W � ȑ z�h`H�Z�  �Ӭ �W � ȑ � �Ӭ �W � ȑ z�h`H�Z�  �Ӭ �W � ȑ ȑ z�h`H�Z�  �Ӭ �W � ȑ ȑ ȑ z�h`H�Z�  �Ӭ �W � � �  �Ӭ � z�h`Hڮ  �Ӭ � � ȑ �h`H�Z�  �Ӭ � � ȑ � � �Ӭ � � ȑ z�h`H�Z�  �Ӭ � � ȑ ȑ z�h`H�Z�  �Ӭ � � ȑ ȑ ȑ z�h`H���  ���! h`�
��~� �~� �`H�Z�Y �7��m6 �6 �7 i �7 �8 i �8 �z�h`H�� �� �8  /ԭ7  /ԭ6  /�h`�� m1 m. m/ ma mb mV mZ )`H�Z�)�JJJJ�  C̊)�  C�z�h`�Z� �"Ȣ ���% �&  H��� �� �] �[����]  X٭b ��I��b �/�W �( � �) �  _� Hҩ ��  �� �ө.�W �( � �) �  _� Hҩ���  �� ��z�`�* m m � �+ �  3� �% � �&  HэY �@0L�
��e�� 
�e��
l 
�+ m m � �* �  3� �% � �&  HэY �@0LT�
����� 
����
l 
�* m m � �+ m m �  3� �% � �&  HэY �@0LJ�
��e� 
�e�
l 
L� � ���  ��LJ� � )� �� �Y �a � �W L���Y �Y �W  �� M� H� _� �� �� �� LԮ ���  ��LJ� � �� �� �Ӯ ���  ��LJ� �� �ڮ ���  ��LJ� �� ۮ ���  ��LJ� �� qۮ ���  ��LJ� 7�* � �+ � �,�W  _� Hҩ ��  �� J��4 �* �5 �+ ��2 �* �3 �+ �* � �+ � �a ���,�W ��-�W  _ҩ���  �� ���  �ө��. LW� �� 	ڮ ���  ��LJ�LT� � ���  ��LJ� � )� �� �Y �a � �W L+��Y �Y �W  �� M� H� _� �� �� �� LԮ ���  ��LJ� � �� �� �Ӯ ���  ��LJ� �� �ڮ ���  ��LJ� �� ۮ ���  ��LJ� �� qۮ ���  ��LJ� R� ��  �� ��* � �+ � �a ���,�W L�ש-�W  _� H� �� 3� �ҭV ����^ � �` L��V ���`  X�LW� �� 	ڮ ���  ��LJ� `�LW� � ���  ��LJ� � )� �� �Y �a � �W L`��Y �Y �W  �� M� H� _� �� �� �� LԮ ���  ��LJ� � �� �� �Ӯ ���  ��LJ� �� �ڮ ���  ��LJ� �� ۮ ���  ��LJ� �� qۮ ���  ��LJ� 7�* � �+ � �a �W  _� Hҩ ��  �� J��4 �* �5 �+ ��2 �* �3 �+ � ��� ���. LJ� �� 	ڮ ���  ��LJ٭\ �<��\ �\ `H�Z�s �s �O

��c � �?�W �c � �c �  _� H� �� 3� )� ��  Oӭs 

�� �c �c �c �s L^ٜ� �� �G

��t � �7�W �t � �t �  _� H� �� 3� Oӭ� 

�� �t �t �t �t � L��z�h` ҭ% J��% �% � ��% �  �ө �W  _� H� M� �� :� �ӭ& � �&  H�� ��,��-�L�� M�s �s ��A

��c � ��s ��s 

��Y i	�c �W � �c � �c � �c  _� H� �� ��`�% )� ��% � � ��% � �& �& � �� �� ��7

��t � �� �� M��t �W � �t � �t � �t  _� H� ��`�% )� ��% � � ��% � �& �& � �� �� ��7

��t � �� �� M��t �W � �t � �t � �t  _� H� ��`�% )� ��% � � ��% � �& �& � �� �� ��7

��t � �� �� M�8�t �W � �t � �t � �t  _� H� ��`� ��% �% �
�0�% � ��	  )ީ� �(� ����  �� � ��  ���% �ɭ �%�. )ީ� � 8i(� �
� ����  �� � ��  ��� �˩	�% �% � �2 )ީ� �(m � �% � ����  �� � ��  ���% � �ǩ�% �% �
�2 )ީ� �(m � �% � ����  �� � ��  ���% � �ǭ � �) )ީ� � 8i(� ����  �� � ��  ��� �Щ
�% �% � �+ )ީ� �(� �% � ����  �� � ��  ���% �� � �(� �� ��	 �/� �
���� 轾�	�)�� � �$ � �s�m � ��i � � ����	 0� ��� m	 � � i � �$ �ǭZ � �
��
�L�ݎ � � � �2i
���� 轾�	�)�� �d� �� ��	 �� ����  �� i
���� 轾�	�)�� �d� �� ��	 �� ����  ��ύ& `H�Z�
���� 轾�	�)�� � � �� i� � i � ʀ�z�h`H�Z�* � �+ � �a ���-�W ��,�W  _� H� �� 3� �ҭ* m �* � �+ m �+ � �a ���-�W ��,�W  _� H� �� 3� v� ��z�h`H�Z� �$ � �s�m � ��i � � �Q���	 0��� m	 � � i � �$ ��z�h`�s �s ��

��c � ��s ��L��W �c � �c �  3� i�& � �%  H�� ��,��-��.�:�/�6�"0�*L�L���%  H�� �!�,��-��.��/��"0�*L��L��L1� _� H� �� 3� Oӭ i� �s 

��W �c � �c � �c  _� H� �� 3� )� ��  ���s L� _� H� �� 3� )� ��  Oӭs 

�� �c �c �c �s L� _� H� �� Oӭs 

�� �c �c �c �s �W 8�"
���� 
���
l 
 m�V ���V  ��L� m�[ �\  ��L� m�a ��9��a �,�W  _� Hҭ* � �+ �  �ީ-�W  _� Hҭ* � �+ �  ��L� m�7�W � � ���  _� H� �����  �� ��L� m�6�W � � ���  _� H� �����  �� g�L� m��b �) � �( � J� 3� i�% LT� i�%  H��2��/�W  _� Hҩ���  ��L�� 8��( � �) � �/�W  _� Hҩ���  �� ��L� m� X٩��] L�`�� �� ��L��

��t � �� ��W �t � �t � �t �$ JJJJ�� �$ )�� �� �0L��)��L=㭂 
����% ���&  3�% m �% �& m �&  H�� �L�⭂ 
���m% �% ��m& �&  H�� �L�� _� H� �� 3� OӮ� ���m � ���m � �W  _� H� �� 3� ��� �� 



�$ �� )m$ �$ �� 

��W �t � �t � �t �$ �t � L�� _� H� �� ԍ� �W �0�0�� ��W L㮂 ��W L㮂 ��W  _� H� �ޭ� 

��W �t � �t � �t 譂 )�t � L�� _� H� �� 3� OӮ� ���m � ���m � �W  _� H� �� 3� ��� �� 



�$ �� )m$ �$ �� 

��W �t � �t � �t �$ �t � L��`H�Z� �@� � � � ����� ���z�h`H�Z� �$ � �s�m � ��i � � �-� ���	 0��� m	 � � i � �$ ��z�h`�Z�5���� ���� ��z�`H�Z� J� � 8�JJJ� z�h`H�Z� 
� � 


i� z�h`H�Z� �Ӡ �2� ��0��� ����� � ��0�z�h`H�Z� �Ӡ �2� ��0��� ����� � ��0�z�h`H�Z �
���� 轾�	�)�� � �
 �@� � � ��
��(���
 i0�
 � i � � i(� � i � ���Ωύ& z�h`Hڪ���




�& ��)& �& �h`H�Z� ��  �� ��8 �A 0N��7 �@ 0D��6 �? 0:�8 �> 0P��7 �= 0F��6 �< 0<�8 �; 0J��7 �: 0@��6 �9 06��L �� � .�]� �B ������T �- T�]� �N ������T � �� A�]� �H ������T  g�z�h`�< �? �= �@ �> �A � �H �N ����`�9 �< �: �= �; �> � �B �H ����`�6 �9 �7 �: �8 �; `�6 �< �7 �= �8 �> `�6 �? �7 �@ �8 �A `H�Z�T � �L~�(� �� � �� �� �爹�� � �&�  %̽��  C̩� � � ��  ���D �� �� H�c� ���  C�h� �� � � ��  ��� �� ��h� �  ������� �&� U�L��
� L������ �&� u�L��#� L���� �I��� 轩�  C�� �� 4�L��� 4�L�����L�� 轩�  C����  4�L��� 4�L��z�h`�� �P� � �˩� �d� � �˩� �x� � ��`�
� �P� �; )�  C̭:  /ԭ9  /ԩ
� �d� �> )�  C̭=  /ԭ<  /ԩ
� �x� �A )�  C̭@  /ԭ?  /�`Z�
����" ȹ��# ��� i7�"z 9�`Z�T ��
����" ȹ��# ���"8�7� z`H�Z8�7�& � �& �� ��]8�7� h`H�A8�7�& � �& �� ��]8�7� h`� �� ��  �� �� � � � � � � � �� �� �ύ& `H�Z�� ���Q�� ���.�� � �뭉 �� � �  �ꭝ � �뭖 �� � �  ��� �� ͋ � [�� �� ͘ � +ꭅ ���.�� � �� �뭣 �� � � � �  E�� �� ͥ � ��z�h`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��a��� �a��� Ȍ� �� �� �� � �'�� ���� ȱ��� � ��� � ��� ��Ȍ� �� ��`�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��a��� �a��� Ȍ� �� �� �� � �#� ��  �� �뭉 �� � � �� �� � � `�� ���� ȱ��� ȱ��� ȱ��� ȱ��� )
��a��� �a��� Ȍ� �� �� �� � �'�� ���� ȱ��� � ��� � ��� ��Ȍ� �� ��`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����Α �� �� �� ͯ �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����Ξ �� �� �� Ͱ �� �� z�h`H�Z�� )?	@�� �� 4��-� �� �� ����� )@��J��� �� Ȍ� �����Ϋ �� �� �� � �� � �� z�h`� �� `� �� `

������ ����� ����� ����� � ���� ���� ȱ��� ���� �� �� ��� ��  [� +� �� ����� `�K��� �L��� ��  �� E���� `�M��� �N��� ��  �� E���� `�O��� �P��� ��  �� E���� `�Q��� �R��� ��  �� E���� `�S��� �T��� ��  �� E���� `�U��� �V��� ��  �� E���� `�W��� �X��� ��  �� E���� `�Y��� �Z��� ��  �� E���� `�[��� �\��� ��  �� E���� `�]��� �^��� ��  �� E���� `LEVELcSELECT$BEGINNER$AVERAGE$EXPERT$GAMEcOVER$CONTINUE$END$PAUSE$b$PUSHcSTARTcBUTTON$VERYcGOOD$TRYcAGAIN$ENTERcSIGNATURE$��%�-�4�>�G�K�Q�S�e�o�y�B H N  PdxB H N p���





-�0�{�̓/����U���<�Ɩ\��X�֘Q��S����2�d�	����_��4�ġ����݄=����-�m����-�m����-�m����-�m����}���ͅ]�]�]�]�]�]�]�����]���݆�]���݇]�]�]��-���=�]���������}�Պ-�m����-�m���퐝�(( P`ppp@@@@@@@@00000000  �PPPPPPP                                  �xZ����   $(($xx (<Pdx������,@T					 @ Yh]eRe�e�e�e*f`f�f�fg������������#�#�#�#�#�#�#�#�4�4�4�4�4�4�4�4����������������������������� �J�K�yϧ�������E�E���������E�����������E�E�E�E�E�E�E�EЛհհհհհ����������������������������������/�D��������������֛՛՛՛՛՛՛՛՛՛՛՛՛՛՛՛�Y�Y֞՞՛՛՞՞՞՞՞՞՞՞՞՞��������R�R�R�R�R�R�R�R�R�R�R�R�R�R�R�R�mׂח�����������������������������֬����������������������������������������� �8�8�8�8�8؇؇؇؇؇؇؇؇؇؇؇؇؇؇؇؇آط���5�5�5�5�5�5�5� � � � � � � � � � � � � � �&�&�����&�&�&�&�&�&�&�&�&�&�&�&�&�&�k�~���������%� �   �   ��     
8:<> �� j� j� �� w6� �� �� w� �� �� ��    �	� �$� �� �	� �� w� j� Y	� j� w� �� w	� j	� w� �� �H�    j	� 	� �	� �	� �	� 	�    _	� q	� 	� �	� _	� q	�    _	� T	� K� K<�    �� �� j� Y� O� Y� j� j� �� ��    �� w� d� Y� d� w� w� �� �� �� �� �� w� � �    ��.� ��.� �� �� �� �� ��    �� �� �� q� w� � �	� �	�   @� �� ��@� �6��� ����@�   h	��$�@�	�� �� �� Y	� �� ��� �	� �	� ���@H�    �	� �	�	�@	�	� �	�    �	� �	� �	�	� �	� �	�    �	� �	� �� �<�   h�� �� �� �� �� �� ���h�   � �� �� �� �� �� ���h� ��h�� �� �    � �� � �� � q� d� � _�    �� �� �� q� w� � �	� �	�    �� �� W�    ��@� ��h�   ��:�*������*	�    �� �� �� �� �� �� �	�    %� _� K� �   \�	��	��	��	   ��	\�	��	}�	    #� � � � � � �   �� �    �� /2�    �
	 �
�
�
	�	�
 � 

		����#�/�5�;�?�C�G��Q�  ���  ���������  c�c�����  ��2�  ����  {�  :�  ��  j�  ��������
�!�8�O�u���  ������������������ 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P��@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____  0@P`p��������  0@P`p��������  0@P`p����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   R� �i�