&�T�6�����ƹT�6�����ƹT�6�����ƹƹƹƹ$�4�D�T�d�t���������ĂԂ����$�4�D�T�d�t���������ăԃ����$�$�$�$�$�$�$�$�4�$�$�$�$�$�D�T�d�t���������ĄԄ����$�4�D�T�d�t���������ąԅ����$�4�D�T�d�t���������ĆԆ��$���$�4�$�D�T�$�d�t���������ćԇ�$����$�4�D�$�$�$�$�$�$�T�d�t���������ĈԈ����$�4�D�T�d�t���$�������ĉԉ����$�4�D�T�d�t���������ĊԊ����$�4�D�T�d�t���������ċԋ����$�4�D�T�d�t���������ČԌ����$�4�D�T�d�t���������čԍ����$�4�D�T�d�t�����$���$���$�$�$�ĎԎ����$�4�D�T�d�t���������ďԏ����$�4�D�                 ��0�����������������0�� �   � ���3�3�3�3�3���    ���������������  �<<<<<<�? < < <<<<�  �<<<<< ��� � < < �?  �?|�\_�p�p��W?|��_ p��W�W}|U��    �p5p5\\ \\\5\5\5\5\\�  �U�5�5�������U������   ��W��ppppppppp���W �  �����\�\��� � � ���\�\������  ?�5p5p5p5p5p�UU�5p5p5p5p5p?�  �W�����W�����W�  �?U5�?      �U�      �?U5�?  < � � \\\5\�\W\_\s\�\\\�  � ׀� � � � ׀� � � � � � � �   * � ?33� *  �              �?�              @@    � ��          ?��  U�G�\��� ��  P� �@�@?� �? � �     < � <��_����? � 0����� ? � P4<40�0�0�0���@?������ L=������C�C�C�G?==�3��  � ������U��0=�������0�0�0�0����C?�?��  @���  ���==�  T����0�0�p���@�  ? �@=�?�0�0�� �@��������      P P  �� P �@������@  @U@�@�C?C=� |U�����강l��  4���?�� @U����  �?<��P��?�/   / / �� TC�C�CCCC�  CC?C�C�CCC?===\?��? �@=������ �P?�4 � � CC=�0P� � _ �   @ PC@        � \?�� � �@?�� ?    � ��Z��l l@  � ��U� � P @ lP�������Zo�����nlPl@l@�����ZAU@���@�P�P�   l l � � � ��?�?�?@�A�A���[����� ?           ��*                �
(�  � �         � � (��
          5 ����                  T    @ @        TP  ?����* �      �S�������%��*            � � ?�?
� #      @V@ J   �            # �  
 �           � (� � � ,          � � , ,�� ,@PP � �@� l � �          P9U9V��       l l  ��� P  @���o�o�l���������[�VU  @j����������V �T�������O��~�ߐ�� | � o��g�fy�v������t���f��|漹|���ttWt���W���5�u���}��P������W�� ��v�yy��nf��of�� � �A@   ^ } of��of��of��|f��vA�U�ՙwf_�G�y|f���f��f���g �^@@^A�Uf_�yf晙 o � | � � �    ff��ff��ff��of���f�� o � � �    �����?�@�@�   �    T   @ ��� � � ����������������[�z�������Z��j�P� �@   U������������_�@�U  _ ��W]�w@@@  u ��P7�7L��p��}_G@   _ T��uTP @      y]��TT�T��W  ���QA  }UWUU�U�U�UWQWA��W�����wWAu���tuuuw]_]�}��u�u�u��@UC�]�]��Wf��W�yPC@�@��uuu�u@wvyvy�w����@w } } }@}��}�u    
��� � � �ll����@@@@@l:�����A�U�������nꪪ�����@� �U����c�m:n�l�����������P@} u TP�z���@ ��\�l�@U      ��p� � �A�Э@� �    T�@   m � t � t � u � @@��EP�    @�@W�U���ut =P�� o  0 � ��]w\\pw�q�qwp� W |�\]t|�p�p����� � d �@P� ]@W��t] _�W] ] _ q�]\��U�_u�uPpu�U�U W _������/ � � � >�>�>l>l      � �U@>@>�����d@@ ��?������@�@?  � � � �@~���g��?   @@=��ff��f��?��_�{�nf��=f>��f���g曙���޻wg��gf��ff��ff��ff��ff��ff��ff���39N?S�ff��ff���f���o߰C�=��T  � W \ \5p��u�� � ���   �P� u � P @ @ @ @\�� \ \U����    t t t �@mT^�_�   *��V�U��u5@@@�U?�?  �?W�                � �   �h B  @@@@ @ @   @� �A    P  * l ���l@k@k��� � � ���+�������������>�=�>����@ o�V���� �� � �������  �  
   � �    �����٣��     � �   
�   � � � � � � = = 5 5                 �����U�9���� �@9yyyA~>���     �� �P����?�?                             ! $ � �   ( �               � � �     �*    PZ�o�����?�   @       �u�� �             @    @    P P             �?��Z�@            9    P @                 @  � 
�       PP
 �      ��* @ @ @   T@A     PP  � � (�    �   �*    ����Ƒ֑�����&�6�F�V�f�v���������ƒ֒�����&�6�F�V�f�v���������Ɠ֓�����&�6�F�V�f�v���������Ɣ֔�����&�6�F�V�f�v���������ƕ֕�����&�6�F�V�f�v���������Ɩ֖�����&�6�F�V�f�v���������Ɨ֗�����&�6�F�V�f�v���������Ƙ֘�����&�6�F�V�f�v���������ƙ֙�����&�6�F�V�f�v���������ƚ֚�����&�6�F�V�f�v���������ƛ֛�����&�                �� ����4�� ����4�� ��ްE�l��:��TA@��0���++��      ??����    � �ZE��� 3��� 3��� 3��F=[�   �����Q�F� F  ? ? ? ? ? ? �?  �?? ? �? ? �?  <<<<<�                PUP@QDUPUP@QDDUPTQTUTUUDDTP@TUTUTTTT  UU @UU TTD UU UU UU UU@U@DU@DU@DU  UU @UU @UU @UUT UUQ UUT UUP UUPUUDDTU@@Q QU DTE DUEAU@@@EEEPEEPQ@AQTDQUDT @ PDDUPU T           @P    EDDDQUUUUUUUUT@@D@TAT@@@@@@ADQDT@ATDADDQDD@TPUDDDUUUUUUUUQEQPU@UP@UAP@EAAAAU@UDPDTAT@UUDDUUUUUUUUEUEU U UUUUUUUUQUUUEPEUUDDUUUUUUTUPUPEDDUUUUUUTUUDDPPTPP PPUU  TPUU QUPP PUP PUQUQUQUQUQUQEQUQTPAPDPE@U@ UUQQDPQDQQDQUUDDUUUUUU@QUUQDDUUUUUUUUUU  @ UU @UEEU TDDDUEUEUEUEEUEUEUEDDDT U UEUEUEDEEDEEUEDPTU UUDDUUUUUUUUTUQDDEDUUUUUUUUUUTETUTDTU DUUTTTTDUTUTUDUTUDUDUDTTTDDDDTDUDUDQDEEQPDPQUUTTTTUPUUDUQDDUUUUUUUUU UDUQUUUU UUTTUPUTPUUU@T  @  @A@EUDDDDDDDDUDPEDPEDEQDDEDEUE       P @D@Q@T U @     @ @D @   @ TP   PPEDDTUUUUUUUUP Q Q  DUPQUQPUTEDDTUEDDDUUUUUUUUD@@QUUUPUDDDDDDDDUUUUUUUUUDUDDUUUUUAQAUQ@UUUAAAQAAPUUUUU PUEDDDD  UUDDDDDDUUUUDDUUUUUEUUUDDDUUUUUUA P UED@UUUUATADAAQADUUUE  UUDUDDDD UU UUQUDDDD    @  D      E@ EP        @  @        @           @    T@ @P         UUTUQDDUUUUUUU UUUDUUUUUUUUUD@EADUEDUUDTUUTUUETUEUUUU  UUUUTUQDDUUPUTUUUUUUTUQ     UUUU             E@E  UUU   @ @E@Q@U@U UEDUTUUUUUUUUU P              UATE Q A E@UPUUUUUUUUUUUUEDUU QUAQPQDE@DATU TUUUADEADEUDPEU UU PUEEUDDDEDDUUUUUUUUUUQUUAQQQQQQUQ TUDQEDEPUU@UUUQDDUUUUUUUUUTU   QETUEUUUUUTUTTTTTUUTTUUU                      Q D P     @ @                 @  @ @ U   U                UUDUDDDDDD   Q DQDDDD @         P   T @ @UEDDDDDDD   @ @EEDDD                                           @ @E       DE   E DQDT@T  D  @          D AD@       D      @D  T@DDE D@  @     D   @@DD@ D@PDD    ADQPE@    QEQQUUUQTDE    D   D @TDQQAD P@D@@       PPAQED@           @ DDDP@D A D@P   QTDD@ DD E ED            DDQ@ T T@@                @     @   @       3 3 3 0           0 3 3 3 3       ��  ��      ��  ��         3 3 3 �  �       �  � 3 3 3 3    
((
��(

(  <�5W5W5\p� ^�n�~���������Νޝ�����.�>�N�^�n�~���������Ξޞ�����.�>�N�^�n�~���������Οޟ�����.�>�N�^�n�~���������Πޠ�����.�>�N�^�n�~���������Ρޡ�����.�>�N�^�n�~���������΢ޢ�����.�>�N�^�n�~���������Σޣ�����.�>�N�^�n�~���������Τޤ�����.�>�N�^�n�~���������Υޥ�����.�>�N�^�n�~���                �� ����4�� ����4�� ��ްE�l��:��DUUUQ��0���++��      ??����    � �ZE��� 3��� 3��� 3��F=[�   �����Q�F� F  ? ? ? ? ? ? �?  �?? ? �? ? �?  <<<<<�                EETEUQDTTTQDTQUUQEETUEQQUDUATDQDQUTUETADATT   EDQQUDQQUETDUUUDDTQ QUQTEDA@D   Q    @@ @  @@A P@DQETQQEP@QUU@EDUUETUQQQ@D    EDTUQEETQEUTUUEU ETUUUUTUQTUUUTUTTUUDUUTEAQU   PUUUTTQUEUU EDPUUTUQEEDTUUETUQEEQDDTUDPEUUUUUADUQUDUEQTUQUTUUDTDPUTUEUUTE UDUUUEUQUDT UUUUUUUUUUUD EDDQUUTUTUUUQDDTUQE@TUQUUQQPEDPQUTEUQUUUUUEUUUQADEDTUEQEDUTTUUUUUQTDAUQUUUUEUUUUUUETUUETQQ@TDEQEU@  @QE@QTDUEDUQUDT DDDEUTQEUUUUQE@EUUUUDQUEDA QQDTPDPTQD DUUUUTUUUUUUEUTEUETQQUUUED@PD EDPD E AA@ UPPTTUUDUUPEUPUQDEA@ UT  E @A E  T PP@  PPPPUEDQUEUUE           UEQTDUEEE       DA      T QPPTEEDEEUUEQ    P  PDUUUPU@QP@D Q DU@ U DQETUUT QTQPDA@TDQQUUUUEPATPEUUA@D A@ @ EDTQTTQAUQD               UQTUTQQDED       TETUUUQEUTUUUUUUQDDAQTQQTDUEUUUQUEQQDATEDDUEUPPU@T QDP AD@TT@D@               UUUTUUUEUQUUUU   TUUUUUUEUUUTEUUUTUQDTTEUTUUUEUPQTEUDDUTU@UTTUQUPPEDUAEPQD@PEDD@  D@    TDD U @              UUUUUUUUQUUUQETUDU UUUQEUUUTUADDPAATUQTQDTQQUPA@P   PU @  @     D      U UUUUTUQQEUQEEPUEDTUUUUT                    @  @P A @@  @@@PT D                   @  @          @             @ P @  D@TPEEUAQ D A@TT U AP@AQ@ DD      @   P    P P E  D      D  @A           @   EEQDEQETTUT   @D@DUUUUUEQ QDQ A     Q@ D  @               P TA T@  EDD  D  P@PUUEDTQADEETUQEUEUQUQDUDUUQEUUTUDUEUQPTUUAUD@@       @ @   D     PDD@             @ T@A @UPD QADTTEUUEUTU@QPUAQED         @ @       @     E Q @ A  P              E                              3 3 3 0           0 3 3 3 3       ��  ��      ��  ��         3 3 3 �  �       �  � 3 3 3 3    
((
��(

(  <�5W5W5\p� ʧڧ���
��*�:�J�Z�j�z�ʧ��������ʨڨ���
��*�:�J�Z�j�z���������ʩک���
��*�:�J�Z�j�z���������ʪڪ���
��*�:�J�Z�j�z���������ʫګ���
��*�:�J�Z�j�z���������ʬڬ���
��*�:�J�Z�j�z���������ʭڭ���
��*�:�J�Z�j�z���������ʮڮ���
��*�:�J�Z�j�z���������ʧʧʯگ���
��*�:�J�Z�j�z���������ʰڰ�                �� ����4�� ����4�� ��ްE�l��:��UUUUUU��0���++��      ??����    � �ZE��� 3��� 3��� 3��F=[�   �����Q�F� F  ? ? ? ? ? ? �?  �?? ? �? ? �?  <<<<<�     @QPPPADQQQQUQTUEUUUUUUUUUUUEE AE@QT A@@ D APPP UUUUTQETDDQEQUTDADUU  U PDQQDTPQPUTDQQQQ  TU@TPT@TPTPTDDPTUTUDPUD TU@TPEPEQEAEPDQD@EED@DUUUUPU@PPPAPTQPETUTEDETUTT PU PUPUPDUTUDTPT @D @@@@E@ @@T        @ @Q@U@P @A@ T UP      @ @AP Q@E Q   U UQTU   D @P@E TPU@U U T T PUUE  @              P  @   P                                        @TU        DUU  UUT EUU UUUU@@  UUUU  UU TUUEEE  UUUUUU  UUUAEEEEEEEEE@D EEEUEEEE  UUQQEEEEEEEEEDUQUT DD EEUUPUUTAPUUDUDEDUEEEDUU          @ P A  @          T Q @   @     @  DQDDD D  D DTUUUU  DQDQUU U UUUU  UUUU  UUUU UUU TUU  UUUUUU  UUPUU TTTTPTQDQ QDQTTTTTTTQQ  UUEETPPTTTTTTTUTUQ EUDQ@DAQA @TTTTTTTUA@@AEAAAAAUUTTEU PUE@PEUU @   P         @@@ TU TU EEU U UPEDEEEEEEUUUUDDEUU P TUUE TATEAU @U TTETUUEEEUPDUPUD UAEUTUUUTTTTEE EDE EDE ED UU@DD@TDT@TDTPUUUUE@TD@DT@TDT           @@@@@U@PTPPQDQUTQUUAPUAUUAUUAUUEUUEUTUTUTUTUUUUPUUUUUU UUQ     @ P @ P @ P DD UDDDAAAAAUETTTTPPQPQQQPTAUPUTAUEAEUQPQEUQUE        @ QPU@U@@@@ U UP      T UU     @D P@@@ D@@@ T          QPU@U@ @@AEQDTTTETE QU UEUEUQUQUTQPPDDTUTUUUUUTUPU@U UQ Q PTED P   DDU@U@EEEUUDEAEEPQQUQUQUEUEUU  @DDEPAQUPEQTTT   DDTDDQUPTQTDQQUEDTQQQUEETTETEAAPEQQQUQUTUTUAEUDUTUQUQUQUQUUUE@EUQTPUQ@UTUTUTUTUQUQUQPEQTTUTTEQ@D P@@@@D @@@T        @  QTPU U@@@ Q TUT      @ @P Q@D U   P @QDU   @@E@ PU@U    @ UUU                                 @@P@ P@D @P@T3 3 3 0           0 3 3 3 3       ��  ��      ��  ��         3 3 3 �  �       �  � 3 3 3 3    
((
��(

(  <�5W5W5\p� ����&�6�F�V�f�v�����������Ʋֲ�����&�6�F�V�f�v���������Ƴֳ�����&�6�F�V�f�v���������ƴִ�����&�6�F�V�f�v���������Ƶֵ�����&�6�F�V�f�v���������ƶֶ�����&�6�F�V�f�v���������Ʒַ�����&�6�F�V�f�v���������Ƹָ�����&�6�F�V�f�v���������                �� ����4�� ����4�� ��ްE�l��:��j�� �T��0���++��      ??����    � �ZE��� 3��� 3��� 3��F=[�   �����Q�F� F  ? ? ? ? ? ? �?  �?? ? �? ? �?  <<<<<�UQEUUPAU UD UU  @UUQETDAEEE@UQ@QUUQUUUDQ UPQUQU DUUUUDQEUUUDDUUUU PUDDUU UEQEQPUU TQEUDTUQUUEDQUQUQ@QQDQQTQDUQUUUUTQQQAQQQQQTQAQQQQ@UUUU@ @ U@ QQPQAQQQAQQTA@ U@ @ U@ @ UUAQQPQEP EU     EEEE  PU UUTUPUEPUET@E@TTUEUEEEEEQQPUUUUPPQUPDEEEEDEDDDDPQPPQUPUUEE@EDDD@EEDD@ @EETEE  UUTUUUEDDDTAA@TAUUUU  UU  UU  UU  PUTEQDUQUQUQUEEUEU@TUU QUD UD @ @UQEEEEDPQADT@UUPTUDDUUPUDDQQEQUUUQUDUAUDP@@@ @UQUPUPEQ@ @@@EQUQUPUQDDQPUPU@TPUUUPEEQEPTEQUUUUAT QATUUUU TQ TP T P TQ T Q TQ T Q TQ@TQDUEUE@T UUUU  UUUU  UPETDEPE @UD @DTDTDETDTDTDTDETDTDTDTDEUE DUPUU  UUUU  UQTTQEEE ETEETETE ETETETETE ETETETETE EUE @U @U@TUDDTU UU @U @UUDDUU  UU  QU @UDU @UU  TUTUED UUTU  UUUUDD  UUUU @UUADT PUUUUUTUUUPUUUUUU UUAUEUUUU TTDQUETUEATUTQUUUPPTUQTTUTTUQTUQ@EUEE UUUTEUUUUU@AU  QUTUU  UUUUQUTU@P UUUU@ @@@ @@@ @@@ @@@ EEPUEE  UUTU P  TETDA@P U             @   @ P   E    EDUUUUU  UU@QQPQPQEQEAAPPUEUU           @U    @ @     @  D D@P@PTDDQUEUUUUU  UUQTUUUQU UAUUUEQEAAPAPPATPATEQEEE EUUAAQEDDEQQ@UUUTUTDTTT     QDUDPTTTTT QT@TE@T Q@TUTTUTUUU@UTATDQUUUUUUUUU  UAQ@A PTDTQUUPUEQPAQUA               U UUUUUUUUUUUUUUUUUUUU DUUUUUUTTTPTUQPAQTAATEUUUETEQEAQTUUU       @    @ @ @ @ @ P TTU@ETPQUUPUTQQTDUUU      DUUUQTPPPQU @ @ P P T TPU TUPTTTDTDTU3 3 3 0           0 3 3 3 3       ��  ��      ��  ��         3 3 3 �  �       �  � 3 3 3 3    
((
��(

(  <�5W5W5\p� �6�j�����ɿ6�j�����ɿ6�j�����ɿɿɿɿ ��� �� ����� ���� �\].147:=@CFILO�� �^_/258;>ADGJMP �`0369<?BEHKNQ �cdyz�������� �RSef{|���������� �TUgh}~���������� �VWij����������� �XYkl������������ �Z[mn����������� �op����������� �qr���������� �st���������� �uv���������� �wx���������� � "$&�a(*,b	 �!#%' %)+-) ��	  ��
  ������|}����~�������{��klopstwx��mnqruvyz���GJMPQVWbch���]\HKNRSXYdei��ILOTUZ[fgj�`a`!%)*129:AB���^_"&+,34;<CD�������#'-.56=>E�������� $(/078?@F����� �� �	

	 ����� �����������fg9:A��o�h;<BCJ��xp�ij=>DEKLS��yzqrkl?@FGMNTU\��{|stmn�HIOPVW]^c�}~uv����QRXY_`d���w���Z[abe%& '(-.!")*/034#$+,125678� �� �	

	 ����� ���������&9��'(:;�#�)*<=�"%�aLM+,>?LMZ�$����bNO-.@ANO[��������cPQ/0BCPQ\����h�m�dRS12DERS]��mljnk�eTY34FGTY^�nkifUV56HIUV_! !gWX78JKWX` ! �����opuv��|qrwx}���{styz~�� �� �	

	 ����� ����������on��QVW`ah��RXYbci��tSZ[dejr��uT\]fgks��PU^_pqlm�JAB�CDK>?�@EL*+2:6*+2F M,-3;7,-3G !"N./4<8./4H"!#$O015=9015I$#(%�&)%�'� }| �	

	 �{y�w �zx�v�������������������������������������������������������`&�&�&�&�&�&�&�&�&�&�&�&�&�&�&�&����"��$�4�D�T�d�t���������āԁ����$�4�D�T�d�t���������ĂԂ����$�4�D�T�d�t���������ăԃ����$�4�D�T�d�t���������ĄԄ����$�4�D�T�d�t���������ąԅ����$�4�D�T�d�t���������ĆԆ����$�4�D�T�d�t���������ćԇ����$�4�D�T�d�t�                �� ����4�� ����4�� ��ްE�l��:��j��U�U��0���++��      ??����    � �ZE��� 3��� 3��� 3��F=[�   �����Q�F� F  ? ? ? ? ? ? �?  �?? ? �? ? �?  <<<<<�                        @PTEUQEQUUUPUUUPTUEPU   U EUUU @Q DEETAUE @  T @UTQ TTTTTTTTUUUUUUUUUU  TQ TQTPT@TQ           @ @ @DTEEUQEUTUQE @ @ P Q UUPQ@  A  E@@@@@E AAPAPPED AT@APUQ@TQTAAU @TD@PP PE AADTA UE@UUUUUUUUEUUTUETTQUUUUUUUUUUUUUUUDUUUEUUUUTUEUUUUUUUU@UQ@DDU  DDUU D PD QUUUUUUUUUUUUUUUUUUUUUUUUEUTTUUU T@@ @@ D T PEDPDA  UTT D UQPEUTA@UP@U@ AEAA@A A A QE U@UUUDU QPE UA  AT TUUUTUUTUPUUQQUQ TAPUUQ@T@T@P UUUUUUUUUQ@EPQEAPPP QTUUQDTAUTUEDAA EUEQQDQPDADDUEDEEEDUADUQTQQEQDDUDUATETUDU@EP@     A @ EAQDDUUQUEUUEUTUUUUU  EUDD Q D D           QDDQTDDAUUUU   T U U QUUETUTTUQUDUQUDETTTTTTUUQQQQTTUTUDUQUUUUUUUUUUUUQUUQETEUUUUUEUUUUUTUUUTEUQU@E@QUDQ DTUUUDA @ E E UEUUTQUEUATTUD@ T  PQQTETQTTUUUUE E D@EUQ@U P   QPUD @DD  TUUDUQUUUTEUETUUUUEEUQEEUEEUUUU PPU PUQU AUU� UU  UUUU QU  UUUQDT          U UE AP DUQAEQ@QDQPDQ @UUDUEDEPU@UADUPTPUDQEAEPQQQQQEUEDQEDTEUEE P@T@UUUUTUQUUUUUTUUUUUUQUUUTUQUTUUUU DETQEUUTUUT U@   @@  UT QTPT@ @T@ ETUTPUDPUDQUUDUQUUUDUUEUTUUUUPUUUUUUUUUUUUUU@DUUUUUUUUUUUUUQUUUUUUUUUUUU   @       A  @@ @@@ D@UTQTQDTPQ @D@U T QTPQTAQATP @EQQDEUU          QTUUUUUUUUUU  �UUUUUUUUUUUU  @  UUUUAUQ PUR3 3 3 0           0 3 3 3 3       ��  ��      ��  ��         3 3 3 �  �       �  � 3 3 3 3    
((
��(

(  <�5W5W5\p� d�t���������ĉԉ����$�4�D�T�d�t���������ĊԊ����$�4�D�T�d�t���������ċĊԋ����$�4�D�T�d�t���������ČԌ����$�4�D�T�d�t���������čԍ����$�4�D�T�d�t���ĊĊ������ĊĎԎ����$�4�D�T�Ċd�t���������ďĊԏ��                ����U���������������������������������������� _ �               ��_U      ����<�<�<�<�<�<�<�<�    ����������������       WU��          ��_U        ��?    ?���     @U��?              ��P� @ @ @�C�O@@�C�C@@@�O�O @ @�@�COOOOO�C�@ @ @ @P_���       � � p p | �  \ �                    ? 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 � U ]��w��p�p��� � �           @PUUUPU P           � � k���%l	l	[�[�[i[U�V&X&X�VVUVU[U[UlUlU�U�VU�U�UUUU     � � �����U]���p�0�0d�e�e�e�eC�CfC�C�C�C:C��    � � � � � �                      ��>(ꨪ���� ���w�w444���^}^W��A~�t]\Wp�]  �        �� �?_��Cq55p�S_���oU[U[UlUlUlUlUlU�U�V�۬����������j���W���|�|�p�p����q�u����_��Q�D�U�U�W�����0����U��tp����]���QGAGG�G�G�G�G�G�W�U����늻�����V�UUp �|�s_}U�AGW]���������]�u��W^W^WWW��z����� ��:����Õ�UUUU9U9U9V9V9U9U�U^UU�U�W�����C��U�W\�uU � ��_���T� ttu���������Uu�Ww��U��@W �U�W��U�U VU��ZUZ�_p��Q��5���V [ l�5�4���@�P���T� �]u]�W����]��u�u@�]tt� � @ @ P PPTT�U�U�U9U9UUQ9E9A�A��E�U9����?��@�]U_�]Ut tUu�O @UU����U���UP P UU��5U<��p�_�U�U�U������:�z�z�z�^�WUUUP@@ AU^:�>�������P�A�A�G�W5]�� 9                                          EUUUUUUU              �0���UP�@}@]Q]W�^]�_��+_���Q��    ���Z�j������                 0 1 1  3 1 = � 5 7 � � �        �    0 0 0?0�?��U�U�W���P@p�p�������������������������������������������������������������������������|uCC_��C�C���                  � _�V���� 5 � � � ������l�k}kw�q{�@ �B�R�b�r���������Ґ����"�2�B�R�b�r���������ґ�����  �?<? ? ? ?<�  �?0?0?0�?<?0  �?? ? �? ? �?  �?<?0?0?0?<�  �������  �?������  ��??< ?<�?�  ��?<<<�?�  <?<�<�?�??<  �?�?�����  �������  <<<<<??�  �?�? � �?�?                ���UG]{��	FFFFFFFFFFFF�	f�]W�V�      ��UU  UU����UU  UU��      �*U� � P �U���?��[�   [�����    ��  ��      �
U&��u�^�p�������������������������p�^�u��ѕ'� � � � � � � ��        
 "   �*U%U  % *U��    U�U]  ]U��     � � � � � � � �T�d�t���������ĒԒ�����$�4�D�T�d�t���������ēԓ @ @ @ @ @ @ @U    ����< < <�<<�� �    ����         � ������ � < < <�<����?                   ���<< ���� <    ��          � �< ��  ���� �      ��� � ? ?         �������0�<�<     <�<�<�<� �<�<0<�<�<    ��<<3��       ����� � �?�  ���     � �� < < < ����     � �����     @ @�C�OL @ @� @ @ @ O�O�C @   @�C�O|||O� ?@�@�C�O  | @  
�
�
�
�
�
�
�
�
�
�
�
�
�
�
�
��ϕ#��������e'(;<��f)*=>��+,?@���-.ABk���/0CDQR��12EFST��34GHUV]^��56IJWX_`�gh#$ 78KLYZab�ij%&!"9:MN[\cd�O	P�lmn�� vu �	

	 �tr�p �sq�o� �d �ek �f �g �h �b[_ �ilm^c\` �jno �]a �$+2 �GQ �%,3 �HR � �&-4 �IS � �'.59@JT � �(/6:AKU �	 �)07;BLV �
#*18<CMW �  �=DNX �! �>EOY	 �" �?FPZ? �A� C�	����������	
��	�?�  � � �	
 � : ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`L�\�l�|���������̀܀�����,�<�L�\�l�|���������́܁�����,�<�L�\�l�|������??????????���������????��< �?�????�????��?????????�? ?�?? � ?????��??? �????��? ? ?�����????�????��????�? ???��<<<�?<<�<<�<<��<   <��<<<��?  �  �?�?  �   �< �?<<�?<<<�?<<<��������?   �<��?<0      �?<??�<�<�<�<<<<?<�<?<0�<<<<<��<<<�  �<<�<?<�3�<<<�?<�< � <<��?������<<<<<<�<<<<<<�<�<�<�<�<�<<<<��<<0<<<�����? < �� < �?���������������
���O�����'�'�/�;�K�o����c���������ˇۇ��ށ�.��.�1�U�y������	�-�Q�u�щ-�����'�g�s�}���ǋ�G���ǌ��G����g�Ǐ'����G� �?  ����������������߬�����U���U� �V� ��� W���U}��U]7pU]������_U?pUUpUU��� � ���?�? �?  ���������������_��_��_= �[? ��< W�7�U}��U]�pU]����?�W� pU� �U5  �  �   �  �?  �?  ����������������߬�����U���U� �V� ��� W���U}��U]7pU]������WU?pUU�U�  �?  < �< �� �  ��  ��������������?p��7p�5p��5�WU�UU�UUpUU5���p}�5pUU5�UW �� <� �<����?P�����@ @ �?[9�\p�p�????P ����P P�}~�z�z�~�P U P���t�]�z]�z]�z��zt���P� U  T @�Ы����t��m��z]��z]��z]��z]��z���zt�����Ы�@� T  �_  ��@����������_��wu�tWUwtWWwt]�ut��u��]�]��WW���tUUut�_u�WW@�� �_  �  @  @  �  ��@���������wu@wu�WUt]�ut��u��]�]���tUUu��}�_�@� �  �  @  PUU       ���      @���~      Ъ���T   Ъ���G�  �����ޫ�  ��������z  ��W��z��� ����z��� ��Ъꩪ� ЪЪꩪ� Ъ@����z ЪPU��ժz Ъ����A��Ъz����G��@�z������@��ѫ���� ��A���^�� ��W��z��� �����z��� �����ꩪ� �����ꩪ� Ъ������� @��������  ��꿪��_   ��ժjU   @U@�         U     0 � � W� t �   � pppp� pttttP ����P @�t�z�z��@ U @�Щt�t�t���Щ@� U  T  � @��Щ�t��t��t��t��t��t��Щ�@�� �  T ���WU��U�w���]�w]�w��wU��U�w��WU�������WU����ת�ת�W��W���U��U����WU�������WU�������W]�W]�W]�W]�W�W]�WU�������WU�WU����wU����w_��]��W�WU�WU�������WU�W}�W���}��}�w��w���i�W��WU�������WU�wU�wU�ww�ww�ww�ww�ww�w]�WU�������WU�W��׵�Wm�W����շy�o^շW��U�������W}�W��W��W�����ww�ww�ww����WU�������WU�����������������W��W��W�WU���� �� ���*�:���:+���+���+���+���+���+���+��ꬨ�:���:������������ ��  ��  �:  �:  �  �      �? ������������:���:���:���:���:���:������������ ��  ��  �:  �:  �  �  �  �   U   � !�a "@!��
B�"B
�(H��P�
@E�)��("��� `ADH�P%  @�  Q  @     � @# �  @   �    @      @       ! �    AD  �  FA�  @@��TUU���o�  k��/b��`�J�b��c��c��c�V�c�
�b��`��/b�  k���jTUUUUUU���-  h�  n�`�:`�`�`[�`k�`�:`�`�  b�  k���jUUUU� � � < � �  �000�0 ?     q ��  0 �  ��� t � t   }   } @w_�W��^���^uWg]�U]]?     q ��  0� � �t � t  }  } @w_�W��^���^uWg]�U]]?    q� ��  0?� ?���7t �5t �} P} @w_�W��^���^uWg]�U]]WU���U���W���U���Q�����?�T�@ 3� ��G ��U�WPGp@   �   WU��DT� Q��O��?��O� ����DD�?POGD@��}T�@Gp    �   V����ZUUX����UUUXUU�ZUUUVUUUUUUUUUUUUUUUUUUUUUUUUU�UU[UUUU�UUkUU��~UU�����WUU���]UUUUUUUUUUUUUUUUU]UU�UUUUWUUUWUUUUUUUUUUUUUUUUUU�W}�W}UU�^�^�]Un��o��[UY�UZ�UVUUUUUUUU�UUUUUU���������U�����UV����ZUUX����UUUXUU�ZUUUVU^UU�VUUU^UU�VUU�WUUU[UU�WUUUkUU�UUUU�V�zUUUUի�_UUUUU�]�UUUU]UU�WUUUUU�_UU�_UUUWUUUWUUUUUUUUUUUUUUUUUU]�U_�UWU{��z��^U�[��[�UU�Vi�ViUUUUUUUUU�UUUUUU���������U�����U @  TU  �}@}�@}�@}�@UU@��P��UU�Z��VU@��@��@�����@UU��Z���@�� UT P @PPUT     T  �w@��@�W@�WP�W�W�TU�@U� U� UU �i@��f@��V���F@eUP�j ��j @�  U  P   P  T  �_  ��@����������_��wu�tWUwt�_wt]�ut��u��]�]��WW����_UutUUtU��U�@��@}��@ �   �_  ��@���������WU��]�WU@WW@_�����}�_��]�tuwu���t�_utUUu�UW@��@}��}���� �_  ��@���������WU��]�WU@�_ }�@����}�_��]�tuwu���tUUutUVu�UW@�� � �  @  P_  �� ��@�@�P����P��@W� ]� �  ]�@WW�]W��UtWU���@W�@WU ]U �� P_  @  @  �_  ��@�����������Ы�@�� �� �  ��@WU�UU�UUtUUu���_t}�utUUu�UW@�� � �  @  �_  ��@���������WU��]\WU��WW�\_��\������uwt_�wtUWu���tUUutUVupUW5���@_��@�@ �_  ��@���������WU��]�WU@�_@�����}�_��]�tuwu���tUUutUVupUW5���@_��@�@͑������������������������������Y�ٱ��˓ۓ�����+�;�K�[�k�{���������˔۔�����+�;�K�[�k�{���������˓˓˓˓˓˓˕˓ە˓˓˓˓˓�����+�;�K�[�k�{���������˖ۖ�����+�;�K�[�k�{���������˗ۗ�����+�;�K�[�k�{�����˓����˘ۘ˓���˓��+�;�K�[�k�{���˓������˙ۙ�˓˓˓˓˓˓����+�;�K�[�k�{���������˚ۚ�����+�˓;�K�[�k�{���������˛ۛ�����+�;�K�[�k�{���������˜ۜ�����+�;�K�[�k�{���������˝۝�����+�;�K�[�k�{���������˞۞�����+�;�K�[�k�{���������˟۟�����+�;�˓K�˓[�˓˓˓k�{���������ˠ۠�����+�;�K�[�k�{���������ˡۡ�                 ��0�����������������0�� �   � ���3�3�3�3�3���    ���������������  �<<<<<<�? < < <<<<�  �<<<<< ��� � < < �?  �?|�\_�p�p��W?|��_ p��W�W}|U��    �p5p5\\ \\\5\5\5\5\\�  �U�5�5�������U������   ��W��ppppppppp���W �  �����\�\��� � � ���\�\������  ?�5p5p5p5p5p�UU�5p5p5p5p5p?�  �W�����W�����W�  �?U5�?      �U�      �?U5�?  < � � \\\5\�\W\_\s\�\\\�  � ׀� � � � ׀� � � � � � � �   * � ?33� *  �              �?�              @@    � ��          ?��  U�G�\��� ��  P� �@�@?� �? � �     < � <��_����? � 0����� ? � P4<40�0�0�0���@?������ L=������C�C�C�G?==�3��  � ������U��0=�������0�0�0�0����C?�?��  @���  ���==�  T����0�0�p���@�  ? �@=�?�0�0�� �@��������      P P  �� P �@������@  @U@�@�C?C=� |U�����강l��  4���?�� @U����  �?<��P��?�/   / / �� TC�C�CCCC�  CC?C�C�CCC?===\?��? �@=������ �P?�4 � � CC=�0P� � _ �   @ PC@        � \?�� � �@?�� ?    � ��Z��l l@  � ��U� � P @ lP�������Zo�����nlPl@l@�����ZAU@���@�P�P�   l l � � � ��?�?�?@�A�A���[����� ?           ��*                �
(�  � �         � � (��
          5 ����                  T    @ @        TP  ?����* �      �S�������%��*            � � ?�?
� #      @V@ J   �            # �  
 �           � (� � � ,          � � , ,�� ,@PP � �@� l � �          P9U9V��       l l  ��� P  @���o�o�l���������[�VU  @j����������V �T�������O��~�ߐ�� | � o��g�fy�v������t���f��|漹|���ttWt���W���5�u���}��P������W�� ��v�yy��nf��of�� � �A@   ^ } of��of��of��|f��vA�U�ՙwf_�G�y|f���f��f���g �^@@^A�Uf_�yf晙 o � | � � �    ff��ff��ff��of���f�� o � � �    �����?�@�@�   �    T   @ ��� � � ����������������[�z�������Z��j�P� �@   U������������_�@�U  _ ��W]�w@@@  u ��P7�7L��p��}_G@   _ T��uTP @      y]��TT�T��W  ���QA  }UWUU�U�U�UWQWA��W�����wWAu���tuuuw]_]�}��u�u�u��@UC�]�]��Wf��W�yPC@�@��uuu�u@wvyvy�w����@w } } }@}��}�u    
��� � � �ll����@@@@@l:�����A�U�������nꪪ�����@� �U����c�m:n�l�����������P@} u TP�z���@ ��\�l�@U      ��p� � �A�Э@� �    T�@   m � t � t � u � @@��EP�    @�@W�U���ut =P�� o  0 � ��]w\\pw�q�qwp� W |�\]t|�p�p����� � d �@P� ]@W��t] _�W] ] _ q�]\��U�_u�uPpu�U�U W _������/ � � � >�>�>l>l      � �U@>@>�����d@@ ��?������@�@?  � � � �@~���g��?   @@=��ff��f��?��_�{�nf��=f>��f���g曙���޻wg��gf��ff��ff��ff��ff��ff��ff���39N?S�ff��ff���f���o߰C�=��T  � W \ \5p��u�� � ���   �P� u � P @ @ @ @\�� \ \U����    t t t �@mT^�_�   *��V�U��u5@@@�U?�?  �?W�                � �   �h B  @@@@ @ @   @� �A    P  * l ���l@k@k��� � � ���+�������������>�=�>����@ o�V���� �� � �������  �  
   � �    �����٣��     � �   
�   � � � � � � = = 5 5                 �����U�9���� �@9yyyA~>���     �� �P����?�?                             ! $ � �   ( �               � � �     �*    PZ�o�����?�   @       �u�� �             @    @    P P             �?��Z�@            9    P @                 @  � 
�       PP
 �      ��* @ @ @   T@A     PP  � � (�    �   �*    ���	��)�9�I�Y�i�y���������ɣ٣���	��)�9�I�Y�i�y���������ɤ٤���	��)�9�I�Y�i�y���������ɥ٥���	��)�9�I�Y�i�y���������ɦ٦���	��)�9�I�Y�i�y���������ɧ٧���	��)�9�I�Y�i�y���������ɨ٨���	��)�9�I�Y�i�y���������ɩ٩���	��)�9�I�                �� ����4�� ����4�� ��ްE�l��:��j��U�U��0���++��      ??����    � �ZE��� 3��� 3��� 3��F=[�   �����Q�F� F  ? ? ? ? ? ? �?  �?? ? �? ? �?  <<<<<�                        @PTEUQEQUUUPUUUPTUEPU   U EUUU @Q DEETAUE @  T @UTQ TTTTTTTTUUUUUUUUUU  TQ TQTPT@TQ           @ @ @DTEEUQEUTUQE @ @ P Q UUPQ@  A  E@@@@@E AAPAPPED AT@APUQ@TQTAAU @TD@PP PE AADTA UE@UUUUUUUUEUUTUETTQUUUUUUUUUUUUUUUDUUUEUUUUTUEUUUUUUUU@UQ@DDU  DDUU D PD QUUUUUUUUUUUUUUUUUUUUUUUUEUTTUUU T@@ @@ D T PEDPDA  UTT D UQPEUTA@UP@U@ AEAA@A A A QE U@UUUDU QPE UA  AT TUUUTUUTUPUUQQUQ TAPUUQ@T@T@P UUUUUUUUUQ@EPQEAPPP QTUUQDTAUTUEDAA EUEQQDQPDADDUEDEEEDUADUQTQQEQDDUDUATETUDU@EP@     A @ EAQDDUUQUEUUEUTUUUUU  EUDD Q D D           QDDQTDDAUUUU   T U U QUUETUTTUQUDUQUDETTTTTTUUQQQQTTUTUDUQUUUUUUUUUUUUQUUQETEUUUUUEUUUUUTUUUTEUQU@E@QUDQ DTUUUDA @ E E UEUUTQUEUATTUD@ T  PQQTETQTTUUUUE E D@EUQ@U P   QPUD @DD  TUUDUQUUUTEUETUUUUEEUQEEUEEUUUU PPU PUQU AUU� UU  UUUU QU  UUUQDT          U UE AP DUQAEQ@QDQPDQ @UUDUEDEPU@UADUPTPUDQEAEPQQQQQEUEDQEDTEUEE P@T@UUUUTUQUUUUUTUUUUUUQUUUTUQUTUUUU DETQEUUTUUT U@   @@  UT QTPT@ @T@ ETUTPUDPUDQUUDUQUUUDUUEUTUUUUPUUUUUUUUUUUUUU@DUUUUUUUUUUUUUQUUUUUUUUUUUU   @       A  @@ @@@ D@UTQTQDTPQ @D@U T QTPQTAQATP @EQQDEUU          QTUUUUUUUUUU  �UUUUUUUUUUUU  @  UUUUAUQ PUR3 3 3 0           0 3 3 3 3       ��  ��      ��  ��         3 3 3 �  �       �  � 3 3 3 3    
((
��(

(  <�5W5W5\p� 9�I�Y�i�y���������ɫ٫���	��)�9�I�Y�i�y���������ɬ٬���	��)�9�I�Y�i�y�����������ɭ٭���	��)�9�I�Y�i�y���������ɮٮ���	��)�9�I�Y�i�y���������ɯٯ���	��)�9�I�Y�����i�y�����������ɰٰ���	��)���9�I�Y�i�y�����������ɱ                ����U���������������������������������������� _ �               ��_U      ����<�<�<�<�<�<�<�<�    ����������������       WU��          ��_U        ��?    ?���     @U��?              ��P� @ @ @�C�O@@�C�C@@@�O�O @ @�@�COOOOO�C�@ @ @ @P_���       � � p p | �  \ �                    ? 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 3 � U ]��w��p�p��� � �           @PUUUPU P           � � k���%l	l	[�[�[i[U�V&X&X�VVUVU[U[UlUlU�U�VU�U�UUUU     � � �����U]���p�0�0d�e�e�e�eC�CfC�C�C�C:C��    � � � � � �                      ��>(ꨪ���� ���w�w444���^}^W��A~�t]\Wp�]  �        �� �?_��Cq55p�S_���oU[U[UlUlUlUlUlU�U�V�۬����������j���W���|�|�p�p����q�u����_��Q�D�U�U�W�����0����U��tp����]���QGAGG�G�G�G�G�G�W�U����늻�����V�UUp �|�s_}U�AGW]���������]�u��W^W^WWW��z����� ��:����Õ�UUUU9U9U9V9V9U9U�U^UU�U�W�����C��U�W\�uU � ��_���T� ttu���������Uu�Ww��U��@W �U�W��U�U VU��ZUZ�_p��Q��5���V [ l�5�4���@�P���T� �]u]�W����]��u�u@�]tt� � @ @ P PPTT�U�U�U9U9UUQ9E9A�A��E�U9����?��@�]U_�]Ut tUu�O @UU����U���UP P UU��5U<��p�_�U�U�U������:�z�z�z�^�WUUUP@@ AU^:�>�������P�A�A�G�W5]�� 9                                          EUUUUUUU              �0���UP�@}@]Q]W�^]�_��+_���Q��    ���Z�j������                 0 1 1  3 1 = � 5 7 � � �        �    0 0 0?0�?��U�U�W���P@p�p�������������������������������������������������������������������������|uCC_��C�C���                  � _�V���� 5 � � � ������l�k}kw�q{�@ ��'�7�G�W�g�w���������ǲײ�����'�7�G�W�g�w���������ǳ׳��  �?<? ? ? ?<�  �?0?0?0�?<?0  �?? ? �? ? �?  �?<?0?0?0?<�  �������  �?������  ��??< ?<�?�  ��?<<<�?�  <?<�<�?�??<  �?�?�����  �������  <<<<<??�  �?�? � �?�?                ���UG]{��	FFFFFFFFFFFF�	f�]W�V�      ��UU  UU����UU  UU��      �*U� � P �U���?��[�   [�����    ��  ��      �
U&��u�^�p�������������������������p�^�u��ѕ'� � � � � � � ��        
 "   �*U%U  % *U��    U�U]  ]U��     � � � � � � � �)�9�I�Y�i�y���������ɴٴ���	��)�9�I�Y�i�y������� @ @ @ @ @ @ @U    ����< < <�<<�� �    ����         � ������ � < < <�<����?                   ���<< ���� <    ��          � �< ��  ���� �      ��� � ? ?         �������0�<�<     <�<�<�<� �<�<0<�<�<    ��<<3��       ����� � �?�  ���     � �� < < < ����     � �����     @ @�C�OL @ @� @ @ @ O�O�C @   @�C�O|||O� ?@�@�C�O  | @  ߵ)�)�)�)�)�)�)�)�)�)�)�)�)�)�)�%��B� ��� �� ����� ���� �\].147:=@CFILO�� �^_/258;>ADGJMP �`0369<?BEHKNQ �cdyz�������� �RSef{|���������� �TUgh}~���������� �VWij����������� �XYkl������������ �Z[mn����������� �op����������� �qr���������� �st���������� �uv���������� �wx���������� � "$&�a(*,b	 �!#%' %)+-) ��	  ��
  ��������e'(;<��f)*=>��+,?@���-.ABk���/0CDQR��12EFST��34GHUV]^��56IJWX_`�gh#$ 78KLYZab�ij%&!"9:MN[\cd�O	P�lmn�� vu �	

	 �tr�p �sq�o� �d �ek �f �g �h �b[_ �ilm^c\` �jno �]a �$+2 �GQ �%,3 �HR � �&-4 �IS � �'.59@JT � �(/6:AKU �	 �)07;BLV �
#*18<CMW �  �=DNX �! �>EOY	 �" �?FPZ? �A� C�	����������	
��	�?�  � � �	
 � : �����������˹۹�����+�;�K�[�                                                          �                       �������              �� �    �   ������                          �       ����������������������ɺɺɺٺٺٺ��               
 
 
 
                      















 	
    					 	 
   
   
       
       ���� �)�2�;�D�M�V�V�_�h�q�                                ������������������������������      Իܻ�������%�-�9�@�M�Z�d�     ��  � ��  �  � �  ��   �  ��  �   ���������ϼ��߼�����ϼ��/�   � ���� �� ���� �������� ���  ��� � ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������
�������l ��� � k�`�	)�)�`�(�!�|�"�#���$ �`� ��b�� ȽY�� ȩ|� ���	��`(08@PX`hp
�)��+� �V� ��=�>�?�@�B��A��C��D �	�P ���`�	)����`��恥���� ����i�!��"�|�# �`�Q ܥ��<�Ȅ4�9`�����������������������������������������
�������l +�7�����A�b�pԎԽ���C�\� � �����` j� �� �� �� �� �� � � +� �� �� �� �� � A� ��`� �!�0�"���# ۩8�" �`�<�����`�<
��m���n��� �� �ĉ��`�<
��k���l��� ���ĉ��`�<
���������� �� ��	��`�<
��z���{��� ��0����`� ��@�ĉ��`�<
���������� ��P����`�<
��<�=l Z�o�v»�����"�XÈå����2�Uĩ�2�(�b������`��2�� �	�2����L�b�

i�������`� �
�2�������


i �b�������`� �	�2�������P�b�����`�
�2��6����������<�b�d�f`� ��2�������Ýb����` 0@P`p�� ��2����LÝ��@Ýb����`$(,048xpic^YY^cipx� ��2����zÝ��


i �b����`@80(  (08@� ��2����
���b�������`� ��ý�Ù2�����Ù���Ùb����`		

ll\\LL
���| � ��2����ĝ��ĝb����` (08 (08��������2��������b`��2�:����
�������b���j`� ��2����sĝ���ĝb����`@80(  (08@8@HPX`hp8@HPX`hp� ���������I���	���`�<
��q���r��� ����`����`��0�H�`���l����� `� �/�C�0�0�
��
�0�/��/�!��"���# ۥ0�!� �" �`� �/�<i�0�0�
��
�0�/��/�!�X�"���# ۥ0�!�`�" �`� �(�=�!�^Ņ"���# ��(�(���`( � ��Ņ!��

ih�"���# ۥ�e ��`$$%��� � �(�$�!�(

ih�"���# ��(�(ř��`�	)�)�!��� �� �<��ŅP ���`�� ��`��B�>�r�����`����` ԥ��
�� -ƥ���� �� "� �� �� l� �� �� �� ��`� ���`8��!i�#���"i�$ �ƥ�0y���i��0� � �� ��Ln� �ǩ � �ܩ� �ܩ�  ���� )@� �����!�� � �ܥ�i� �ܩ�� ���� ܩ �H敩�W` ��P ���`� ����������� )�	�� �ƥ�	挥�ŉ��`������W`���:ǅ�Cǅ���b8��/e����0e� �ߥ ������%����������L`  �����0� � �� �ǩ � �ܩ�� ` �ǩ � �ܥ�i� �ܩ�� `��0��� �� �ǥ�� �ܦ���� ` �ǥ�� �ܥ�i� �ܦ���� `���� ��`�����
���ǅ��ǅl ����$�$�`���� )@� ��慦����`���`8��!i�#���"i�$ �ƥ�0&��0	 F� ��L2� �� Fȩ�  N� �� +� �� ��`��� ��`� e=�=�=�
�(�
�=�>�>�
�� �>�?�?�
�� �?�@�@�
��	�@ A� ��`�@�B��?�A��C �ĥAi�A�
�	8�A�B��V`�����"Ʌ(��U��Q�� I�� �0J������e��!����!� � � ��υ)���be(�b����� ���)�2�2`��� � `    

���r���������d ��来�)����`0S����ɍ1�	)

� ���F�� il�� i�a�x���a8��!i�#���"i�$ �ƥ������E�` !"#���P0��
���Ʌ��Ʌl ������`� � � �$����� }ʦ<��Ʌ  b�`���	��� � �������ˢ � � ������ �ʩ�  b�`�� � ������ )����إ��	�1�� � ������¥����� � ������)���С`����ʅ!� �e!� �4J� �ʦ ����!�b� �����ʝ2`  
�	)?i(�!`����ʅ!� �e!� �3J� �ʦ ����!�b� �����ʝ2`� � �$�䉐� �ǩ ��� �� �� ܩ����P ��`�)@�`�r8��!i�#���"���$��� �ƥ�0?� � �ܥ�0	 �� ��Lf� �� �ͩ ��� �ܩ�� ��  Nȩ�� �� +� �� ��`�)�|�)�W���'�0���	)��d��� � �ܩ�0��� ���`�	)�)�`� � �ܩ�	� � �ܩ5�0��� ���`���	�ͥ	)��d��\� ��8� ��������Ɉ�G�	)��d��=e���� ��� � �ܥ��`)�悥�)�������`��\̍0��e�� ���`  66      ��
��}̅�~̅l �̅��� �� ��`�	)��7��!�) �-��V �ǩ�  �ߦ 0��0�`����i�`��� � ��`�	)�8��� )@�% �ܦ��8�������� �	)���V� �����0��`��
��ͅ�ͅl "́��ͥ) �L �ǭ 0� � �ܢ��8���y͝���yu͝`�}͝0��� ����؆���V��� � ���`bjrz���!�D�	)���V�	)��1�� �ܦ�����8����ri�`���� � ����0�` ܩ ���W�`���� � �� �ͩ�� � ��� ��`���� ��`��
��΅�΅l �|��ͥ) �N �ǭ 0� � �ܢ��8���tΝ���ypΝ`�xΝ0��� ����؆���� � ������V�`bjrz���!�S�	)���V�	)��>�� �ܦ�����8����ri�`���� � ����I�����΍B��0�`���`�	)��$����� ����� )����� �� 	�挥�ŉ��`����
��i� �ܦ���υ���� 0D��ŏ���� �Ϧ���e ŏ��@I�@����
�
�@I�@�
���be!�bL�Ͻ�ŏ��������0� sѦ���8� ŏ��@I�@����
�
�@I�@����b8�!�b �Ѧ�����ϝ2���` �|xt�|xt 	
���� � �!`����LKн0�!�����!���ŏ�	�!�!��� ���e�
���Ѕ��Ѕ����� ��e�
��eЅ�fЅ�����!`�e��!� ���@�	� I�i� `w�w�w�w�wСССС��������c�S�?�+���������������  ��������������  �������������������  ����������
����������		

�������  	

�������  ���� � �!`����LҦ�����ŏ�� �����08��LЦ���х���� 0"�bő��b8��b� I�� ���0J�`�b�
�� I�� �bi�b���0J�` ���������e��!� ���@�	� I�i� `���i�a�/i����0i��`�!i�#���"i�$ �ߥ �:������V �ǩ � ��� �ܩ�� � � �ܩ ����
���҅��҅l `�Ҭ���������Ң� ܩ�F�` ܩ�G择 �� ��	��� ��ҝ0����` ��� �ͩ ��� �ܩ�� `� ���䥜��EƜ���� �ܩ� ��`�����`�C ��`� �W�� ��䉐�� ��� )������� Q�LJ��挦�䉐�`��i� �ܤ���Ө���b�!��� �� ��������� �������2�3� ���!�bi�c� ����� i� ��г��`   ������H� ��`����GƋ �� ��`����FƐ`�F�ԅ �	% ���W`????�&� �7ԝ��H�����"�<ԝR�����I�
�� �`<FPZd��0� � �� ���` �ǩ � �� ���`� � �ܩ ���`�� �� �ͩ�0��� ��  ���`�	)�(� � �ܭ�8������ ���
��)��0I�0`�	)�(� � �ܭ�i�����l�)��0I�0��� `�C0�`�D���4�9` ܩ�4�9` � � �� A� � �ũ��`��"� �����'���I����<��ŅP ��` �ͩ ��愥�)�������� `���(�	)�!� � ��枥�)�����Ս0�H�`��Ս `� � ���4�9�<`7878������������������������������������������������������������������������������������������������������
��օ�օl �r�	�ץD�!�h�"��# ۩���!�p�"�y�# ۩(�0�1� �`�x�a�;������� ��$�B�H�r�0������` � �� �� ��`�	)��`�a��� �`�	)��� �ܭBI�B���`��� �=�>�?�@�B��A��C�D�<i�4�9`�	)?�Ɓ0���!�p�"�y�# �`�� �ܩ&�B���� �	� �W�`�	)��� �ܩ'��`�	)���`��
��5ׅ�6ׅl 9�vע �

��^י0�fי`�nי���� �����`)*)*)*)*0H`p`H0   @`h`@ �� }�`�	)� �ע �0I�0��� ����� ��`� �� � ��`����`��
���ׅ��ׅl ��ة3�0�@�`�p����� ���1�B�`�r�0���.�H�`�x�@��� �������` � ?� i� �� ��`�	)��� � �ܥ�I����=؍0��� `34�	)��� ��惥�)����a؍B���`11111112�	)��� ��愥���� �����؍H���`./0/.�	)�)�`�(��� ��`� ��؝X��؝���؝����(����`,+-8HZd`b�� ��`����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������& `�ɍ& `� �!�"���#�$ �` Uۥ!JJ

�!�#JJ

�#�#8�!JJ�%�%�$8�"�&�&� ����%�� s��&��`�!eJJ��@��"�e�0 s��0��`�i0���`��!� ȥ"� ȥ#� Ȅ` U� �ۥ;
�� ��/���0� �/�!�# �۱/�" �۱/�% ���#�� s� �ۥ!�#�"��`��%��&`�/��0`�%��&`���`�I����<�� ����E�F�G�H`� ��`�  I����I�%��`� �#�!��"��#e"�#�!��`� �#�$�!��"��"�!�#���$`����/�� )�  �� �����`�/������ )�  �� �������  ��������� )�  �������`� ������`� � ��� )@�� � �� �`��0����
�'�݂�(��`�!���" Uۥ�%��& Mݠ � ��/�%L/ݱ%�/ �� ���'� sۥ�%��&�
�'�(��`�
��\݅/�]݅0` x��0Pp���� @`��� 0`��� P���@p�� 0`��� P���@p��`�!)
� �$���" Uۥ�%��&��0����
�!�݂��"�0
����/�-���0�.� )�� �1���$�_ �ީ �'�(� �/�# Mߥ#
&(�$��'�# �ߥ#�%�1�(�'� �(� �$ �� ���!�˥'�# �ߥ#�%�1 sۥ�%��&�
�!�"Т` �ޠ �/�# M� �ߥ#�% �� ���1�!�� s��1��%��&�
�!�"��`�� ��`�/�/����0`�� )
�� ��ޅ+��ޅ,l+ ����ߥ-�/�.�0�8�"�)��
��L�� 5ߤ*��e
��0e/�/��0`�-�/�.�0�"8��) 5ߥ*L�ޥ-�/�.�0�"�) 5ߤ*��L�ީ �*�)��*e
�*��0�)��`�� )�,� ��#jjj)���#

)0��#JJ)��#***)�#� `�H�
��\݅2�]݅3� �1�2=�ߕ)����� �#=����#)�#���� h�`�0?���� � )@���!����� `� � �%�/�#���#�%`��!���"��0�$�����%`� `�!8��%`� � � �* �X�Y���Q�V�W`������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � xآ�����&  R᩠�  � � � � �6 7��9�� ��ԥ6���9� r�LM� �� � � ]� ���6L,��� ��� ��������������`�9�$� �9�4���0�P �� � �� � �  �� ��`� �� ��0��` ���������������
���T�� �%��&� � ���%L��%� �� �ۥɐ���X��`��%� �:�:� �;� �!� �"�: �������`�4�w�& �4
��e��f�� � �/�*���@�0�0�) �۱�# �� ���)�0����)�) �۱�# ���)� ��L<�ɍ& `��������������������/H�0H�4
��?��@��#)�
���%ȱ�&� � �� �%�/ �����
� �� ��L��h�0h�/�/i�/��0�*�*��� �*�0�/iX�/��0� `�/i.�/��0`�4
�����l  � � � � � � � � � � � � � � � ��� �$�&�T�6�����&�T�6�����&�T�6�����&����"��6�j�����
�6�j�����
�6�j�����
��ϕ#�H�H�H�6��	�6 �� ���ah�h�h@ ���J�N�O�P�Q� �R�S�T`�P
����J���K`�Q`�O���N�O�S`�P�S�� �� �J�LȱJ�M�R�L�U�R��ȱL��R�������Q� � � ����R��ȥT���T�U�RL�����R�ȱL�U�T�RL���R�ȱL�RL��HJJJ�S�R�hL��XȱL� � �� h)� � �� ��� � ���� �S� � �� �RL��n�V0)

����V�Q� �b�R�d)� �c�S� �T� �X�X�Z�d�M)x�IJJ�e�b��c�=��9�d0 �b8�e�b�
�c� �b�c�b� �c� L�eeb�b���c�c��� �b�X�� � �W0

����W�i�( �j�) �Y�k�* �Y�	�Y�� �* ` y
 o� {o_: D�i�- � o �
 o
  K�W���U�A�'�s���������� �� � �	� ��� � <� �� < <	� ��� < �� �� � �	� ��� � h	T T���� ���0 }@ T@ } }	@ @T@ } �T hT � �	T ThT � }@ T@ } }	@ @T@ } � �@T�����<�\<   �A� ��o�����_��9�+�j� �� �� �� � ���w��� ��7� �� �� � � � �]�	����g���� � � �� � �@� �t�M�G�#��� � �� � �� � � �@����� � � � � � �  � � � ��� �� � �� � � �� � � � � � � � � � � � ��  � � � � � � � �K�E�7���G���g�{�"�q�����E�������Z�F���2��� ��	� � � � �o�=�Q�/����+��� �!� � � ��-�����[��0��#� �A��� � �� ������R����� � � �� � � � ����� � �� � �� � � � � � � ���C� � �@� � � � �� � � � �� � � � � � � � � � � � � � � �����������S�r��!�#�� � ��C���������@������ � � � �� ���;�w������ ��� � � � � ���'�I�`A�!�#� � � �� � � � ��\��S�A���� � � � � � � � ���@�� � � � � ��� � � � � � ����� � � � � � � � � � � � � � � � � � � �� � � � � � �� �  ���1T 1@ ���1 1T 1@ @T}1� 1T 1@ ���1 1T 1@ @T}1� ��@�� �  T !�  ��@�� ��!@ !�T�@�  T  � �@���@ T 1� @   [�[�T}T@T@� ��! ���@T}�!}T@!} }�����}T�����!  @���}T@ �!}  T}T@T@� ��! ���@T}�!}T@!} }�����}T�����!  @���}T@ T}!�    G�G��� � � ��} }� � �� � � �� �� �@T} 	} } }T@ 	  ��T T� ��� �  �T}�� � � ��} }� � �� � � �� �� �@T} 	} } }T@ 	  ��!T}� ���A@@   Q�Q�!@ T@  @ } � } � ��� < � < �0 !@ T@  @ } � } � ��� � � } �0 "< \< � � � � � !� �� } "�` "< \< � � � � � !� �� } �p   -�-�@� �@� � � �!!!.!@	T	@	T	@	T	@	T	@	T	@	T	@	T	@	T	@	T	@	T	@	T	@	T	@ y�y�T	@��� �	@}	T < T	@��� �	@}	1�   ���1}�!}!h!@ �   �0�!@ �A�@ 1h}!h!@ !  !1@h!}!hA@@ 1��!�!�!}!�  !}1@!h!}A�@ 1��!�!}!h!   �0��! �A@@ 1}�!}!h!@ �   �0�!@ �A�@ 1h}!h!@ !  !1@h!}!hA@@ 1��!�!�!}!�  !}1@!h!}A�@ 1��!�!}!h!  !1@T!@!�A�@   �����@� ������� � ���� �  ����� � �   �    ����#X` #X` "�` "�` "�` "�` "<` !�` !�  !�  !}  !T  !@! � � � � � ��qk_UPG?85/*( # ]�]�� �� ��}� �!�0 } �} �}T@ T } < � �� ��}T }!�0 @ T �!}  @T}!T @ T@ T@� @T@ } �} �}@T �}@ � �� ��}T �@ ��@T @T @T�!}`   ���& ���Q�V�W� � � �* �X�Y� � �< ��Z�[�[� �\�]�a�^��& �a�^���^ �� ?�\����]����ai<�a��`�Z��Z`�Z�\�>�]�:��8�\ ,�i0�_�i �`�\�����_����_�i0�_�`�i �`���\���  ��\�a�.�]�*�D ,����ȑ���� ��i0��i �����Z� �\�_��a�Ș g�\�a����\`�\`�[��[`�]�K�]�G��8�] ,�i��i ��i0�_�i �`�]�����_����_�i0�_�`�i �`���]��� ��]�a�0�]�,�D ,��ȱ����'��� ��i0��i ���ߩ�[�]�a����]`�]`



}��_���i �`�J��� ,��e��i ���_���`� � ��@�� ��������`H)��G�hJJJJ�
ei@}W�` 0`��� P���@p��      

�� �|� � �����`� �/ ���� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� � �