L��L���1��;��7�/�9I�9� n� ���	� �` !� <� t� ܙ �<�� �`�9���1
��X��-�Y��.l- ހR��א��B���߇g��z�=>?@IJKLMNOPQRSTUVWXglmnhijkopqr{|{|}}~~����������������������������������������������������������������������Ʃ � ������ P碖� � ������������'�/�)�����
��d�����L����(�A�$�"���#�!�;��'iH�'�(i �(���(���'���/�'#��

� ��, 㢩n�P���Q �LƁ� � �G�K��=� �C)����F�J��P� �d�#�<�$�2�/�  ?� ��擹F�� ��
 ��LÁ

�  � ��/�/�H�.�)�)�	��$�"�#i�#�!LP�� �)���#�!�$i�$�"LP� �� !� <� t� ܙ 򙥢� j� � � 	��1`� �� 	��3��2� �;������ �� ��H��` 0���>��)��1�1�> ܙ� ����`�)@���� �� $� 8� ���	�1�� �`� ���������� �� O� �� {� ׃ u� � t� � �� �� �� ~� -� �� ԏ���'���#�@�������=��� ��1� �����Ƙ��� <���� t���� ܙ��� �`�����������������������������.<�`     @ �	t�Q@ddQ@����7��)�1榢 � �)��}���0



� �� �*�� ��䥐�`�*���"� �}���*�	� ��� ���*�� �Ͻi��~�� � �� � � �ȑ� �i0��i ���H 좥�)�����+�i��#�i�$ ��+�#��$� �h�L��i��~��H��)



�� � ��/� �����Ƚ�����/�˥/���i���i��إi0��i ���  *来�)�5�<��/��!���e;������ ����/8�!�! 좦!� �	�!�/� ��`I� i+�+�/�U���� �L*��?��@�
�
�A)����A�2�<�A�?�
�@�����@�;�@�? n� ���� �
�1`�` !
��)��!��)�������8�Ņ� Y����)�� �`�<���e;��#�� ��)e ����\��⨥ٚ��ڄ�� ���<����F����?�Ĉ������ѯ���F��;������0������������� �����Q����M����U����1� ��`@Z@@ �' ��((��8�JJ���8�JJ�


ee�`�:�:�	�� �:��� 6� ��`�����)��<��`��!���e;������ ����/8�!�!�!� �	�/�!� ��`�/�������i8�0�������ڹ�����i8�0��Ő����� � �U������(� � �ȑ�(��i0��i ��� ��������1�`慥�)�� ���������� ���"���! � ��`�=��1� ��`��1`����>� �B�C�D�E�F���������1�%慥��
�7� ������	

in� Т ���� � n���� ׈�1�1��` ���1�`�YƟ�����3�2`��=�<�A� �B�C�D�E�F���@����>������1�<��܇�? !� <� t� ܙ ������
� �`�A�&�<�A�@	� �3��2`�@i�+ 㢩���[� �`�0���� �3��2`	
� �� �/ 㢦/�z��+0�e�i�+�
ią�[� ��/�/��ة���[���+�	�@�<�A �`����  ����� �/ 좦/�͈��+�
iʅ�[� ��/�/�
�� ��`��)�
�������`� �P�0�F�d�N��� )��	�
)���䓐�`� ņ�LO� V��
�.Ň��z�i	���0٥.i�.Ň��Z����Z�x ��L;�� �������`������F�����d� ������ i���
i���<i���2i��L;��8�	���0��.8��.Ň���Z�� �Z��x ��L;�� �������`���� �����F�����d���� i���
8����<8龙��2� ��L;��
Ň�� V�� �-ņ��xȱ�0�-i�-ņ��Z����Z�x ��L;�� �������`������� ���F�����d���� i���
i���<i����2i��L;����0��-8��-ņ���Z����Z�x ��L;�� �������`������� ���F�����d���� 8����
i���<i����2i ��L;�� 8�JJ��
8�JJ�


ee�`��)���ŉ������) �` � � �`斥�)���)����� ������`� 8�JJ��8�JJ�


ee���0��)��

� �H�^��"����! � �h�L�� j�� �ƕ�!`� a�L���� j�����"�7� �L����8����� �L����i���i �L��� �L������� � ��i0�����`栥�)���)�
������` ���� �����d8��d 4�L��������� k�Lˌ��� 4������"�7ޖ޾L��ު��8������� ��L������i�����i ��L������L����8�JJ���8�JJ�


ee�`�� ��������.�

i��-� �-�� ��-�i0��i ���`�����H

��� � ��� ��i0���h�`<��<��)����� ������`� �&�����"���
� �ƕ��`� �P�L4�� � �	�Ri� �K�
��	�Ai��:�F���P0�8��Pж���PЯ�P8��PФ��(�<��2� ��Lč�ē�LЍ�����H

�� � � ���� ������ � ��h�L���i0��i ��ҥ�)�� �������`���&������"���� �����d8��dL����ݖ�	�iݖ���ݪ�	�iݪ���Ƚ�������.�H

i��-� � � ��-� �����-� � ��h�L���i0��i ���h`�ld��� �P0�䓐�`�P�朩�(�2��<� �� ��L4��P)�սP)}F��%�� �2�"�<�!�H�F�� ��L�� � �h�L4�������� �P��䓐�`� 8��0�������
8��0��ؐ�����`���������� �*���䥐�`�?8�0��������TŇ���`��
����-���.l- $�P�z�z�� ������(����i0����i ��ƌ���)���� �1 !�`� ������(����8�0���Ǝƌ���)���� �1 !�`�:�:)��������� ������i0��i ����ƌ�� �1`����ƍ`�`��
������ ��� ����  �������ǐ�撥����1� �:��`0484840�:�:)�;� ������2���H�P�0攽2�"�<�!h� H�H � �h��䓐��h���` 6�� �P�
0� �P ���䓐� ��1� �������`� �� ���������� k�Lf�0��� 4�Lf��F�J�
� yB �B �
��
�B �C i�C ȹB ��`  ($(,4048@<@DLHLPXTX\���������������푕���������������H�2�"�<�!�F



� �Z

e }(����� � � ��L0� � �h�`� �P0��䓐�`��(�<��2� �� \�L?�� �������`��8� 0����8�
0����� �

�� ��������� Lc�� � ������(��i0��i ���`� �P�,0*�x�� �x ��Ln� ���
�����-����.l- �䓐�`��6�p���ד�Z�� �Z ��L(i)�(�n�
�<8���<�2� �2 ��LZ����Z ��L(i)�(�n�
�<i��<�2i �2 ��LZ����Z ��L(i)�(�n� �<��2 ��LZ����Z ��L(i)�(�n� �<�<����2 ��L��n�F���(i)�( ��L)��`� �� O���� t��:�:)�%��  㢩 �+������ � �� O���� t�`�������� � �ȑ���i0��i ���<i� � ��� �/�)�A�$�"���#�!���(���'�/�'#��

� ��, 㢩n�P���Q �L��� � �
���


�  � ��/�/�H�.�)�)�	��$�"�#i�#�!L�� �)���#�!�$i�$�"L� �� j� � 	��1`� ���@�� �������Z��`Y@@@� &*&$( 㢩 �'��(�'���$���#� ��+�#��$� ��(��'���#�#��#i��#�$i�$���'�'����@�� ��#�+ �@��&��'�+ �Y�����%�+ �Y�����)�+ �`�"+�",�-�.�-���""".��123�.../-�0���0�.�0�0�0�-�58.��97��"..�6�-�-�-�"8�6�"��"��6�".8��0�<�""�-�-�-�".��;�0�:�8"�:�0�0��6�0�VUSSRPPPPOMMMMMLLLLJJJJJJIIIGGGGGGFDVVVUSSSSSSSSSRRRPPPPPPOOOMMMMMMMMMLLJJJIGIGVUSSSSRRRPPPPPPOOMMMMMMMLLJJJJJJJJIIGGGGGGGGGGGGFD���������������������������������������������������������������������������
��������������������� $O$+2 㢦<�5��(�2��'� �/�!�'�0����������+<��
)�+�!�0�1�/�/�;��@��!������� �+��@��!��+���+ ��'�(Ш`		 � �+�%���&��(� �'�'�
iF��B�����+�	�<�+ ��(��'��`>BFJNRVZ^bfj>?@?@?@?@?@?@?@?@?@=[eeeeeefeeeefeeeeeed@>@>@>@>@>@>@>@>\\\\\]\\\\]\\\\\?=?=?=?=?=?=?=?=bbbbbcbbbbcbbbbb@=>=>=>=>=>=>=>=>=>?^______`____`______a 	
 (88HXXh|| 㢦<����/� �#�@�$��'�( {��<����/���#�A�$��'��( {��<����/���#�A�$��'��( {��<����/���#�Y�$��'�( {�` 㢩��/� �#�[�$��'�(�( {�` 㢥=�'� �/�/
i��[��'�����+ ��/�/��	�'���'LG�` 㢩[�����+�?�!�
��
�!�+��i�! �!�+�[��� ��+�@�!�
��
�!�+��i�!�[��"� �[��$��!�+ �` 㢥>i�+�\���� �` 㢩 �/��'�\��/
i���'�Ai�+ ��/�'��`  (.26:  $(,.4:@FHNTV 
$(.28<@HNRV\bhntv@@DFYY@@SUSUSU@@SU@@SUYY@@@@@@YYDFJLSUYY@@JLYYDFSUDFYY@@YY@@DFDF@@@@DFDFDFDFDFYY@@DFSU@@SUYYYY@@SU@@YY@@@@DFYY@@DFSUSUSUYYSUSUYYSU@@DFYY@@DFYYYY@@@@YY@@SU@@SU@@DFYY@@DFDFSUYYDFSUYYSUYY@@SUSUSUSU@@SUYYSUYY@@SU@@DFSUYYDFDFSUDFSUDFSUDFDFSUDFDFYY@@DFYY@@DFSUDFDFYYDF� �� � �&� �&
� ��  ���&�&�&��� ���&� � ���� �&�  �&� �&� �&��� �& � �����& �� �&��� �&� �&��� �&��� �&�� � ������ �&� �&��� �&�&��� � ���&��� �&� �& � ��� ���&�&� ��� �&�&� � �&�&� �&� � �&�� � ���&� � �&��� ABGHEFABGHCDGHABCDABGHEFABABABEFCDCDCDEFABGHEFCDGHGHEFYZEFstyzuvststyzuvyzuvyzwx��uvyzstuvwxwxstyzstwxstst��wx��uvyzuvyzwxuvyzwxuvstyzwxYZ��wxwxststwxst����uvstyzwxstuvyzyzwxuvuvwxyzwxstuvyzuvyzstuvwxuvwx��yzstyz��wxuvyz����uvyz����yzuvuvyzwxstuvwxYZ��uvuvyz��uv�<��,�T�;�?��/�@�8�/�(�/�蚅�����+ ��/�(��`�;���/��8�/�(�/�X���^���d��+ ��/�(��`�;�+��/�,�8�/�(�/������������+ ��/�(��`JJOOORRUADFFIIJJMMPPRSSVVXDDDFFFGMMPPPRRUXSUUVVVCCCDDDFGGGJMMOPRSSSUVVCCCCDFGGGGGIILLMMMOOOORRSSUUVVV��$��
��������������������������������������
"���������"����� $

$" 
  
"
" "" 
 







                                                       * 0   F                     �<��>���e;�����2� ����/8��! 좦!� ��,�+�/���U�� ��!�/� ��`              
                                       "   0           8   >




















SSSSSSSGGGGGGMMSSDDJJPPPJJJJJPPPPPGGGGGGGMMMMMMMDDDDDDPPDDDDDDDDDDDDDJJJJJJJPPPPPPP�����������������������������������������������������������������������������������  &.6=UUUUUUW]]Wbehmhmrxrxrxrrxrxrxrebebeb�����������������������������<���`�%�e;��(����� � � ��*�䥐�S�� �~��?�Ѡ�T�$��i�w��~�ʡ����ĥ��`��[�� ������������`	
 � �/ 㢦/�����+�
e/iɅ�[� ��/�/���`
 㢩 �/�/����+�
e/i΅�[� ��/�/���`��%���&`���%�̅&`�+�%���&`�%��&��+)



e��i ��+JJJJe���-��.� � �� ��)�)% ��) �)  ���E)�)LC��%)������-���.�� �i0��i �е`� � �/����+� 
e#��$� ��(��/� � �'�ܩ � �#i��#�$i�$��`��������)��LR���)��L�� Y������'��(�� � � ��� ���(��i0��i ���`�
�4�	�	 ��� ���Ȧ;�@朩��Bi�B� �B�
�	�
�B�C���
��

�  좥�!��" �`��)��m Y����I��E�H�^�������� ?�h�ȱ�����^�������� ?�`��i���i ���(��  �`ȱ������H��(��  �Lv�L� Y��H������^�������� ?�L�� ��( �h�ȘH������^�������� ?�L(��� ��(��i���i � �hiH�������^�������� ?�L`��� ��(��i����i� �h�ȱ�����^�������� ?�`�� ��(��i����i� �` Y��H������^�������� ?�L���� ��( �hi	�������^�������� ?�`��i����i��� ��( �`�������5��>�I���=�=����=�`��	�早�`�?i�?�`���`戥�������`扥������`�>�>�
��	�>�`AAAAAAAAADDDDDDDDDGGGGGGGGGJJJJJJJJJMMMMMMMMMPPPPPPPPPSSSSSSSSSVVVVVVVVV��������������������������������������������������������������������������,�R�P� �Q� � �R � ����� � � �P�+�"��!� �� �,��,)��!�!�ݥ!i~�!�"i�"��`� �	�
�	� �
�� 

i� �


i�
`  %+38: 
#&)/4:?DJSY\b !!(,26:AKQW]bjp̩ҩ٩ܩ����������
�����#�,�4�;�?�E�H�K�P�V�[�`�f�k�p�s�w�|�������������������������̪ت������������������#�+�0�5�8�;�@�E�L�S�Z�c�e�c�k�q�t�c�c�c�w�|�����c�������������c�c�����c�ū˫ҫիثҫիث۫ޫ�c���c������c�	��c��c��#�+�3��c�7�;�@�E�c�c�c�J�O�T�_�e�k�r�c�c�y�����c�c�c�c�c�����������c���c���������ìƬɬЬ׬ݬ��c�c�c�c�c����c�����	����#�(�.�c�1�8�?�H�c�O�c�c�U�U�c�Y�]�a�e�j�p�x������������c�������̭ԭ������c���%�%�%�*�/�/�/�c�4�:�c�c�c�c�c�c�>�A�E�K�c�O�R�c�Y�^�a�e�c�c�c�c�c�h�c�o�v�c�{�������������������2�3(3�3#�(8�!2!�#3�2"�6&�(8�������6(2��$��4��#�3�4$�!4�2%�&7!�6'1��$42�"�"�2�(8��7(1��8(�8(�&6�3$1��(8�2$2�$4�4$��1%4�2�2$��5�%�7'�"24$�2"�"2�2"�2"�3�"�4%�&8"�7�'�&8"�24��&�241�'�62(�6�&��&6�#3��4$�6&����8(�3#�#3�!4$1�4$��"2�5%��6&���3#�#3�4$�!%51�"5#�#3�!11!���#3�"4"��&6�3#�!3#1�1#2���#�3��!�1�1#3!�!��1�1"2!�$2�2�3#�#3�����2"�(8�%5�6&��$�4��2�"�����21#�"2�21!"�%1�4�%5�2"�"2�"2�"2����1!�"2�1!�2"�3#�1!�!1��#�3�"�2�2%5"�3$4#�1�"�2�!�6&�4$�$�4�"2���2"�#�5"�#4!�$4�2�#�3#�1�3$�4$�&6��1#3!�!3#1�4$�2"�����2"�#3�1!�#3�3#���!�1�&6�4�2�"$�2%3���1"1�5%��%5���#3��!%51�$4�4�$��&6��6&���4$�2"��2�"�'2"7�%4$5�#6&3�8(�8(�8(�#�#�3�3�"���2�1��#2���"��6&�2��!8(1���"��6&�2��!8(1�$4�4$�22"&4�322"&1�$422""�!422"%�3#�3�#��3#�"�2�5&1���!1���$�#3�4�3#��3�#�1!�$4�$4�$4�"2����2"�$8$��2�"��#4!�4$����H�H�;�<��(��yu�
����-���.�$�y��
��ꨅ-�먅.��yg�
�����-����.��-"���� ������-)

�n�h�h�`JJJJ��ZL� 	 #%(*,.02357:=>ACDEGHIJLQTVY[^`adfghjmprt                                                         		

		
  		
 	
	
	VSAVDSSVSVSASVSAVJAAVJADADDVAVDDVVDDDDDADSVSAAVAVAVVADSSSASSASVDAVAAVVAVSVDAVDDSADSASAVSSSSVSASASVDADDSDDSDDAVDAVSDDD���������������������������������������������������������������������������������������������������������������������"""
""""""""""""""""""""""""""��
�����-����.l- ����ǲ��ݲg���� �`� *��
� ��`�= <��@���=�� �����` ߇�0�`�> ܙ� ���` א����� [��<����P��	��� ���PLĲ  ��.l9l9�.�   � 0 \ \ _�^�z�����3�ôǵ׭?���׫>����� �    �� ? 1 1     � 0 \ \�_�^�z��  55��?�ï������� � � < < <���??3 3 < < <  ��3�^�_�^�^�z��  5 5���?���� � � L L p � ����?�        � \  \ \��;�� 5 5 �/���Ǭ߫�ǫ׫������ �    �3� ? 1 1     � \  \�_��:�� 5 5 5 ��?�ë���������� < < <���:>3 3 < < <  � \ �_�^��:�� 5 5 5 � ��?����<�<� L L p � ����>�?      ��W�G�W�W�_���  5 1 � � � �   � ǀ��;�� ���?�        � W�W�G�W�_���W  5 1 � � � � ���_  3 �  � �� ;  ��?      � W�G�W�W�_p�� = � � ���: �C������ΰ�  : :  3 � � �� � p \   ; � �? ������� ���k��� �      � � � � ��� ? � p \�O� ; � �? � ����^ � � � p o �    ��� � 3 0    � | ^?N�0;�� �? � ����� � � � �  ��:�?0����?׿;��   � 0 _�]p�^�z�����?�õǵ��>���<� � � � �    �� ? 1 1     � 0 \0\��^�z�� 55��>�������� � � � < < <���??3 3 < < <  ��3�^��^�^�z��  5����?���� � � L L p � ����?�       � l \ \ \���:�� 9 5 �/���Ǭ��Ǫ���?��������:0�? 1     � l \ \�_���:�� 9 5 4 ��>�ë�ת���������<�< <�0�? 1     � l \�_�^Ӟ�:�� 9 5 4 � ��>���������|<�<p � ���~5W�        ��[�W�G�W�^����  5 5 � � � �  � � � ǀ��;�� � ������ <      � [�W�G�W�_����  5 9 � � � � ���_  3 �  � �� ������ ?      � [�W�W������ = � � � � � � �C���������  : � � 3 � � �� � p�_�_�_ { � �? ����������� � � � < �  � � � � ��� ? � p�_�o�� { � �? � ������ � � � 0 � �    ��� � 0 0    � | ^ ���;�� �? � ������ � � � �  ��:�;0����?׿;��   � L \W㧼[���� 5 5����;�>w�_��l�wi_l���  �ڮ5]	�b�X3�    � L\W���w��{� 55� �3�>������l�7E_,      K�7�	�b�       � \ \�7����� 5 5����;�>s�_��l�wi_l���  �ڮ5]	�b�X3�    � \\W�W�7��{� 55� �3�>������l�7E_,      K�7�	�b�        � � � � � � �  �<  � 0 �?  �0 0� 00�  � 000�?0  �� � � � � �  <33�00000  0030�03<0  �000�  �000�    �0 � 00�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`L ��1����権 ��`�1
��'��-�(��.l- =�u�ACA�
�
2 � ��F���������<�:���+��2�.��<�1�� �4��
�7��P�
�n�1��`� � ��*���� �	�c�� ���H����	�� �� �/�/�c�)

i<�+�D�$�

i��# ��/�/�	�۩ �/�'�4�+�'���#�~�/
e/iG�$�i� � �*����?�

i
�T ��'�/�/���� �/�0�+�'���#�~�/
e/iG�$�i� � �*���"�?�/

i
�T ��'�/�/���`����������       ��P�0�>��)�権����`� ��� � e� �� ؈ d� =� � 
� ޅ >� �� �� ׂ � H� s� �����������Ƙ�@��`権��`斥�)���)����� ������`����� � ��i0��������!�5� �L����8����� �з��i���i �С� �Й栭P� 0��)���)��<��� �������` ԃ����i�����i ����<����)�� �������` ԃ���������ޖ޾��<����)�� �������`������"�� ���祚��	���������� �Lꂥ<��� �*�����`� �~�#�i�$� ����i��� �*� ��:攥���,��=��P� ����� ��`�����
��D�i���~����������H�$�4� �<��0��8��������L��T��P�+ ��H �h�L,�������� � ��i0�����`    
  		<��<��)�`��ŉ�K����E�) �? ੘�%�̅&� �+��(�!��"� ��(��+�()��!�!��!i~�!�"i�"�ԥ��� ������`� �&�����"���� �ƕ��`LV��P��0��<��T ���� JɃ�������Э��8����*о����������8�
JJe���8����*В� � �<
�� y�� �
�y��� ��
y����y ����� � ��˰ �<���������P�
� �F��L������� � � ������� Lm��i0������������<��@�P�;09���5���1� � �<
�� y�8�0����|���
y�8�0���`ـ����� � ���`�<�B�P�=0;��)�5���
�,���)�������
��tL�����<���i� ��L��`� � �څ�	�R����K�
�� �������� i��i���
i�����<i����2i���<i����2i��� �������`���"�� ���� �L��� �������� i��i���
i�����<iB���2i���<iI���2i��L����ݖ�	�iݖ���ݪ�	�iݪ�桩 ��`������� � � ������� `�i0����<��-�P�(0&��)� ����g������Z� �
����M`� ����A� ��� � ��������-��� y;����
i���;�m<���2i������L�� "',3 	


 
	 	
 
�<��`����L�����}�� ������.�� � �.�ʇ���O�������!� ��������Ti���ii���!����a���!���Ti���ii����.�.� ��暥���� ��`�P��0������)�쥠��� �������`������ ���!��������C��`�<��9�P�402�)�+�2��<��<��H� � ��������i0������`�(� � ��������i0������<i���2i��� � �ȑ��ťi0������04880�<��L���H��)�>�k�$���#��1� ����(�#��$� *��#�#�(��()��#i|�#�$i�$��`�^��+�4������%�̅& �����6��2���.���*�A8��0�������V8��0��������`��(�#��$� ��(��+�#�#�()��#i|�#�$i�$��`�<��&���"���Z�P�0����� i8��0��`����攩�� i�?��T�M�i�?i��~���U� � �����*`� � ���� � �*�
�*�� ���~��i� *��T�U�*Ɣ���� ��?�A�A�T�V�~��΀�i�k`�T���+�l�%���&�~i��~��ii �i� �`�� � ��������i0������`�<�)���
��c��-�d��.l- ����������݋������+�J���_� �1�_�B�`��n��`� �<� ����n�`� �<� ���`� �
�<i��<�2i �2� ���`� �<� �	��`� �
�<i��<�2i �2� �����n`� �<� �����n`�
�<8���<�2� �2�
���`� �<� ��
� ���n` 
���������������� 	      	  
	 X\� � � �* ����� ����� �<��&�2�$�<�#�F�� ��L{�����+ � ��F`���� �� ԃ���� 숦<�b�� �<yd����2yx��������������
���`8 484048484 4808 048 48 4004848404048�� ���%�̅&� �������
������ ������2��3`���5�� ���������ν��$���#����5��+�� �� � � �#����� �#i0�#���$���4��)��/��(� �'�#��$� ��(��/Lr��+�(���#�#�ޥ#i~�#�$i�$��� �<� ���`� �<� ���`�<�#�2�$ ��� �<� �"���`` 66
��    �P��0Ǧ<����-q�й�l�%���&�c��(�e��/� ��FI�F��l�+�<i��#�2i�$��2�$�<�#�)��i���a��+� �'�'
e#��$� ��+�(��'�'�/��#i��#�$i�$�Х<�`�F�g��+�<�#�2�$��(�#��$� ��#�#�+�(��(�
��<�#�2i�$�֭�
i��+�<i��#�2i�$��(�$��#� ��(��+�#i��#�$i�$�� 8�JJ��8�JJ�


ee�` $(,(�<��6�P�10/�)�7 ��F�F)�F��������+�2�$�<�# �`������罭���)����ƫ�<�#�2�$ ��`�܅%���&` H��G�$���#�܅%���&�<���+��(� �'�'
e#��$� ��+�'�'�	���(��#i��#�$i�$��`                                   � � p p��3��      ������                                                                �_��� � � � � �^��_� 7 7 7 7                                                                 ������\������S����7�5���ַ�                                         � � � �      ��������C���+�������������ɷ��4�������      ���������         ? � � ������������ � �����������WUWa�b���3��������z{��������������������������$~� �������?�   � � �          郩��Η�� � 0 _��G�������w�{������?�?�?�?����k�j�Z���� 7 7                                              ��w�������������?�7�7�7��2�5�9�6                                                       � � p p 0�����u���������7:�8w�w]W{WzW�C                                            0 0 � �        ��чч7\7�p��C���G�G6�5�00                                                               � � p p��3��      ������                                             < �                Wu��� �   � ��֞�y� 5 6 6 9            � � �              �������� � �      : � ���:���/�n�_\�m�\�^Sn���7�5���ֺ� � �����:��� :                      � � � � � � ���������G����-���^����鵹�����:�ί���:   ���j������         ? � � �������� W � � �
�VhZ���f��`�j�﫳�����9����������2�2�,�������T%�I�iIeJ�¤~*
R��=    � � �          郩��Ϋç�ܬܫ�>�7�w���-ލw�{������8�6�1�?����k�j�j�����7�>��                    � � �    ��:�:����� �wMǝ�-�7lw\��9�2�0�4��2�9|5�6���� � � � �     � ���� ;                           � 0 0 0^����w+�+������5:t8���N�M�MzC�C                                            0 0 � �        ��W՗՗7\7�p��C���W�W6�5�00                            ���������������w�w�w�w�w�w�w�wU����������z�z�����_~�WUUUU�U�������_����������U�V�Z�j�k������UUUU����p��p��UUUU�������3���3����j��U�}�׼׳���?��?��?��?�ꬪ�����������Uw�w�w�w�w�w�w�w�^�^�����竷��k�U�U��m�N�6�7���UUUUUUUUU����N�Թ��������n�[�p��p��p��p�����3���3���3�����}�U�U�}�׳׼�}5?�?U5U5�?5?�������[���6�6�w�w�{�n����3�m�m�uquq���VWV��W�UUUUUU�U������UUUUUU�V�[�.��5y5yM]M]CWDWŕu�U���嫹V��n�0��UUZUoU�����朻���Z鯾�k��_6p���?��?��?���?��\���p�_WUWU��֯u�ulul]l���?�ƱƱűűű��?��kkk[[����Ϭ�����l�l����?�������?���k�k�[l[l[l[l���?�ƱƱƱűű��?�����������?����:??��?�6W��S�pp��3��s�3|�omUm�����ƱƱűűű��?�^�WTUS�S�NU��o4UU}U�UU���U���l�?�������?���_�O�;��3�[l�����Űſűű��?���|�\�>��_W������?��U�����������z�_WUWU�?:�6�5�5�5�=��?�������S�S�S�S����N:N:N9N9N9N��?������������N�NSNSNSNSN���?:�:�9�9�9�9��?�������S�S�S�S����N�N�N�N�N�N��������??��?�6W��S���Sup��3���s�3���?�9��?���ӔӔS�S�S�S���^�WTUS�S�NU��o4UU}U�UU���U��l���N�NSNSNSNSN����_�N�:��39�9��?�����ӰӟӔS�S�����|�\�<��Ny����??��U���l4l4l4l4l4�p�p�l4l4l4l4l4�l4l4l4�p�l4l4l4l4l4�        �p������ � � � �  ; � �? �����>�:�:����p��� � � � ��:�:�:�:j:�:�� � � � �  ;����? � ������������������� ��:�:�:�:�:�:�� � � � �  ;����? � �������������� � 
 �  �:�:�:�2�"2" 0  � � � ������>�� ? � �/������������������ ;�?? 1 1     � � �������s�� ? ? ���>������������>�> < ��:�?�:�?< < <  � � ��������2�� ? ? ? ���>�������N�N�r � � ��׿��?      ���������������  ? 3 � � � : ��l�����������������C�     � �����������l�  ? 3 � � � � ���^��s�����<�� 3 �?�*� �      � ������������� ? � � ���3 �C�C��̪<��< 0   ? � � �� � � � �  ; � �? �����>�:j�����p��� � � � �j��9�6�ڪ�:�� � � � �  3 � �? � ���:�:�:j9 � ����z / �    �������3�0�;< � � � ��03�� �? � ���:�:����  0 p � � ��:�?������Ӫ3�<�; < � ��Z���lk��? ��@:95�����W��lk����Z � �����5�9@:��?  ����V�l�[\C � ���9���C[\l��V�� �W����9���   � ��Z���lk�0�  �p5��<p���l����� � �����7>�j3�#�<<    ��|�l�[\G0S � ���9�?0����������_ � ��� ��4   ��UE��eeeee��Pժ�A�A�A�A�A�eee��UEUE����A�A�A֪�P�P�������W���������DU�ZQYQYQYQYQY�����WW����QYQYQY�ZDUDU��������lUl�l=lU������:U9�99U9�:��WUGGGGG\��U������9�������������������:�:�:�:�:�:�������������������������:� � �������������? ���:�:����������������� � ������:�:��?  ��������������� � ����:���ꫫ������������ ������:����   � � � �  ;����? � ����������,           �:�:&2&(      � � � �  ;����     � �  
                0                                           � �         UDWD  @  DDDDDuT�QQGDSQG�Q�D5QUU�� ��5 5�5�UUU���W�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU          @  @ � �    DDD^^U�U��ꀪ �  QUUUU�����
� �MDQGDQDD�G�5�5 �5 �pp\_U�U_�@_=@�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU  @  @    D@1�T�TSDNQN      (��E�@U@ePfPJ�J�jDQ�ީ:��e�:e�� |� ? ��D�QpD�QUUWU|UU}UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUDDDDDDUUUUUDNQ:T9U9U:U~���U�U)U��"�J��D�HTUD�eD��D9Qy����:p��|\jGp0�W�����UUU�T=QT� � Q�U  � � � �P�U�UUUUUUWUWU^U^UWUV�Z���>�GUUE�����D�WD\qDtq�D��D�����U�U5D�Q�TU�U���� �����>��U��z��=0w� s�Ϋ0�TWQ�T�UUU�UuW]\������UUWU]U^UWUWUUUUUUUUUUUUUUU]u]�mU�U��ժU�U�Ut�^D^QWU^�^W�U5U_u� W�  �0|��� PW�����ݻ���PŪ)��G���@�p��[����*\�rUrU�U�U�U�U�VUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUU�UU�UU�5 7�=p0<p p?�ѫG�DDQUUUUUUUDDQUUUUUUUUUUUU�UUUUUUUUUUUUUUU[UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U_=���UUUUU5 ��� �   �� �U1WUUU�_7�      U�U� 5        ��?            }U�_ �          UUUUWU�U _ �    UUUUUUUUUU�_p ��U�U�U�T-al�����UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUEEULT0UqT0ULUULUUUUUUUUUUUUUUUUU�+�F+kD��J�D�UUTUUUTUUD��j�UUUUUUUUUEU�D��UUUUUUUUUUUUfU��UUUUUUUUUUUUUUUU���U�U�UDUEDaD �0�O�2�ʈ)f&SUDUQUTUQUTUSUGUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�������D�[�j��D����2���c��h�ff��f��)fʙʦ���ff��hjc������(τ�af����(�#�����h*�(�#�#;;�ULTUqT1UqTUGUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�����*EkmE�����3�<?�� �
�U���(;;<;�� L
0(�(��������!<I������ ��mW[gGgG:�:lNlS[�Q�P	UUGUUG\MN9O�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU��U��U�UUEUUUUU��*�)�þ�ݯ��
u�u��z��F������޿ު�  g���κ>����@�B�ҎЎ��o'o�J��BN09�x�4�t�3�ӵ�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUEUUUU�����k���    � 0�?�\�+��� 0�  0UU�� <� � 0 ��Uo�[�] � � �����v�u6�o� }� �����,���)R�� �� ]U{U^U\Uz]]w�]_]UUUUUUUUUUUUUUUU�W�Wm]m]t5\�WUի^W���]խ�uUߪp�UU������������_UU��W���_����UU:�5W:��|�|U�����������uuu������������]���ZU��UUpW�U:W�U�UuU_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_UUU�W\�_�^�WUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUkf��k��͵�����ըVUYU������������UUUU�����������
UUU�_�\�_�z�z\{UUUUUUUU]UmMm5m�UUUUsUU]U]�}�]UUUUU�fՀe?��ffUUUUUUff��`��� �W�^�^�v�p
_�U_Uu��ufՙUgU�UgU]��4?�9t6i5i]�]^��*\�W�Uuev�yfv�__U{U��UUUU�߫�=T�SuƵŵ��n�l_�]k}��f_�]g~�]���Wu���]yU��g����e���W�W�T^U^UzUvU�UfW�]e^UuU�UWU�U�U�U�U�����UU�ߪު����ߙu�Uu�_�^�^�_�_��������UU���~�[����wUu�w����go����_U�������vUuU�_]����������T�T�T�S�S�T��ę]e]�WeWYW�U�U�UU�U�UWU�U�U�U�U�����U����o�o�o�k�_�_z]�_�^�^�_�_�����U��߫ޯ߻�������^����n�g�������������䷓��mz-�-�M��m�m�������;�;�;�;���tUtUtU�U�U�USWS^U�]��_�������������[U[�[�Z�Z���_�_y����ץ�e������z����᭑c���9�峔��j�1a1����e��>�0�署��͐Ð�R�I� �����:����2�3E>���:�yd��f��f�yjr�嵑�B�F��U[][��V
U�U��� �R��eeX���B�M�0��� �$�$[%[a<	<���:�:��iE)������`��C����S�S�:�9(�ZCD�9U9F9R����#�#ZΪ\_�W�W�U�U�UzU}[�Z�U���jժ_���B$	!�H�������W�@�E��jZ�U��_���l����Z�kJ��տZQ��rA�@V����p�7������������f�Y��%�'������Z��d��� �z�__U^UWUWe�Z_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUիU�UUUUUUUUUUUU��UUUUUUUUUUUUU����^�WUUUUUUUU�p�_uu�_UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU     � \���_��           �Z�              ?        � � � � �               �           ��__�     � ��5_?�5_:L��W0�0�0U�������Zի�n��U���j��k� =�� � � � �0��������������j�C:<�    ����W���V����U諥:�?���U��T�� � � S � 0 �����Z����Z��Z����j����������}U���z�z�N�C�@�U��?��������j����z��V��Z����Z֪j���� � � ? 5                  �j<��� < �      ��j�j��:�: O L ��U�U��幕�U�WU��j������ > � ��=�=                      �? � � � � �    �             � � � � � � �  �������m�m�m���� � : � � ?            �  �  3        � 3  3 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`�3������!���"���� ��%���&� �!�$� ���!�#� ���!�) ���� �/� �!�����)�+LU� ���!�+ ���!��+��, P�� ��/�8�� �$�#i��#��$�#��$���$��8� 
e#����,�� ��L=�`�!��"`  �����        ��� �� �� 	�   	  �� � ��          � �� ��     �  �              	     ����� �  �	        � ��	��� �  �      � � � � �� �!  �   �         � � � �   	  �	 � � �      �   �  �  	�   !� � � �"            	     ����� �  �    � � ��� � �      �� �	� ��   � � �	��             �	������ � 	      ���������	�  � �  � � �	� � � � �!   �        �   	 �������         		 � ��   	��  �  �  	    !� �  �   �  	�"          �������  �        � �	�	�  � 	���� �   �  � �����	    	 	     �    � 	 � ��   �      �      � �      	 � �  	 ��      	� 	�   ��	�	�� �     � 	����� � �       ���������       �� �	� �	� !     �	   	�   ��􀀀 �  � � ��     � �! ��� � �  �	� �  ������"   #                      ��  �!  ��		�   񃃃�    	�   � ���         " 	�	   �  �� �� �    ���  �	�����       �	��� �� � !   �    �	�	���    	�	 �     �� � 	   � �	      ��            	   � �     �       � !          ��      	��      �����  ��   	  ���           	   ��  !  ���	         	�	����! ���� �  �     �  � ��� ��        ��� ���   	� �	     �       � �	�  � �	� �  �         � �� ����� 	� ��	 � ��    �    �    !  �� ����" �   �  � ��     �  ���  ��	� 	�  ������ 	  �      ��	� 	   �    �!  ���	��  	  �    ��     �� 	���  	  ��	          	�	  �� � ��! ��	�	��  	  �  	    �    �� � ��  �� � ��    �  "          ��  �   ��  ��   	 ��   �� 		  �	�� 		  �    ��!    �� 	�	�          ��  �� �    �� � ���	  	�   �������� !        �������� � 	��	 � � ��� � � � 	� � � � ���� � � 	 	� � � � �� � � � �� �   �!�         ���������         􏉏�����      	��	��	� 	��	��	�!       �      �� �	��  ��	� ��     � ��� �     �	����   ��		���       !     �      � ��  �� 	 �  ����� �  		    �  ��� �  � ��� 	      	              �  ����	��  ����	��            ��	��   ��	��  !      �      �  � � � �     �	�  �	�� �     � �  �	� �	�     � �!�	�   �  	      �  �	��  	 �� �� �� �       	  �  �	�� �  � �� ��! �   �" 	 	�		 		 	   		���� ����     �������  �      � �����! �     "�        ���	� �      �  �����	�     � �  �	� � �  � �	���             ���	  � �   !  � � �� ����   				� �� ���     	  � ����� "      � � 	�	    �     �������  �        � ������ �       �������� !            �   �	� ���� �	� �����	�        ��	��	�� ��	��	��        �   ��� 	  ����� �  �  �  �       	���			���	     	� ����� �         �        �������� 	 	 	 �   	 	  �  ����� �     � � ���� � �  !   �           � � � �  � � � �  	 	 	�	  � ��� �  � � � �  � � � �               ��������	         	��������         ��������	                 �    			    ��	�	�   ��			�       �  ������      � 	�������	   	       	                 �     	 ���      ���  	             	     !       �      �	!����� " �	   �  ���� �	    ��	���	�     �� �����#	      $����������        �������� �	�    �  ���� � �	�     !���	���	�"    �    �      	        	     �    ������ �       �  �������  !    	�                           � 	           	     	 �     !    �  "         	 	 	 	���� ���� 	 	 	 	 ������� 	 	 	 	 ��������        !          	�	�  ���� ��       �  � ��� � 	�   �  �� � � � !  � ���  "��  	        � �����  �     � ����� �  �	�	� � �	 	  �  ��������!                 ��	��	����	��	��        ��	��	�� ��	��	��   ��       ��             �������! � 	 	 �  �	�	�  �	�	�  ��	 	 �  �������        "    �     �   �	�!  �� ��     �     � 	����� � �      � � � �         �       �	    � ��� �����   				 � �������      �      �	    				 �   	    			      	    				�			 	   	 	 		  		 	  				     � �    � � 	 � ��� �� 		   	 � 		��� � �� �   � !�������      	����������        !���� ����        ����	  	   ��� ���� ��  " �	 	         !�� ��  	 	 � �  � ��	 	  	 	 � �  � � 	 	 � �� � "            �    ��� �   �  �   � �	�   � �	�    � �	�   !� ���   ��  �         �      !  �   ��  �  �		   �   		 �  ���� �   � �         �������           ��������         ��������         ���������   	  	  �<�
�����!����"�ǐ� � � �-��.�!�-�!��"�-��.��H�� � ��`
���ޒ@  �VY\_�nqtw�PWZ[`cfilorux}�IQ[[[adgjmp[[[~��J
"[[��K #[[��L	!$[[��L[T%(+.147:=@CF��NSU&),/258;>ADG��O  '*-0369<?BEH��
���b�!���� ������/he�MM|�]^��������k�svv�RX������z{����� ���� ���������@  ���	��
��
��
��
��
��
������'-39�?
{�  (.4:�@
|�  )/5;AGMSY_ekqw}�  *06<BHNTZ`flrx~�  +17=CIOU[agmsy�  ,28>DJPV\bhntz��  ������������������  �
!�#%  � 
" �$& @ �P��   .<� 
!/=J� "0>K� #1?LW� $2@MXb� %3ANYcl� 
&4BOZdm �	'5CP[enp�		(6DQ\foq�
)7ER]�*8FS^�+9GT_i�,:HU`j�-;IVakUUUUUUUUUUUUUUUU            ��������                            U�U�U�U�U�U1U1U1U1U1ULULULULS���37U<U������@��1\<����CS�SuS�CULUU0T��  �          UU�U�U�U1U1ULULULS�Ӭӳ�ӾS���ԭt�t��Wt�]�����U]UW�WUW�W�W���z�z�ާ^�_�wT��_]U]�_U]Uu��U���Wm}k�ZUUUU�U�����5�4 � � L   0 0 0 �      TUSUOUOUMUMUMUSUSUSUTUTUTUSUNUOUNUNUSUSUOU7U5O�?�@?UuUUzU�U�U�U|UpU�UW�WW�UUUUUUUUU�U�U�U�U�U�>�9   4 � SL050�    4 4 5                     �  S � ��^0�0�L�L�L�L{L]LU0U0U�k0�0�LULULU�W�~�갪UUUUUUUUUUUUUU�UqU\U\U����U�U�U�U1UEUUUUUUUUUUUUUUUUU��3?,���Õ�UU:U:U�U���唥S�S�N�O�N�:�:��^_^UWUWUW_�_UpQp��U  0 � � � � � � � � � � ����T0W0W�|��0 0 0 �L=L�OU����տU��������U�U��������^�^�W�W�UUUUUU�U_�zUUUUUUUUUQU ��}UU�����������WU�ZW���0�<���1=1�LU�U0U�k�e�VU�Ul�l��ղU�VȖ [ [ ��          UW}U�W �0 ? 5 � s=� @    @@� 8�?���8�8�8�?���U�ի��ժ_�p�p���p�_U�WU�U�_�z�_�U_�U]UWW}~��W�^�z�z��UUUU�� ?� \���U�UUUUUUUUUU U�@?ZժZ������������������ꯧ���V�U�U�U�U�U�U����گ��g6�9�5ZU�oU�U�ZU�V�[ � @ @           @ UUUU�U?�    @ �@iPV�eYY     @TW��߷��z���z���U�U^W�U}UWZWkW�׷}�^�V՛U���_�U�U�U�U�W����������^�^�^�s�s��>�; :  CU<U�T*S�O�N�S�T�T�T�T�S�S�N�N�S�T�T�S�SSS�T�T�TeUUUUU����WWUVU[�m�m=�   5 4 4 5 5 EU_ � @   VU      @U_�
�EZU�돫a�X���  0�7�UuUu}]W�UyUz�n_�U{U{�~����_UU��ꪪ���������_UUU��= �p<\�WUUUUUUUUUUT�:�:090��������9 9                          U�_u��U�TTP� � � � � � � � � 5 � ? : : :  0 � � �]W]�5U?U�U�U�կ����������U�UUU�_�z�^�WW�U]UW_�pU_�ի������U�TUSUMUMU5W5W�W�\�lUlUlU�U�U�U�U�U�V�YlV�Y�f�Y���Wܪ�����W����<W � � W � �                    UUUUUUUUUUUUUUUU      : ? 5 5 � � � � U�_UU���:�:TUSUMU5U5U�T�TUSUSUSUMUMUMU5U5U5��U�Vz[z�UzZz�U�Z��Uު>�    ����                   ��������������������������������������������������������������������������������������������������������1
����-���.l- �~�� �:���1`fi����%(+.147:=@CF&),/258;>ADG'*-0369<?BEH������������������������������������            *� )�%��2�3��� �<� �B�C�D�E�F���������>`�:�:)�<��%���&��(急�)����l��/��#�/���+�C��#� P��#�#�/�(���`��)��|��/�$�(� �'�J�$���#�/���+�'
e#��$i � P��(���/�'�'��ک �'�#i��#�$i�$�ǥ1
��U��-�V��.l- ��W�������� �  ����� ��   ��������� ������� �  �������� ����������  ��������� ������� �  �������� ������� ���� ��������� DDDDDDDDDDFGGGGGGGGGIJLLLLLLLLLLDDDDDDDDDDFGGGGGGGGGIIIIIIIIIIIJLLLLLLLLLLDDDDDDDDDDFGGGGGGGGGIIIIIIIIIIIIJLLLLLLLLLL��������������������
�������������������
�
�������������������
�
  J)*� �:���<����P�����Q�1���+��%���&�G���Ҝ� P�`�:�����:)����P� �+�ΤPLٝ�1� �:`�:�:��0��� �:�P� ٝ�P�]��+�Ҝ��G�� P��P�Q�� ���1`�C ʐ �� ���3��2���<�T��?� �@�����<�A��=� �������V������������`�����:�:)����P� �+Lݝ�PLٝ* ;�<���� ����� ��<��`	 !�<��� ��� �מ�@��� ��`�1
��@��-�A��.l- i��'�c�����������������������������������%���&�B�$�D�#� �'��( 墩B��T��<i��+ P�D�$���#�	�( 墩V�$���#��( 墩Y�$���#��( 墦<�L��+�Y��������� P��1`
�0���9�<����uB�B�
��
�B�C������B��<��
�� ���1`��3�2�<`� ��@��$� � �(�. ɢ�G�����U� �@��. ɢ� � ��U��( ɢ�1`���%���&� �+�I�$�#��(� �/�/
e#��$� P��+�/�/����(��#i��#�$i�$�Щ ���������1` (- 3=FPYbf=ktF���F�������@CEUW[BVYVX[UWYVYVYUWYUWY[VX[�HDJ����B�����B�B�Ă�"
 

��������������� ����� ���������� ���� ������������������������������������ ������������������ ������������������������������������������ �������������������������������������������������������� ��������� ������:�:)�A�������e���1��-����*�1� ��� �+��
}��ՠi ���%���& P��`欩 �������欢 �/��HH�Bi�H������(h�+�/
i��[� P��/�(��`�0���4�����`�)��(� � �������.�ՠ��� ɢ��(����1`� � ���.�����i0������`� �/�/
e#��$��'�O��+ P��'�/�(��`                  ��\�L��eT\P���j�j�V\ \Tld\�����  ��� ���������L�P@P�U�����i�@�O�L�\ΜΜ��� �� ���V����@�@�����j̪ͪ�Z����Yͪ��� ���  ���Z���A�A�A�����ll@\T���L�L���  ��  ��@�@�E��P���� P @ @P�������UVA@@��  �� @��j��������ê���T� ����ϪΩΩΩΪ��� ���  ��l \ T���l@ L�����Al@l@��  ��  �� @ j ��A���_� @ T�UA���[_��|�����  ?T��U����A�A�@ΐΕΪΪϥ��������� ���� ����?��� 3 , Ti\i�j����L�L�i, 3 �@�K?����  ���j���ZdT@��0�0�5l6�6\51�C@ @U�j�����  ����?����i�T8005V9�:�:�:�:Q:E558V����?���������^P
��^P��
^P��
^P
����
^P�����������^��^�P�

��

PP
����^.,^-,�/�*������P�
��mP,�,
-�,.P,.�,
-P,-P,
.�,�/�*������^�����S���
���P�
x�8xP8~�
�P��������P�

�P
��
�S
���S
�P
P�

�P���ꪪ����P�
���P�
��
���P��P�
��
���P���ꪪ��(��.N�(�B>{A;(��;({�;(�B�(���A��A��������;�z�?N�((�B(��((B�(�B(�B(��((A���O��*��������(�B����(�B-,�.(,�.,A-(/��(���
������;
{P;��8
��8xP8��8
xP8x�8
�P8
x�8��������������>�_��S���

���S��_�о�>�����⪢����P����
����P�
������B�P;�P/
.�,
�P������ � 0 0 L L � �������0�0�0�L�L�L�L�L�L����������������������������<<<<./� ���������������S0� 3       �  C��0��C�����������������     � � �      ���_�_�<�<  ���������������WW��                    � ?� P@��������������?�?�?�?�             ��??  UT���������������������������������     ��  UU������������� � � � ����������������  ���P1u� � � 1 1 1 1 1 � � � ����1�1U� ��           ��0TL�@�?0�         ��  > � � � � � �� CU��u�	��������L�L�L�C���������� .���������  UU����_�����������.�� ����        � � 1 0          ��?  ��0]0����� � S C L L L L C � �����0��C���    �  �  _ ���}�}������� � � �               � �P TU�u������������  ��                    �  �_��_����������������������������� � �       �����       � � � � � �       0 � 0���������������<<,< < . �� <   �        �?�?�? ? � ��   0 1 � � �1�1�1�1�1�1�������������������������� � ���������������������C��0��� � � �  0��L�U�  �    ��������U� T� ���������U ��?   �<3�0300�  � � � � � � �  �<  � 0 �?  �0 0� 00�   �0�?   �?  � 00�  �0 �00�  �? 0   � �   �00�00�  �00�? 00�  � 000�?0  �00�00�  �0   0�  �000�  �?  �  �?  �?  �     �0 �?0<�3  000�?000  �� � � � � �  �     �   0�30        �?  <33�00000  0030�03<0  �000�  �000�    �003�3  �000�0  �0 � 00�  �?� � � � � �   000000�  0000�   000�033<0  00� 00  00� � � �   �?  � 0  �?        �                  � �  
��� 0   < <             < <     0� 0      ��  ��    �0 0��   �   �*�*�*�*�*�*�*� >             ��  ��  ��  ��������� �       ����������      �?�?�?     ����������������  �?�?�?      ����������      ?�?�?�?�?�?�?�?��?�?�?   ���?�?�?�?�?�          �?�?�?      ? � ���?���������������������,�23�23,��������Z�������Z��^Z������^Z���Z��^Z��^Z��������������^��^��ZZ��Z����Z��Z����^.�.^-�.^/�*���������nZ.��Z.�.�.�.�.�-Z.�.�.�.Z.�-Z.�/�*�����������[���[��[�������Z��x�������^Z��������������ZZ���Z��Z����[�ꫥ�Z����Z��ZZ������ꪪ����Z������Z����Z��Z����Z�����ꪪ�������j��ni���j������{i��{i�������j��i�����������ii������j����j��i���ji�������k����*�����j���i�������j��.�.�.i-�.�.�.i/���i���
��������{i���j��{����j��x����j��x����j��xi���������������z־�o֯�֫ii�������֫�֯�~������⪢��������i���i��j�������B��;�˪/�.Z.��Z��������� CU��u>�9������  UU����_���� CU��u���������  UU����_�� � �������                  ����  �GGGGGGG�  ����DD��    ����������?� �����W?�����������������?�� � �?�����������    ��DDDD�� �̫ͬ���0�0�0�0�0�0�0�0�0�0    ��UUUU��  ���3�s�3�s�3�p 0�O�3�s�3�s�3�s�3�s� p�0�s�3�s�3�s��  ��������    �0�0���\�W� ��           � � � � � � � � � � � � � � < < < > . . /   @������������������1�4�4�4�4�4�̼�����of��of��of��of��of������        ����.        ���� ���������0�0�0�0{{�z�^�^�������W�W�U�U�U��쪬��U�U�U{U{U����������ff��ff��ff��ff��ff������    ����ff��ff��~~���ý�ff������    ����ff��ff������33��ff������    ����f���f���g���g���f����?�    �U{U{U{U{U{U�U�U�U��������������WUWUUUUU������UUUUUUUUUU������UUUUUUUUUU������U�U�U�U�U�������UUUU��5353535353��WUWU��gf��������U;U;U;U;���{��? ; ; ; ; ��{U���������W��     ��WU��UUUU��3333333333��UUUU��ff�������� ; ; ; ;��U{��? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U{�U3U�_�s�s�s�s�s�_�U�U���fÙ������� ; ; ; ;��U{��? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��    ����                ���������� ; ; ; ;��U{��? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��UUUUUU��UUUUUUUU                �� { { { {��U���? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��      ��        UUUUUUUUUUUUUUUU��U{U{U{U{������? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��UUUUUU��UUUUUUUU                ��U{U{U{U{������? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��      ��        UUUUUUUUUUUUUUUU��U{U{U{U{������? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��UUUUUU��UUUUUUUU                ��U;U;U;U;���{��? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��      ��        UUUUUUUUUUUUUUUU�� ; ; ; ;��U{��? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��UUUUUU��UUUUUUUU                �� ; ; ; ;��U{��? ; ; ; ; ��{U�� ? ; ; ; ;��U{��? ; ; ; ; ��{U��      ��        UUUUUUUUUUUUUUUU�� { { { {��U���? ; ; ; ; ��{U��  { { { {��U���? ; ; ; ; ��{U��UUUUUU��UUUUUUUU                ��UUUUUUUU������U{U{U{U{U{U{U_UUUUUUUUUUU������U{U{U{U{U������WWW����� � � � � � �  � �������/�?�?�?����������������U�U�U�U�U�U������U�U�U�U�U�������                / / / > > > < | � � � � � � ����������//??/?.?>?<�<�<�<<�>�>�>�.�/�� ^U^U^UWU������  տժժժ�����  _U^U^U^U������  �?�:�:�:���z��          ��UU��          ��UU��          ��UU��          ��UU��          ��UU��          ��UU��          ��UU��          ��UU��   � � � ���U���  �U�U�U�U�����  ��ժժժ�����  W�W�W�W�������  �������������� �UUUU_U�U]_���_��UUUUUUUUUU_U�_Z�UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�UUUUUUUUUUU��__�UUUUU�U��u_�u_zM��W5�5�5U��ըը�Zի�n��U���j��k�U}�W�U�U�U�U�W5��������������j�Cz=^�WUWUWUWU^ե��W���V����U諥z�]�^�^�_UW�W�T��U�U�USU�U5Uտ���Z����Z��Z����j����������}U���z�z�N�C�@�U��?��������j����z��V��Z����Z֪j��W�W�U�U�UUuU_UUUUUUUUUUUUUUUUU�j=�ճU=U�UUUUUU��j�j��:�:UOUMU��U�U��幕�U�WU��j������U~U�U��}�W}UWUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU�U�U�U�U�U�U�UU�������m�m�m���_�U�UzU�U�UUWUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������`���y����3�3���3�33���������������o�[�PPP[�o��� ����� ����� �����������������������<��������������0���0�������������������� �?�?�?�?�?�?���?�?�?�?�?�?�?��� ����� ����� ���������������������� �������������� �����������������������������������������<������������������������������?���?������������������������<��������?�?�?���?�?�?������������������������������������������������������������������������������������������������������������������٫�گ���������«�����]�������������]u�������������( ( ( ( ( ( ( ( ��������V��ƿ��ƿ��ƿ��ƿ��ƿ���V謹��������������UU  ����������������������������������������������������  UU����������( ����                    ����(           ����   ( ( ( ( ( ( ( (           � � (  ����            ������������   (�*�*����* * (       ����                * * ( ((((((((((((((((  UUUU                                         UUUU    UUUU    UUUU            UUUU    ����    ����  �?��S{������p�\��?�1�6�����ׯ7j>L��������^W:���[5n1~��߭ݻ=v� � � � ��� � � �  ? � �         � ���?�����?���        � � ��� � � � �   �� ?          ������������       @��G|�]U\��g�gY?�/Z=�u6Y�d�b�g�g���T]J|��W@�a�Y�V�6�uZ=�/? ����z�U�Al�k? ���9U���P���[[�E�U�i�n�� �i�T�A�Y��饺�/�
��[D'��תייә�?W�U�����������әәǙ��gD������������P�Q���������[�[�[��[����?��V��V��F�����[�[��[��������V�V��F������kkkkkkkU��@�@�@�@�@�@�U���\UuU�f��Tn��T��T��T��T��T��T��T��TՕ�T��T���TgՙtU]U������ff��UUUU��j�Y�fgY�UWUWQ�Un�U��WUUuћUk�Uk�Uk�Uk�Uk�UW��W�Uk�U5U]f�Uv�UkUUUUff��ff������U�U�eٙ�eک���WY����� �`�X���_w �AW�|WB|��U��AתՑ=�Ց=|FW|FW��Uw������=�թ=��Uתݪ����?�ժ��� �����d� ����W�W������ ��۪�e�e����?��WUWUW 0���0��U������������0�PC���������T���������?[�[�[�[�[�[�[U����?�����U�������U�U�����������������U�Uժ�����[U[�[�[�[�[�[���U�����?�������WUWU�?�����?WUWU������������T:P:T:P:T:P:T:P:  ������UUUUDD    DDUUUU������  ���������I�I�I�I ���{�;�{Իջ���������������������_�/�-�-{-{K����������������{K;;�{�A���:[?��������������  ��k5�:�?�? ������F��������V���V����z�����y���FFF�:f5f5f5�:����:��A�����F>FF���FFw�t��]������ FFFV���  ��k�k�k�k�k�k�kU��W�_����_�_�U�kUk�k�k�k�k�k���U�_�_����_�W��������U�����������������Uժ����������WUWW�W�����WWWWU������ ���W�WTGPAW��^���^՞ڝ�^����l�l�l���'b'b��_�����_���  ��'b'b��l�l�l���  ��_�����_�AGPTU�W��G ��^՞ڞ�]���^�����'b'b��l�l���p��_=��^�Տ���p���l�l���'b'b���ߟ�_�^���_��?���[�[����[U�����?{;{;����U���[U[U����߮ܮ����U�U����w�w;�?�?����f����,�� ���f����:�8�? �TUGUWU[[E[���E��D�Q�T�U��?��SQWEG�SdGF? 4?���ӱӴӵӱӓQgGASPT�����Ӵ�����u?�? ? ��������WU ��Ǫ��  ��UU  ������ǮǮǮ��ǺǺ����]u����C�S�����^���~�~�~�����V����@�H�@���!��Ǫ�� WU������������  UU��V V ����TjT���UU  �����jj�?U� ��Ӫ����F�F���Uש�����ӾӾӿӵӶӶӶ����v�����6�����ӵӿӿӼӼӽӿӪ���  UU��P�P������� �U��?jj���0 pU����   � U��ߠ����``� WU���� � ҁ��Ӫ�U����?�������������������������૪��������WU�����������U����?������?�?�?�?���  ��  ��  ��  ��  ��l��� ���<�<  �?P9�7 77<3<3���<� ��l����  3 7 7�7P9�?�     � �U��\UCC  ? ���N/??@\U���U � �  ??N/�/��?     �_�<క��p��  �/0<U]4\��\��\�\���  U54U54]55�?    ���d�Y�����  �7@7P77E7�7lUl}l�l�l}lU��  U5�6�6m5U5U9�     � 0 0 � � � �  ��3 0�?��� � �𨬪������  ���.�:�:�?�?    � l<�����=    ?�4<9C�d�  C��0d��L7��  � �/k3�1p�    0���0������ ��  ��0�6?7�<�<��� ����� �� �  �<�8�0� <       � p�0 �p           0 � \lU���� � �     ?Q0�5E;�� �    �?p�L�L*�8�0�      : � ���@   0 �      *�:�:�:@5�     ��<����������  ? /�?�?�?�?�?��������<�<�0�  �?�?�?�?<<    �<�Ǭ���]|   1 1?�?�6�?�?|�| �U�����<  �?�?�6�?:?1    �l9k�����k�l9���;��?�?����7�,4p��1 7�� � � � 3�1��<�pl8           � l              9  [ k � �        9 : >                 � � ��   ? ��R@P�V�� � � � �    �>��� ?      �����\flekV[k?��ߥ5U9P:P9D�P�E�kAlU\f\j���@�P�D�U9U5�6��?�l8l8l8,0,0,��,+�l8l8 � p � | �|���� ��3��=�?�<�Ӫ�>����� �    �� ? 1 1     � p � |�||����  : ? �=�û������ � � < < <���??3 3 < < <  ��s̮�?��=|���  : ? � �?���j � � L L p � ����:�?      � � | � ���~�� = 4 �/���ǽ޷��]�_>����� �    u3� ? 1 1     � � | ����>�=�� = 4 = ��>|�w��]�_� � � < < <u��:>3 3 < < <  � � |�����>�>~� = 4 = � ��>���] _ � L L p � �u���>�?      �����p�p������^  : 2 � � � � o o � ǀ��?��� ??��?? �      � ������������W  ; 2 � � � � ���^  3 �  � �� ?   � �      � ������������� ? � � ���5 \C[�[������  7 ; ? � ���   � � � ,  7 � ? �����>�3�� ���k��� � <    ��� � � �� ?� � � � �  7 � _? � ��~z�� [ � � p o �    ��� � 3 0    � � � ��07�� \? � ���~�� \ � � ǀ��?�  70����?׿;��   � � | � ��?�6�� = 4 �/��<�� �Q�S0�0�       4 < 1 1       � � | � �� ��  = 4 �#�38                                  �����w^�w]s��/? ���=p�t�zݸ��=\��� � � < <  �7?;\� �      � p � ��}���������?w� { { � � ��3�� �����<�� ?   � � |����L?L7� = 4 � ��<7pwp��~ � ��>� ]W�?0�8 ; � � � ������������� ? � � � � � u\\\�p������ ���?�?�
 ?     � � � <��70װ|? ����2�3�����������<     � � � � ��� ?����������������?������������������3������������������������������������������������?����������������� ���p���\�|�\�L3 �W_;�:�6�:�2\3l�\L��UpU��  �:�>�:�:U;U�   ���p���\�L����0 �W[;�:�>:>�0��\L
ܥpU��  :2�:�2Z;U�                                                                    ��pU�U\�L\�l3  �UU;�:�>�:�2\3L�\�|���p��� ��:�6�:�2W;W�   ��pUܥ\
L���0  �UZ;�:�>:>�0��\�L���p��� �:2�:�2[;W�                                                                   ��pU�U\�L\�l3  �UU;�:�6�:��\3|�\L��UpU��  ���6�:�2U;U�    ��pUܥ\
L���0  �UZ;�:�>:���0��\L
ܥpU��  ��2�:�2Z;U�                                                                    ��pU��\\���;  �U_;�:�:;;�;��\\��pU��  ;;�:�:_;U�    ��pUܥ\
L���;  �UZ;�:�>:2�;��\L
ܥpU��  :2�:�2Z;U�                                                                   � 0 ��\p_�_���� � :?������}>�ת�� � � � �    ��� ?     � p ��\p_�_���� � :5��?�ï�ת<� � � � � < <���?� > < <  ��3̾�_�_�_�~�� >����?���� � � � � � � ����?�        � \ \ \ ��/�?�� 5 5 ���3�3�0Ǫ׫��������  :� ? ?     � \ \ \���/�?�� 5 5 5 ���3�0ת>�<;0�0�0��< <�0? � ? > < <  � \ \�_ޟ�/�?�� 5 5 5 � ��3�0Ϫ�������0� � �>0�         ��W�U�W������  = 2 � � � >  � � � � ��?�� � �?3��?�        � W�U�U��������  9 6 � � � � ���^  ? � � � �� �?��?9      � W�U�U������ = � � � � � : �C��������  :  <  � � �� � p l ��<0�� s? �UU�?�7�7� � � ����      � � � � ��� ? � p ����7 � �? � UW���� � � � \ � �    ��� � ? ?    � p l ��;�� �? � UUV� �� � � � � � ��?�>0����?��3��  ��p�p-p��{�W{}{� 8 8 � ��>}�w�w��vGt\0�    ^��>�;%	@    ��p�p-p��[��pw�u 8 8����;�>w�w��]�^GT      V�T=�;�4      ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������L��LP�L��L��L��L��xآ��� � ���& �� �� �� �������� �!�2���  � � ��� �  �� u�� ��2� �3���  � � � � ����L�����e-e.ee���2����T���&  ��3��� � �; P�L����  ��3�����&   ��3�D�& �J�0����e<� �� �1�2���3�  �L7��� D�L7��� �L7��� ����$ƨ�3���& ��� ����ƨ�3���& � /��2��� �2Lv��ɉ��� �
��%��&��+)



e��i ��+JJJJe���-��. ��`� � �������������-���.� �� �ܩ ��`�i0���`� � � �* ����� ����`�  I����I�%��`���`�� ��`
 =�慦������'� ���)�������V��L����L�� ��`�������)������� ��`���"��)�� � �� U�����惥�)�� ��`��������)Ш������ ��`�����)�� R� �� U�ƆƁ����иƂд�����	��)�L0����� ��`�����)�� �� �� U�懥�i�����i ���@�����	��)�L0� ����� ��`�����)�� b� �� U�Ƈ��8�����ƂLl⥑�摥�)��� U�` ��`���L ���������(� � ������(��i0������`��)���)�
���L��L*� ��`����L��La� 	 >BFJNRVZ^bfj���#���$�������y�㨹��(���%�̅&� �/�(e/�+�#��$� ��#�#�/�/��)�ޥ#i|�#�$i�$��`� � ��iJJ���8�JJ�


ee���JJ�


ee���0���0� `� � ��8�JJ�L#� � ��8�JJ�


e���8�JJe���JJe���0���0� `� � ��iJJ�


e���8�JJe���JJe���0���0� `�� ��  � ��������`�敩 �����

iz� ��y�� ��y�����"�� ����!8龝�� �����!y����y��`H�H�H�2��� ��  �� ���2�5 �� �h�h�h(@���& ��� ��� � � �* ���  P����[��� �����5����& �5Ť���� �� z楢���쥣����5i<�5��`���Ơ`栥��>�]�:��8� g�i0���i ����������������i0�����i ����㥢���  祢�a�.�]�*�D g����ȑ���� ��i0��i ������� ���_��a�Ș �祢�a�����`�`���ơ`���K�]�G��8� g�i��i ��i0���i ����������������i0�����i ����㥣��� 祣�a�0�]�,�D g��ȱ����'��� ��i0��i ���ߩ�����a�����`�`



}�煥���i ���J��� g���e��i �������`� � ��@�� ��������`H)����hJJJJ�
ei@}��` 0`��� P���@p��      

�� ��� � �����`� �/ ����� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                  ��	��ȱ	�� �����0����J��� ����� �* ���`��� �y� �  �ޥ
����	���
`� ��� �������
����`
����	���
�
��	�ȱ	���� ���� ��L*� r�L*� R� 0]���JJJ���� ���Bȱ�3�

��3� �)�6� �� �!JJJJ�$�)pJJJJ	�0 	� � �`��-�>�����k�L���*��$8�'�$���)�* 	� ��`� �-�$ 	� ��`�*���'}$�$����)�* 	� ��`�-�� � 	� ��`�*�Ž$8�'�$��!)�$LA�!)�$���ǽ)�* 	� ��`�*� 	� ��`����)���0��)pJJJJ	�0�

��)�%�38��3��6� �3�6�3� �6� `�3e�3���6�6��ީ�6���3�ҥ�

��)�JJ$	J� `�����-`
ee������)�*�JJJJ�'��-`�����e`���ȱ������.�@���*��� �y� �  `��ý	��	��LR���ȱ��	�LR���ȱ�LR�
qe�����ȱ���LR�05

������� � ����)� � ���� � ��� � ���c��S)x�OJJ�����C��?�0&�8���
�� ���� � �� � Lt�e�������ܩ ���� � � �0

�������( ���) ����* ��	��� �* `f���_3y��1 o�z_� � �- \ ~ � / ��?��������Y�#���������o���X�\X�\�\��\�\��\����h��h�h.�h.h.�.��� �@  � �0   � �  � p� ���P XP �P \P �P �P 	h h@  h h0   	h h  	h ah  ��)�7���  ��  ��	��	��	��	@Tp � �  ��  ��	��	��	��	.@p �   	@T	}�	�� � �	��	��p �   �A� � � � � � � � � � � � � � � � � � � � X X � � X X X X � �  � 
� 
�x  
 
   ��3���
�
�
�
�XX �X�X�X 
�
�
�
�XX �X�X�X ����
�X ����
�X ����
�8 
� 
�X�X
�X   ��   E���A��� � � �  � �}  	�
\� � � �  � �}0  � � � }	T 	T T.0 � � �  }	T 	T T.@   �P� � � � � � � �  L � � � � � � � �x  � � � � � � � � � � � � � � � �  � � � � � � � � �x n � � � � � � � �   �����	h	@		h0�  ������
�(X�3�  ���2N��TT!T �� � �T�T!T ��!T   �� � � �  � � �  � � �  � �0   _���2��! 	  ! ! �!h��0 �0��@�!!h!@ 	@ @ !@�h� �@! 	  !!  �!h��0 � � �@�! �! 	 @ !}�h�   �"�  !�  #X  "<  "  !�  "�  "  "<  "�  #�  "  "<  #�  "�`   )��2�� �!� �!� ����}!@ }!h }!h }h���"� @ � @ � @�@�� � � � � � ����� � �! �! �h�!@ }!h }!h }�}h!@ � � � � ������ ��� �� � �@��� �  �  � � � � � � � � X < X "<  FX � #� X � �   � < � < � < � � X < X < � X � � X � X � X � X X � � � � � � �   ������� ��s���( ( ( ( X X X X 
 
 
 
 
< 
< 
< 
< 
� 
� 
� 
� 
� 
� 
� 
� 	� 	� 	� 	� 	� 	� 	� 	�   ��� � � � �8 �8 
�8 
�8 X8 �8 
8 
<8 	�8 	�8 	@8 	T8 	�8 	� 	� 	8 	8   �����@ 		@	T	@1  �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������H���