        0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l��� �փ����  =000000000000000000(00000  '(000��  (0000000	0000	000	0000	000	000	0000
0
0	000000
0
0	000000
0
0	00000000000                        �c%������  6''$%0''$%$0))&'0'&&$%"%$0$%$0'&&'0$%$'&$%0��  3$0$  $  $0 "  " !0! 
 ! 
 
"� 0 "  "  "!00! 
 ! 
 0 "  " !"!0"  "  ��ņ����  6� 0 � 0 0� 0  0 � 0 0� 0 � 0 0 0  0 � 0 0��  #00000	0
00
0000	0	00
00	0000000000	00	00
00	00	0
000
00	000
0	000���Ǉ���  :
'&0'00&00'&'00&+ 0 +0��  '!0
0!0$00#"
0������  :('���  ''&��� ���������  ��� ���b��/���� 2�� Z�o�Iw� z������� ��� ��L��`�������������_^FNNEzz#W4W2Yw� ��� V��Z���� ���
��� V��"���� ���L���(H� � Z� �z�����e����������C��������`e����h:м`��� ���Jjj(**HJ~�~�~�~�J~�~�~�~�hJ~�~�~�~�J~�~�~�~��ж����`            x   �   ?�  ��   ��   �� ��� ��?� ��� aÁ� aÃ� aÃ� Ã� �Ç� ���� ���� ���  ��  ��� ��� ���  ?�  �   �        �   �  �               � ��������  0�                   p   | |  | >  ><>  <><  80  ?0  ? g�� ����� � |p 0w� 8�����~s�  s�  � 8��������g   w   �   �  ��` /�p x<x |x|~ <x|g <y�g�s�c��`��`� � �?  �   �   �    @      ��]0` � ^��\�L����	 h� z�L��� q� ����}��]0 ����`�[)���������]�)��)��8�� �]`�\�������� ���])��]��])�`��])�	�]���]`��])�	�]���]�[)�\�)�`��]�)���)���])���
��])��]���]`�������]`�����`��]	�]���]�[)�`��]�)���)���])����
��]	�]���]`�������]`��])ߑ]`��]	 �]`��])��]	�]���]�[)�`��]�)��)��\���])�L���������`��])0��8�
��])�]���]`�i�����]`��])��]	�]���]�[)�`��]�)��)��\���])�L@��������`��])0�0��8�
��]	�]���]`�i�����]`��]0` L���])JJ�Y��])�V�����	��])�]`�\����L�������])�ީ f��� �]eYɗ�� �]`���
���� X�L�������	��]	�]`�\����L������])�ީ f��� �]8�Yɗ����]`���
���� X�L���])�Y��]�)�Z�����8�\���])��]��]�]`��])��]��])��]`���
���� X�Lh�� f����]eYɇ����]`�������]	�]`���
���� X�L�  f����]8�Yɟ�� �]��`         ������ ��� ��� �� �   � �]i�P��]i�Q�	�R�R
��Q}�}����P}
�}��� b��R���� B��R�`�)��XdY
&Y
&YeX��YFYjFYjFYj�XdY�JJJJ&WJ&WeX�FW&YFW&Y�Y�A=����JJ��JJ��JJ`�0��ɏӏݏ  �� !�   �()�34�   �mn�rs�   �op�tu�   �  �  �  ����]0� �\���[)��轷������Le��\�����[)�α�����Le���]�)

��k�ȱk���]�\�) )`JJJJJ��}�������]����])�� ��� �]�ȱ]��	���_L�� <Z�\��������])
���kȱ�l`�7����L��`��]0`�����&����������������������]��[)��L��)��Y�):0Y�] D�)�H)@��0	 h� z�L2� q� ��h)�L����]0L��`dY �X ��)$EX)<

�Y ��)	Y��]`�T�H�\�*
����P���Q��P� �]�U�P�Wȱ]�V�P�X ^��h:�`��n���m�V8�X�dm�X8�V����$m�\��n� 
�8`�\�8`�n�����Lˑ���8` 5�$m�\�L��n��
�����2��8`8`�PeQ�o��m��\��o���ee�e�ef�f� eg�g8`�$m�]LB��P�)@��)�LO���$m�]L\��P8`��R��S�T���W8�U�R�t�X8�V�S�m�V8�X�S�dL����U8�W�R�R�X8�V�S�K�V8�X�S�BL����X8�V�S�0�W8�U�R�)�U8�W�R� L钥V8�X�S��W8�U�R��U8�W�R�`8` �����]�`���)��[)���ک�\�� Xé���������]��]}�ɠ�
�� �]����]`�\�`� Xé���2�����]�
��hh`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      	                                                                      	                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   game6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       mx                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        b@�w0�                                                                      0xxx0 0 lll     ll�l�ll 0|�x�0  ��0f� 8l8v��v ``�     0```0 `00`  f<�<f   00�00       00`   �         00 0`�� |�����| 0p0000� x�8`�� x�8�x <l�� ����x 8`����x ��000 x��x��x x��|p  00  00  00  00`0`�`0   �  �  `00` x�0 0 |�����x 0x����� �ff|ff� <f���f< �lfffl� ~``x``~ ~``x``` <f���f> ������� x00000x ��x �flxlf� ``````~ ������� ������� 8l���l8 �ff|``� x����x �ff|lf� x��p�x �000000 ������� �����x0 ������� ��l88l� ���x00x �0`� x`````x �`0 xx 8l�           �00       x|�v �``|ff�   x���x |��v   x���x 8l`�``�   v��|��`lvff� 0 p000x  ��x�`flxl� p00000x   �����   �����   x���x   �ff|`�  v��|  �vf`�   |�x� 0|004   ����v   ���x0   ����l   �l8l�   ���|�  ��0d� 00�00   �0000� v�       8l��� �փ����  =000000000000000000(00000  '(000��  (0000000	0000	000	0000	000	000	0000
0
0	000000
0
0	000000
0
0	00000000000                        �c%������  6''$%0''$%$0))&'0'&&$%"%$0$%$0'&&'0$%$'&$%0��  3$0$  $  $0 "  " !0! 
 ! 
 
"� 0 "  "  "!00! 
 ! 
 0 "  " !"!0"  "  ��ņ����  6� 0 � 0 0� 0  0 � 0 0� 0 � 0 0 0  0 � 0 0��  #00000	0
00
0000	0	00
00	0000000000	00	00
00	00	0
000
00	000
0	000���Ǉ���  :
'&0'00&00'&'00&+ 0 +0��  '!0
0!0$00#"
0������  :('���  ''&��� ���������  ��� ���b��/���� 2�� Z�o�Iw� z������� ��� ��L��`�������������_^FNNEzz#W4W2Yw� ��� V��Z���� ���
��� V��"���� ���L���(H� � Z� �z�����e����������C��������`e����h:м`��� ���Jjj(**HJ~�~�~�~�J~�~�~�~�hJ~�~�~�~�J~�~�~�~��ж����`            x   �   ?�  ��   ��   �� ��� ��?� ��� aÁ� aÃ� aÃ� Ã� �Ç� ���� ���� ���  ��  ��� ��� ���  ?�  �   �        �   �  �               � ��������  0�                   p   | |  | >  ><>  <><  80  ?0  ? g�� ����� � |p 0w� 8�����~s�  s�  � 8��������g   w   �   �  ��` /�p x<x |x|~ <x|g <y�g�s�c��`��`� � �?  �   �   �    @      ��]0` � ^��\�L����	 h� z�L��� q� ����}��]0 ����`�[)���������]�)��)��8�� �]`�\�������� ���])��]��])�`��])�	�]���]`��])�	�]���]�[)�\�)�`��]�)���)���])���
��])��]���]`�������]`�����`��]	�]���]�[)�`��]�)���)���])����
��]	�]���]`�������]`��])ߑ]`��]	 �]`��])��]	�]���]�[)�`��]�)��)��\���])�L���������`��])0��8�
��])�]���]`�i�����]`��])��]	�]���]�[)�`��]�)��)��\���])�L@��������`��])0�0��8�
��]	�]���]`�i�����]`��]0` L���])JJ�Y��])�V�����	��])�]`�\����L�������])�ީ f��� �]eYɗ�� �]`���
���� X�L�������	��]	�]`�\����L������])�ީ f��� �]8�Yɗ����]`���
���� X�L���])�Y��]�)�Z�����8�\���])��]��]�]`��])��]��])��]`���
���� X�Lh�� f����]eYɇ����]`�������]	�]`���
���� X�L�  f����]8�Yɟ�� �]��`    �� ������ ��� ��� �� �   � �]i�P��]i�Q�	�R�R
��Q}�}����P}
�}��� b��R���� >��R�`�)��XdY
&Y
&YeX��YFYjFYjFYj�XdY�JJJJ&WJ&WeX�FW&YFW&Y�Y�A=����JJ��JJ��JJ`�0��ɏӏݏ  �� !�   �()�34�   �mn�rs�   �op�tu�   �  �  �  ����]0� �\���[)��轷������Le��\�����[)�α�����Le���]�)

��n�ȱn���]�\�) )`JJJJJ��}�������]����])�� ��� �]�ȱ]��	���_L�� <Z�\��ԅ�����])
���nȱ�o`�����L��`��]0`�����&����������������������]��[)��L��)��Y�):0Y�] D�)�H)@��0	 h� z�L2� q� ��h)�L����]0L��`dY �X ��)$EX)<

�Y ��)	Y��]`�T�H�\�*
�����P����Q��P� �]�U�P�Wȱ]�V�P�X Z��h:�`��q���p�V8�X�dp�X8�V��N��J$p�\��q�8`�\�8`�q�����L����8` 2� �$p�\�L��q��
�����2��8`$p
�\�!�q�
8`�q��\���ee�e� ef�f� eg�g`�$p�]L?��P�)@��)�LL���$p�]LY��P`��R��S�T���W8�U�R�t�X8�V�S�m�V8�X�S�dL����U8�W�R�R�X8�V�S�K�V8�X�S�BL����X8�V�S�0�W8�U�R�)�U8�W�R� L咥V8�X�S��W8�U�R��U8�W�R�`8` �����]�`���)��[)���ک�\�� Xé���������]��]}�ɠ�
�� �]����]`�\�`� Xé���2�����]�
��hh`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      	                                                                      	                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                   �&lib\sachen.obj >  t �`4�&��&��&`�&��&4�&��& 8��     ���&L�&lib\sv.obj u � ~�|�&|�&��&��&��&��&��&  9��    Ÿ��&��&game6.obj >�  t
 <2��& �&�& �'�&D�&��& �Y[d    2�@�&��&move.obj <2 � 2���&  �'$ �'� �'\�&d �'��& �Oe    �k��&�&defind.obj � � �AH�&� �'� �'�'��&� �'��& toU:    u[��&\�&game6.lnk ~ �؋ ����&��&��&    ��&    ��&  N)�    ���&�
�&        ��v �&��&stage_1.obj  &�  ����&$�'(�'��'<�&h�'��& �."�    �vd�&��&stage_2.obj  J�~ Dt(�&��'��'�'��&��'��& �2Y)    v���&<�&stage_3.obj  �u �ll�&4�'8�'��'��&x�'��& 1�V)    P��&��&stage_4.obj  ۋF -	 ��&��'��'(�'�& �'��& ��)�    � 0�&��&stage_5.obj   u � ��&D�'H�'��'L�&��'��& �&�    >�t�&�&stage_6.obj  ,  a�8�&��'��'8�'��&�'��& ��)�    ���&L�&stage_7.obj   u ��|�&T�'X�'��'��&��'��& @�)�    [���&��&stage_8.obj  ~�W u���&��'��'H�'�& �'��& �)�    =@�&��&stage_9.obj  �� ��E�&d�'h�'��'`�&��'��& &�    �1��&�&stage_10.obj v� �� ���H�&��'��'`�'��&8�'��& *�)�    !���&`�&stage_11.obj �  �W� ����&��'��'��'��&��'��& �6U:    �1	�&��&stage_12.obj  u �~� u+��&�'�'��'8	�&X�'��& ��)�    ��`	�&��&stage_13.obj �� t�   	�&��'��'�'�	�&��'��& �*�    �6�	�&8	�&stage_14.obj [�� ��$ F�h	�&0�'4�'��'�	�&x�'��& ��)�    �&�	�&�	�&stage_15.obj �� 6�	 <4��	�&��'��'0	�'
�&	�'��& [�)�    �	8
�&�	�&stage_16.obj .�1 �� �	��	�&P	�'T	�'�	�'�
�&�	�'��& ��)�    ��    
�&LK @GAME6.LNK �	        @
�&    lib\io.obj 	 U� [�lib\io.asm  5i[ P�6t
�&�
�&�
�&    (�&    �
�& P[Vd    �{
�&��&        ���
    �
�&AS LIB\IO.ASM -OLIB\IO.OBJ Q        �
�&    lib\screen.obj   �� u�lib\screen.asm   �~  t	�& �&$�&    ��&    �
�& �~�    ��    (�&AS LIB\SCREEN.ASM -OLIB\SCREEN.OBJ �        X�&    lib\num.obj  �$P F�Plib\num.asm  P�� �1[��&��&��&    D�&    �
�& @�pc    ~    ��&AS LIB\NUM.ASM -OLIB\NUM.OBJ  u'        ��&    lib\mustbl.obj � �� �[+lib\mustbl.asm �  � P�,�&<�&@�&    ��&    �
�& s��    '     D�&AS LIB\MUSTBL.ASM -OLIB\MUSTBL.OBJ         t�&    lib\music.obj *   �  P�lib\music.asm �� �PQ N�Q��&��&��&    t�&    �
�& ��Y5    �F    ��&AS LIB\MUSIC.ASM -OLIB\MUSIC.OBJ �        �&    lib\checksum.obj [�> %c~ �*lib\checksum.asm *%  � �X�&l�&p�&    �&    �
�& [:��    P�    t�&AS LIB\CHECKSUM.ASM -OLIB\CHECKSUM.OBJ �        ��&    lib\sachen.obj � �5u � lib\sachen.asm � � @�F��&�&�&    ��&    �
�& rʺ�    ��    �&AS LIB\SACHEN.ASM -OLIB\SACHEN.OBJ �        <�&    lib\sv.obj   	�v �|�lib\sv.asm ^ �]� �샄�&��&��&    �&    �
�& ,(��    �    ��&AS LIB\SV.ASM -OLIB\SV.OBJ         ��&    game6.obj q� � �[�game6.asm �^ �� ���&�&�&    `�&    �
�& �V[d    厜�&�&g6_bgd.pxl G & �vL�&X�&\�&    ��&    ��& %�#�    F�S�&            �F�&��&`�&g6_spr.pxl 1 [�v �6,��&��&��&    < �'    ��& �P��    %�    ��&AS GAME6.ASM -OGAME6.OBJ &�&�W�+����]�&        ��&    move.obj �F ��u +��move.asm �F =�� �F( �'4 �'8 �'    � �'    �
�& �Oe    &�    < �'AS MOVE.ASM -OMOVE.OBJ t        l �'    defind.obj � ��V �^�defind.asm � �F �V�� �'� �'� �'    @�'    �
�& FlU:    �&    � �'AS DEFIND.ASM -ODEFIND.OBJ �        � �'    stage_1.obj  �V ,%stage_1.asm  �^� �&,�'8�'<�'    ��'    �
�& &%"�     R    @�'AS STAGE_1.ASM -OSTAGE_1.OBJ F�         p�'    stage_2.obj  ��t �}�stage_2.asm    �  ���'��'��'    P�'    �
�& �0X)    ,    ��'AS STAGE_2.ASM -OSTAGE_2.OBJ �[        ��'    stage_3.obj  7P� ��1stage_3.asm  1[[ �}6<�'H�'L�'    ��'    �
�& QV)    F�    P�'AS STAGE_3.ASM -OSTAGE_3.OBJ ^�&        ��'    stage_4.obj  ��F �F�stage_4.asm  �F� F�@��'��'��'    `�'    �
�& ��%�    F�    ��'AS STAGE_4.ASM -OSTAGE_4.OBJ ��        �'    stage_5.obj  ,% �&stage_5.asm  �� ,%L�'X�'\�'    ��'    �
�& ���    ��    `�'AS STAGE_5.ASM -OSTAGE_5.OBJ �        ��'    stage_6.obj  ��1 ��stage_6.asm  ��v �|���'��'��'    p�'    �
�& &�    F�    ��'AS STAGE_6.ASM -OSTAGE_6.OBJ ��        �'    stage_7.obj  ~�2 �Fstage_7.asm  F£ %�6\�'h�'l�'    ��'    �
�& %t&�    �    p�'AS STAGE_7.ASM -OSTAGE_7.OBJ tu�        ��'    stage_8.obj  �& W�stage_8.asm  �H �x
��'��'��'    ��'    �
�& ��&�    t    ��'AS STAGE_8.ASM -OSTAGE_8.OBJ *%^        (�'    stage_9.obj  � ��stage_9.asm  �px 1[[l�'x�'|�'    �'    �
�& �X$�    t&    ��'AS STAGE_9.ASM -OSTAGE_9.OBJ t        ��'    stage_10.obj �� ��W  �stage_10.asm ��& X& ? t��'�'�'    ��� � � ��� � � � �)��� ũ)����� � ������i��i ���� ���e � ���������	 ť )��������)�S����L������������� ��������� ������i ���Lƀ@@@@@@8  0@P`8@@@@@@p�����Т �*�	�,8��,�����p��*�	�,i�,���������i����ɀ�L]�d � ɴ�
������`

��h��*�i��.�j��2�k��6���)�-i�1�5���,�4i�0�8� �+�/�3�7`	
+,)*78'(56%&34#$12!"/0 -.                     � �              �     D3�L0�L3@� 1DD33DD            � 1@L�03D1���1 D 1��0�1� 1  � 1�@  D 1� 1� 1�D13@���3 D3��03��13�L13D3�3D    D 1�13��13��13@D 3@L 3@L3�L33 �  �           �          �  @    ��L 3�1�1� ��0� 1� 1� �1���� 1� 0�L3@�   �0�3L  �D1� 1� 1� ������13�L13��13���    D3���13��1� 1� �L33�L33�L03�L          ��           �    @�03�03�� 3 ��L           @  � 3��L���� @�3�L0� 1�  L 3�0�  � 1� 1� 1������ @�03��13�L13���3�    D�1�L13��13�� @L 3@L3DL3�L     �   �        �          0 �      DD13DD3 � 3�0�3D 03�D1� 1� 1D 3���@1� 1�0�� 1 D  @�1�   1� 1� 1� 1D ���@13��13�L13��13DD3D    �3D13��1�@1� 1D 33�L33�L13�L3@D� ��@���������`�����[������d ��� ������ �� Y������������ i<� ��`

�� ���� � �����`� �/ ������`������@�]�<��8�� �ĥi0��i �������������i0���i ��������  	����a�1�]�-�D �Ģ���ȑ�� ��� ��i0��i ���ߩ��� ���_��a�Ș �����a�����`��`�����`���M�]�I��8�� �ĥi��i ��i0��i �������������i0���i �������� 	����a�1�]�-�D �Ģ�ȱ����'��� ��i0��i ���ߩ�����a�����`��`



}:���;�i ��J��� �Ĺ>�e��i ������`@�@� ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�  ������ ��??�  ������ ��??�  ����� ��??�                  ?������� ?   ?��������?�?   ?����������?   ?���? ����?   ?���? ����?   ?���? ����??   ?���������??   ?����������?   ?���������?   ?�� ������?   ?�� ������?�� ��� ������?�� ������������?�� ���������?��?�� �?������� ?��                 ������?��?��  ���������?��  ���������?��  ? �����  ?�  ? �����  ?�  ? �����  ?�  ��������??�  ���������?��  ���������?��   �����?�  ��   ���� �  ?�   ���� �  ?�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   P @ C |  �
U�UUUW�   ���
�
�
W*�    Z X P P P�� _  �eUU U � %    h������������*�
 � ��
�
�*�**     ` � � � � �     	 	 & � �        � � T �      � ����
�
         @ P        ��
�
�
�*�*    ��
�
�
�
�*��0��� � � � �    � 0  
 � �     � � � � �� �       
 �         � � @ ��*�*�*j*Z�W�         
�&�* O������j�W�S�    �
�&�&�*�*�O������[�W�S���)�&�����*�*�O�*�*�*V�R�B� � �@�@  �      �
�*i*j)ZT0  � �@�@        �
�*i*i)jZ=
0(                 �`	X	X
�
�
�
�
����  ������  ���
�
�
�
�
�
�
�
U�U�������������� XX� \_T

��W��?�������9����n�l:n�n��?Wիꏪ����vն��������������W�������       @@DD          U  @  T      U   T  @                                                        	
    !"#$%&'()* +,-./0123456789:;<= >?@ABCDEFGHIJKLMNO   PQRSTUVWXYZ[\] ^_     `abcdefghijk         lmnopqrstuv          w  xR   yz                                                                                                                                                                                                                       �            ��UU            �U	             ��V            � U*              ��     ��Z�U�UXUXU `�ZVUUUUUUU D UUUUUUUUUU@    U%UUUUUUUU T P  `UYUUUUUUUUUUTU%U�UUUUUUUUPU A � ZViUUUUUUUUUUUUUUUUUA    
  U�UUUUUUQU T    *�VUUUUUUU            � �            �U?   �@U@U@U@U U  �Z�UUUUUUUU @��UUUUUUUUUUUU@ 	 �
U%UUUUUUUU            	 XUVUTUVVVVV      � ������� � ���������� * * �
�*����������P        ����      �*�*������TP          �  �*�����*�*�
�
 @      �
�
�
�*TP             _�W�U|U\U_UWUWUU�U�UUUPUPU UU  ��_�U�V�V�Z�Z  ? �UU=U��U     � � � ���    ������      ���������*PU@U@UUU U U U	 	 	 	 	  % % VVVVTU`U�U�U������ � � ���
 
 * * �������������*�
�������� � � �������*�*���������
��������
�
�
�*�*�*���� � * * 
 
 �*�*������������ � � � � � ���WU�U�U�U�V�V�V�ZUUUUUUUUUUUUU�kPkPkUkUk�k�Z�ZPUPUPU@UUUUUU����������*�*�
��
�
�����������*�
�
��� � *  U U@U@UPUTUT�U�% % 	 	 	      U V V X P �    �� U U UVV�����*�*��������� � � � ������**�*�*�������� ������*� � � �  �����������
�
� �
����������    ��*�
��� � �  ���������
�    �j^�~���W _ � �UUUUjU�Z��U�U?��V�V�V�V�Z��_�|�UUUUUUUUUUVժ�j=�
��� �      ����������      * 
@
@@P T U UU�U%U	U	UU� ) X              ������ �       �� 
           �              �           �����
        � ��
�        
 
 
 
               ��              
           �����*( �        � � ��U�_ � � �� � * U�?  
    ���            * � @U              	                  � � � �      �����������������������**    �*�*�� � � ��*�
 
 *�*�*�*���������������� * 
 � ��
�*�*�
�   �*�*�*�*�������� � � � �
�������*�����*�
�
(
 
 �������
�
�
�
�*��
           �� � � � � � � ���������*�
������*�� � � � �����������������
�
�
�* � �������
�*�*�*�*�*�*�
���
�
����  ���� � � � � �  
 
 
       �*�*�*�*�*������               �
�*�
�         ������          ���*                           J���؎	 M� 2� Kɩ � �   � 0�  ����& �
� �)��� � 2��� ��څ������ׅ�:��ͅ��`dZ���̍���h�<�idedfdgd ddd\��� L� \� � >� �� Q� 4��� ]��[ � � �� � �� � � �� � �� � �� �� ��\�\��� ŭ��ίd\L��``����������� ���� ������	���!��������
���"�����������������&�'`�Z
�Y���������� ��a:�XȄVdW�Wi�W����P���Q�V�


� �P�V�V�8�


��P����P���P�V�X��Y��)�	�����


�����8�


��`������������������]��[-�	��])�]`��]�])���])��	�����]`�\
��
m�_���]���^` 	 �c�A��dPdQ�Z
��<��=��P���.����� �6�S�P)��SS��SS��SS�Q�AS�A�P���P)��Q�Q�dб`PRESS START BUTTON Copyright 1991,1992�  Thin Chen Enter.����������� �é �� ]ɩ�������� ����������� ��� ��� �� ���� K�L2�d��������4�ĜT��t����$���D�Ԫ�Z
��<悔=滛L��SCORE �STAGE �� �)��� � 2���� ���	��s��� ���Z �Ǫ)��JJJJ ���L�� ��j �hi��j���j�i�h�hdi��;�i��� � V��h �� ���: ���i ��L���[)�`�[)�`��� ��l��� ��d(�g�'�f�&�e�% �ǥ0 ���/ ���. ���-L���e � �� z��P�����`�� �� å )��P��L\���� �ǩ�� � V��`L��`���`�����`�`L�� ��Z
� ����������`GAME OVER��颇 ]ɢ �)��� � 2����	��ͅ��� ���<e � ����P�� å )��P����L$�GAME CPMPLETE !�You have defiance�all SIXTEEN STAGEs.�CAN`T BELIEVE you�DID IT, But you�just did it !!!!!�In the last�We appreciate to�buy BALLOON FIGHT�that`s has great�meaning to our�company. So,�THANK YOU AGAIN !� �   PRESS ANY KEY���!	��`���� ]� ���e � �� Kɢ �)��� ũ�������� �� ����e � ������ V��i �� ���  ���X ���  ���  ���2 ���0 ���0 ���  ���= ���  ��L�� 2�����Z���ZLm���e � ����� ]ɩ����&��� ���xe � ��� ��L$�TIMES = ����	�[)�ΰ��` �ȭ������e � ��L(ɜ)�,�/�2�5�8�;�>���+�.�1�4�7�:�=�@�Z
�����b����c� �b�'�(`,'�`�(��'�(� �(��iL��d��*� �¨)�* � �)�� ��)�*`
 ,'�`dV�d�)�+��+��V��(��iL��b�


i�Rȱb�


i�Sȱb�U��d�)��Z�V����H� �)��� �h ��h��L[�X��Y�Y���P���Q��P d��Y�Y�`��P)�P`��P)�P�X����Pi�T8�S��S8�T��0`�� �Pi�T8�R��R8�T��`��	��P�S�
`��P�S�`��P	��P�X�5��"��� �P�R�`i�P`� �P�R�`8��P`��P�S�`i�P`��P�S�`8�ɟ�� �P`����'�3�?�K�W�u�a��k��������������G�e�Q�o�[�y���������������"#� ��"#� ��"#� ��#"�@��#"�@��#"�@
��"#� ��"#� 	��"#� 
��#"�@��#"�@	��#"�@,-�78�FG� ,-�9:�HI� ./�;<�JK� -,�87�GF�@-,�:9�IH�@/.�<;�KJ�@12�>?�FG� 12�@A�HI� 12�BC�JK� 21�?>�GF�@21�A@�IH�@21�CB�KJ�@�ij�\]� �ef�bc� ,-�kl�bc� �ji�]\�@�fe�cb�@-,�lk�cb�@
�VW�bc� �QR�\]� N	�XY�dc� 
�WV�cb�@�RQ�]\�@	N�YX�cd�@�ef�bc� �gh�^q� �eh�`a� �fe�cb�@�hg�q^�@�he�a`�@�QR�\]� �QS�^_� �TU�`a� �RQ�]\�@�SQ�_^�@�UT�a`�@?�?�K�W�c�m�c�m�c�m�w�����������������������  �������   �������@vw�|}���� xy������� z{������� wv�}|����@yx�������@{z�������@vw�|}���� vw�~���� vw������ wv�}|����@wv�~����@wv������@���$�-�6�?�J�U�`�m�z���������										
	
		

	
	

		

					

����� �'�4�A�B�I�P�Z�[�k�~� 	  
   	   	
	   	
  		 		 �}|����@yx�������@{z�������@vw�|}���� vw�~���� vw������ wv�}|����@wv�~����@wv������@���$�-�6�?�J�U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                @vw�|}���� vw�~���� vw������ wv�}|����@wv�~����@wv������@���$�-�6�?�J�U  �  �`�m�z���������										
	
		

	
	

		

					

����� �'�4�A�B�I�P�Z�[�k�  �  �~� 	  
   	   	
	   	
  		 		 �ύ& L�����1ͩ��  � � � � � � � � � � � ��" ��d`� ��@����'� ����0e�� e����`�


 n��
e�� e�`d
&
&
&
&��
&e��e��@e�`H� ��hHJJJJ ��h)	0�:���H�Z�Z�Z ��z�z�z�h`8� d
&
&
&i ���e�� Z�� ��� �� ��0e�� e�z����8��~����`����������N�N*N*L9�N*N*N�N*N*LQ�N*N*N�N*N*Li�N*N*N�N*N*L��N*N*` �U�L��� V�� ��������������� ��L��`

����� ���6����C����,0)�*��,��)��+����i�nL��ȩ �)�*�+�,L�����e�nL������������  I�� �
>��`�H�H�H�H� �� � � � � � � � � 	� 
� � � � � � � � � � � � � � � � � � � � � �Сh�h�h�h�`��e�E����&E�m `��L������ ����������� ���L�­�`��� �	� �� ���`�	�+� �
� �����
m�
��� � � � �	`
�
m�� �sÙ
������	`@:� 8� 8�6�06�.�<$p8v�8 :� ���)����� �������i��i ��i��i ���ة)������ � )�����ɨ��`�Z��J�"�JJ����e"�#���i �$�H� �#hz��#�$�



e��i ��JJJJe�� �ĥm��� ��ȱ��i�� e��i0��i ���� �Ĭ$�#`�����0�� iɪ�骍�`H)���ąhJJJJ�
ei@}�ą` 0`��� P���@p��      )AYq�����1Iay������@ � � �Z�	�)��
�*���+���,�L�)
��	�%�
�&��'��(Z ��z�)�	�*�
�+��,��+)*� ��z������Љ`�)�%�*�&�+�'�,�(�')i��')Ji� �0� d!�%�'m:H���!E � h �ĭ(JJe��i ��&�



e��i ��'J�jJJJe��()�#� � �,'p�����0�� �ڪ�������#�!........��߬ �Q����e ��e!��m ��i ���L�` @��P�� `��0p��D��T��$d��4t��H��X��(h��8x��L��\��,l��<|��A��Q��!a��1q��E��U��%e��5u��	I��Y��)i��9y��M��]��-m��=}��B��R��"b��2r��F��V��&f��6v��
J��Z��*j��:z��N��^��.n��>~��C��S��#c��3s��G��W��'g��7w��K��[��+k��;{��O��_��/o��?��H��
���


�h ĭ���`��8��
��i
�%�



%`�|�%�ȥ&�ȥ'�ȥ(�Ȑ�(�%�ȅ%�&�ȅ&�'�ȅ'8&-&.&/&0�����`            
      (   P   d   �   �     �  �  �  @  '   N  @�  �8 �� @ �  5 @B ��  	=  z ���  -1 Zb ��Hژ��?
�h�3h�2`�N�O� �NH
���ȍ���ȍ�� ����G`l������Ȣ �N� �����`� �N� �����`� �N�( ��������N`� �1�Y� �1��)�� �+��� �+��"�� � � �( ����`d1 ɢ!���+���(�Y�1��` cɥ1��`�t1���-�+��Lɜ+�:�;� � �:�2��������?� �<�G�,��B�C�D�1`�1�`�B��L�����C��C�`� �B�Dm+�C�?�
�<�	�<�� L�˽̪�2�8�3�9�B� �80LN����LQ����Lj����� �?����� ̱8�Dm+�C �L����� ̱8�K�88�K�8�9� �9L�����Lq�����,�,�,}̨�/�8�0�9 �L�����- ̱8H ̱8H�,}̨�8�/�9�0�,�,h�9h�8L�����' ̤B�̠ �8�M������8i�8� e9�9�BL����� ̱8Hȱ8�9h�8L�����2�̹O)��O:�O� �P� ��8���̦B�<L�� � �L������B��)��O)�O�O�O ̦BL��ɀ�(逼�

���̙M��̙N��̙O��̙P ̦BL�ɤB�G��̨�H̝ �|̝ �O� �P�  ̠ �8���̦B�< ̥B
��8�2�9�3�B��G��G��`�A��>��>�L�ˠ �6���� �AL����� ̱6�W�68�W�6�7� �7L��

� ̱6���̅> ̽�̍( ��̍) ���)�* 	�* L��   �8��9`�6��7`H���K
�LhJH��mL�LhnLnK��L�K`X���<�Ĭ}T@��־���pk_UPG?8(�\��h.�ʴ��xeZKC< 3m.                                   t   q  
  ?<�� �P  а� �@� �� �p� Ё� ��� ��  �@� � � ��  ��� �P   xH�Z� ��  � '� �ɭ E��e��E*�z�hX@x,$ ,% X@�������������������� ? ?   ? ����������� ������ � ? ? � � �����0�0� � � ����?���� � ����� �0����� � ����� � � � � � �?� 0� �    ��� � � �    ���?� 0� �   � � � �    � �� � � �    � �?�         � � � �     � ����������� � �0����������������? � � �� � ��� �������������������<�� � ��� �������������������<�� � ���  � ����������������<�� � � � ���������������� ?����� � ���  � ������������  ?�� ? ? ?3?  �������������� �������������� ?����� � � �  ��������������   ? � ? ? ���� � � ��� � �����? ?   ? ? ?���� � � � � ����� ? ? ? ? ? ��?��� � � � � ����      <��������������������������� �0� ����������������� ? �     ���������������������?�?���?�?� � � �    � ��������?�?���?��� � � �    ��� � ���� � � ��� ? ?   ? ? �� ����    ��   <  ? ������ � � � � �����? � ���� � �3� ���������������������??   ?  ��?�?����������?��?   �   � ��<����������?����?   �  � � ����������� � ���0���������� �???   ?  � ��?���������� �3?   �   � ��<���������� ���?   �  � � �?���������� ?  �  ? �������� � � �������        ��?�� �������������      �?�������������������     ? ?<������������������ � ? ? ?  � ?����� � � � ����?�  0 � �   ���� � �0   ? ���������� � � � ?������� � �  �������������� �������������� ?������� � � ��������������  ?����� � � ��������������  ?����� ��  � ������������� �������������������������������� ������ � � � � � ������� ����� �� � � � � � ������ � ������ � � � � � � ���� � ����� ���� � � � � ������ � ����� �����?��� � ��������������������?��� � � �������������������?��� � �  � ����������������������� � � � �����������������?�?�?�?�?�������� � � ����������?� ���� ��� � � � � �   � � �����? 3  �������� ��� � ��?�����? 3  � ��������� � � ��������������������������������������������� ? ?   ? ���������� � ����?���� � ���� � � � � � � ������������������������������������?�� ?0 � �������������� ����?�� ? � ? � ��?�� ? ������������� ���?���?�� ?  ������������ ��������������������������������������?�<��� �   � � � � ��� � � � � � � ���� ����?� �� � � � � � ������?       ��� � � � � �0���������� � � ������������� � ��������?���?������ � �� � � ����������?���������� �� � ������� �0� � ���?�?�???�<�� � ������?������� ��?�����?�?�� �  ������������ ����������?�?�?���� �    ��������������?�?��0        ��������?�����?0         ����?���   ��?0� � �   < ������ ? ?��?������ � � � � ������� �? �?�������� � � � � � �����                   T U@U@UPUPU@U      Q U   P T U U@U@U U U  Q E EUU U    @ P T T U U T   U EUU  U U UUU U @PUTETUUUTUTU  TYYeeQYUY  @PUTETUUUTUTUVYYQeUeYTVYYeQeUYY@PUTUTUUUUUTUTUTUUUUUUUUU        \ V u E      0  %   @U U W \ U �  �  1  %     T P � \ U �  �  0  %     T P C \ U �  �UU 5  %     T P A T U U U U        PU@  \ U �  �VUx %    TUPU� W@U@w@D@wYT,  	    VT8  %    PU@  T U U U UUT      �u�W�� W�W�W  �/�� 5 � � <  �W���U`�@U�W��5 � � � � � ? �  U@U@U@U@U@U @ U U U U U  T �U��|�X�PU�����  ? ? 7 = ?  ?         \ v E u      0  '    U@UPPUTUTUPUPU                @ @ P P @  TUUUUQUUU     @ @ P P @ @TUUUUQUUUU  Y e$��ee T U@U@UPUPU@U@U e��QUR�U� U�W���U�W�W   ��� �� <  @U U # T U w D w   0  %     @  0 ��PU�]Q�]UUW  " 	    @0 ��PU�]Q�]P�UWT� ! 	       0�@uPUpW@TpWUT� � " 	   YV, � %     U T0 ��PU�]Q�]eYW� " 	    U0H��PU�]Q�]P�e[T� ! 	    U T��@uPUpW@TpWeYP� " 	    U���U U�U�_   = ? � � � %     P���P����_@U�C� /  = = = 1   ��\�V�TY\�?� �           P���^�PuU�U0� �? �        w W���_�W�W W�7 = � � � �5 � @PUTUTEUUUUTU  \ V u E�u�W��0  %   �/�� PU@  # T U U ]VT    % ,VT  ,  %   PU@  # T U ] QVT    %   TUPU@  T U ] QYT    %  ,TUPU@  T ] Q ]VUT,  %  , W              5                Q ] � p P � � ����UUU     Q � | T T t � <� ��/� � � 5    ] U � p P � � �� � ���UW/   ] U � T T t � <=��� � � 5    U U � T T t � < T P � � T U ] Q      %  , T P � � T U U ]      %    T P @ � T U U ]UU    % ,       0 T U ] QUUT,  %  ,    @ @ � � @ T    ��
�
�
�
�     �  �`0QpU    � ����� � ���� � � 5   @ULW�U � �      � ) � �Q@    @ULW�U U T      )
�%eU         � � � ����� � �
 * � � ��� �    � �����������   
 ) & � � *  � � � � � � � �* � �jj
�
�� � �  �����T��V*      �� � � @ � �@�P� Z* 
    
 
 * �  � � @ � �@�P� Z�� � � @ � �@�P�* 
     
h
� � �   @ � �@�P�� *     
h
� V T T T P�� _  eUUUU � %    X P P P @ C |  �
U�UUUW�   ���
�
�
W*�    Z X P P P�� _  �eUU U � %    h������������*�
 � ��
�
�*�**     ` � � � � �     	 	 & � �        � � T �      � ����
�
         @ P        ��
�
�
�*�*    ��
�
�
�
�*��0��� � � � �    � 0  
 � �     � � � � �� �       
 �         � � @ ��*�*�*j*Z�W�         
�&�* O������j�W�S�    �
�&�&�*�*�O������[�W�S���)�&�����*�*�O�*�*�*V�R�B� � �@�@  �      �
�*i*j)ZT0  � �@�@        �
�*i*i)jZ=
0(                 �`	X	X
�
�
�
�
����  ������  ���
�
�
�
�
�
�
�
U�U�������������� XX� \_T

��W��?�������9����n�l:n�n��?Wիꏪ����vն��������������W�������       @@DD          U  @  T      U   T  @                                                        	
    !"#$%&'()* +,-./0123456789:;<= >?@ABCDEFGHIJKLMNO   PQRSTUVWXYZ[\] ^_     `abcdefghijk         lmnopqrstuv          w  xR   yz                                                                                                                                                                                                                       �            ��UU            �U	             ��V            � U*              ��     ��Z�U�UXUXU `�ZVUUUUUUU D UUUUUUUUUU@    U%UUUUUUUU T P  `UYUUUUUUUUUUTU%U�UUUUUUUUPU A � ZViUUUUUUUUUUUUUUUUUA    
  U�UUUUUUQU T    *�VUUUUUUU            � �            �U?   �@U@U@U@U U  �Z�UUUUUUUU @��UUUUUUUUUUUU@ 	 �
U%UUUUUUUU            	 XUVUTUVVVVV      � ������� � ���������� * * �
�*����������P        ����      �*�*������TP          �  �*�����*�*�
�
 @      �
�
�
�*TP             _�W�U|U\U_UWUWUU�U�UUUPUPU UU  ��_�U�V�V�Z�Z  ? �UU=U��U     � � � ���    ������      ���������*PU@U@UUU U U U	 	 	 	 	  % % VVVVTU`U�U�U������ � � ���
 
 * * �������������*�
�������� � � �������*�*���������
��������
�
�
�*�*�*���� � * * 
 
 �*�*������������ � � � � � ���WU�U�U�U�V�V�V�ZUUUUUUUUUUUUU�kPkPkUkUk�k�Z�ZPUPUPU@UUUUUU����������*�*�
��
�
�����������*�
�
��� � *  U U@U@UPUTUT�U�% % 	 	 	      U V V X P �    �� U U UVV�����*�*��������� � � � ������**�*�*�������� ������*� � � �  �����������
�
� �
����������    ��*�
��� � �  ���������
�    �j^�~���W _ � �UUUUjU�Z��U�U?��V�V�V�V�Z��_�|�UUUUUUUUUUVժ�j=�
��� �      ����������      * 
@
@@P T U UU�U%U	U	UU� ) X              ������ �       �� 
           �              �           �����
        � ��
�        
 
 
 
               ��              
           �����*( �        � � ��U�_ � � �� � * U�?  
    ���            * � @U              	                  � � � �      �����������������������**    �*�*�� � � ��*�
 
 *�*�*�*���������������� * 
 � ��
�*�*�
�   �*�*�*�*�������� � � � �
�������*�����*�
�
(
 
 �������
�
�
�
�*��
           �� � � � � � � ���������*�
������*�� � � � �����������������
�
�
�* � �������
�*�*�*�*�*�*�
���
�
����  ���� � � � � �  
 
 
       �*�*�*�*�*������               �
�*�
�         ������          ���*                           P���؎	 M� 2� Qɩ � �   � 0�  ����& �
� �)��� � 2��� ����������ׅ�@��ͅ��`dZ���̍�dedfdgd ddd\��� R� b� �� D� �� W� ���� c��[ � � �� �� �� -� 4� |� � �� � �� � ��\�\��� ŭ��ίd\L��``������k�;�l������� ���� ������	���!��������
���"�����������������&�'`�Z
�Y���������� ��a:�XȄVdW�Wi�W�����P����Q�V�


� �P�V�V�8�


��P����P���P�V�X��Y��)�	���x�


���y�8�


��`������������������]��[-�	��])�]`��]�])���])��	�����]`�\
��
m�_����]����^` 	 �c�A��dPdQ�Z
��B��C��P���4����� �<�S�P)��SS��SS��SS�Q�AS�A�P���P)��Q�Q�dб`PRESS START BUTTON Copyright 1991,1992�  Thin Chen Enter.�� ������� �é �� cɩ�������� ����������� ��� ��� �� ���� Q�L2�`�𔀖���0���P���p� ��� ���@�Ъ�Z
��B悔C滛L��SCORE �STAGE �� �)��� � 2���� ���	��y��� ���Z �Ǫ)��JJJJ ���L�� 
��m �kl��m���m�l�k�kdl��;�l��� � V��k �� ���: ���l ��L���[)�`�[)�`��� ��r��� ��d(�g�'�f�&�e�% �ǥ0 ���/ ���. ���-L���e � �� ���P�����`�� �� å )��P��Lb���� �ǩ�� � V��`L��`���`�����`�`L�� ��Z
� ����������`PERFECT !�NO BONUS !�GAME OVER��颇 cɢ �)��� � 2����	������ ���<e � ����P�� å )��P����L*�GAME CPMPLETE !�You have defiance�all SIXTEEN STAGEs.�CAN`T BELIEVE you�DID IT, But you�just did it !!!!!�In the last�We appreciate to�buy BALLOON FIGHT�that`s has great�meaning to our�company. So,�THANK YOU AGAIN !� �   PRESS ANY KEY���!	��`���� c� ���e � �� Qɢ �)��� ũ�������� �� ����e � ���l06���� V� ���ee�e� ef�f� eg�g � X��e � ����dl�<e � ��dP�k08���� V� ���ee�e�ef�f� eg�g � X��e � ���P��dk�xe � ���P��2�����Ӆ��� ���ee�e�'ef�f� eg�g � XÀ�����݅��� ����e � �� 2�����Z���ZLk���e � ����� cɩ����A��� ���xe � ��� ��L*�TIMES = ����	�[)�ΰ��` �ȭ������e � ��L.ɜ)�,�/�2�5�8�;�>���+�.�1�4�7�:�=�@�Z
�����b����c� �b�'�(`,'�`�(��'�(� �(��iLJ�d��*� �¨)�* � �)�� ��)�*`
 ,'�`dV�d�)�+��+��V��(��iL����b�


i�Rȱb�


i�Sȱb�U��d�)��Z�V��w�H� �)��� �h ��h��L��X��Y�Y����P����Q��P ��Y�Y�`��P)�P`��P)�P�X����Pi�T8�S��S8�T��0`�� �Pi�T8�R��R8�T��`��	��P�S�
`��P�S�`��P	��P�X�5��"��� �P�R�`i�P`� �P�R�`8��P`��P�S�`i�P`��P�S�`8�ɟ�� �P`���������� ��*��4� �>�����������������$��.�t���~���������"#� ��"#� ��"#� ��#"�@��#"�@��#"�@
��"#� ��"#� 	��"#� 
��#"�@��#"�@	��#"�@,-�78�FG� ,-�9:�HI� ./�;<�JK� -,�87�GF�@-,�:9�IH�@/.�<;�KJ�@12�>?�FG� 12�@A�HI� 12�BC�JK� 21�?>�GF�@21�A@�IH�@21�CB�KJ�@�ij�\]� �ef�bc� ,-�kl�bc� �ji�]\�@�fe�cb�@-,�lk�cb�@
�VW�bc� �QR�\]� N	�XY�dc� 
�WV�cb�@�RQ�]\�@	N�YX�cd�@�ef�bc� �gh�^q� �eh�`a� �fe�cb�@�hg�q^�@�he�a`�@�QR�\]� �QS�^_� �TU�`a� �RQ�]\�@�SQ�_^�@�UT�a`�@���� ���"��"��"�,�J�6�T�@�^�h���r���|���  �������   �������@vw�|}���� xy������� z{������� wv�}|����@yx�������@{z�������@vw�|}���� vw�~���� vw������ wv�}|����@wv�~����@wv������@����������������
��"�/�<�K�Z�i�										
	
		

	
	

		

					

������������������������� �3� 	  
   	   	
	   	
  		 		 �}|����@yx�������@{z�������@vw�|}���� vw�~���� vw������ wv�}|����@wv�~����@wv������@����������������
��"�/�<�K�Z�i�										
	
		

	
	

		

					

������������������������� �3� 	  
   	   	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                \]� �QS�^_� �TU�`a� �RQ�]\�@�SQ�_^�@�UT�a`�@���� ���"��"��"�  �  ,�J�6�T�@�^�h���r���|���  �������   �������@vw�|}���� xy������� z{������� wv�}|����@yx�������@{z�������@vw�|}���� vw�~���� vw������ wv�}|����@wv�~����@wv������@����������������
��"�/�<�K�Z�i�									  �  	
	
		

	
	

		

					

�����ύ& L����7�