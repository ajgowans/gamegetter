� � � � � � � �   0@@P`p��������  @0@P`p�������� @ 0@P`p�������� @ 0  � �����     � � � � � �     � ��� < �    ��� ���     � � � �� �     �  � ���     �  � ���     �� � < < <     ��� ���     � �����     ���� � 0     � �3���     � Www_W�    ? ? �? ?     � ���      �<<<<�    ������    � �� �    ����    ������    �< � �    �0 �<<�    ���� � �     �<�<<�    �<<� �    <�����     ����<��   �\��|\�  0 � � � � 0    0  0     ��<�<�<�<�     �        �0< < ��?    �?0<  ?0<�     �0�?      �� � <0<�     � ��<�<�    �?  ���    �?�<��<�<�    ��<�<�? <�    �<�?�?��     ��?03�?�<�   �p5p7p7�5p5�  � ��0<���   0 � < <�0      ?�������� ?     < ? < < < <     ?�� � < ��     ��� < ��� ?     < ?�<�� < <    �?��? ��� ?     < �?���� ?    �� < <       ���� ?���� ?     ?���� � � ?    ������ ? ?      ?�������� ?    ?���������� ?   ������   �  3 � � 3�                   L��L��	L	�	�	
L
�
�
L��L��L��L��L��H��
J��
J��
J��
L��L��L��L��L��L��L��L��L��L��L�
	
	
	
	            
	
	
	
	            
	
	
	
	            56 (	
78 )*  9:  +,  ; BC -.CC<@AD!/0DDD=DD"#12 >?  $%34        &   '(   56)*   78+,     9: -. B C   ;B/0C@AD!BC<D12DDD"#DD= 34   $% >?       &    '( 6	
)* 8  +,  9:BC-. B  ;DD/0CD!C<DDA12D"#D=  34 $%>?        &   @U PU TU UU       PU TU UU @U PU       UU @U PU TU UU BDDDBDDDBDDDBDDDBDDDBDDDBDDDBDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD�DDDD�DDDD�DDDD�DDDD�DDDD�DDDD�DDDD�DDDDBDDDBDDDBDDDBDDD����DDDDDDDDffff    DDDDDDDDDDDDDDDD����DDDDDDDDffff    �DDDD�DDDD�DDDD�DDDD����DDDDDDDDffff    UUUUUUUUUUUU����UUUU����ffff����ffff������������ffffDDDDDDDDDDDD����    DDDD��������ffffBDDDBDDDBDDDDDDD����    DDDD��������ffffDDDDDDDDDDDDDDDD����    DDDD��������ffff�DDDD�DDDD�DDDDUUUU�	  U	  U  U
  e	  U  U	  U	  �	  �  �	  U  U	  e  U  UUUU   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @�  U  U	  e	  U  Y	  U
  U  UZUU�IDDUVFDDTUEDDfUFDD   @   @   @   @   @   @   @   @UUUUDDDD�DDDD�DDDD�DDDDADDDADDDADDDADDD����������������
   
   
   
   QD�DDQD�DDQD�DDQD�DD����������������  ��  ��  ��  ��
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
     ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ������  ����������*���*���*�������*���ZY���f������f������  ���������  � @� � �� ����
��J��JQ���
��RE��U@��P����������  �����������������������"��j���J���I���j)��U������  ���������  ���U���U��jU��ZU��ZU��fe�����bfe�����bfV�����bfV�  ���������  ��*��V���UU�bT�b�bP�"X�ba�bQ��Q�����*�  ���������  �RUU�RUU�R�U�R�V�R�U�ReV�R�Y�ReV�R�Y�ReV�R�U�RUU�  �����                                                                UUUUUUUUUUUU TUU @UU   U                 P   U  @    @       TU TU TU TU TU T        @P UD@ UP T T  U UU UU UU TU UU UU UU TU TU TU TU TU TU TU TU TUUT AUUQUEUUUUEUQUUUUUTUUUDAEUUUEUUTEUUUUUUUUUUUUUUUUUUUU TU UU QU QU QU UE U UU UU UU UU UU UU UU UU UU                    P   P   T  T    UE  F  U  UUE UEE@  @  @  @  @  @  @  @@ @P  U  U  U @ T U TU@@P@@@@      P     @  @  @  @  @  @  TP           @  @@    P     @             @A@ @ P@ @@ @@ @@ @@ @            @ @   A   A   @   P   @   @                              UEUEA UPQPQTEUDPUU Q AT  Q QU@QEP@U@UUUUTUUTTDP DEUUTQEUTUEEQEEEEQPAUEU T @ D  E EA  AE  UA  UU  U  U  U  U   D   D   D   D   D   D                  P                @PE @          T   U  EU T  TU QP UAUQUEUQPU UUUUQUEU Q                  P P U UPUQATUU   TE     D @PU @ Q   Q  Q    E  TAAP UQPPQPUU QPT EPA  T   @E @  @UTPUUTUUU@UTU@T                        D   TDQ@ETUUT U PU TU @E @E U@PQPU                              @ @@@ DDDPADAUADAUAQUEUEUQUQUUUUUUUUUUUUEUDUUQEEEDQEQTETTDUTUTUUTUTTUU      UP  P  P                  T  D  PD@ UEE@PTT UEPUT@UUE@T UPPEEPED PD PUD A    UUTU  Q  UUT DU UUU DP TT  TT @P  @@@@U@U@PEETUEUD@ DD  TTTET EU UEUUUQAE  Q       UD TUQ UP                              @  Q PD @D  TEU @P @U @ @ @ @ @ @PP@UA@UU@DQ@UA@PUUPPUA@UU@   @   @   @                @  E QDAP EUPEED@AUATAQ@A A A A               @ @@ @ E@ P D@ @ ET UQ UU UU UU UU UU UU UQ U U E U U U U U U@U@@ET@QD @UQ @P PU PU PUEUQUPTDTUQUUQQUUQQQTUUUUTUUUUUUUUUQUUUUU TU UU UU  PU TU TU UU  UU  UU  UU @UU @UU PUU PUU PUU TUU UU UU@UUQU QU UU QU  AQ      @  P        @  @  @@  PUUPUETUUTUUUUUUUPUUQUUU TUU                                PPE UP@U @                                                 @AQ   PAU E  TEUPUTUUQAEUQQT@TUTPEPQUUQTD U     E   @  UTTD PQ D DDQUQDE UU@TU@ T   @@ @                                  @    @  @@@TPDU@UTT                  P    A  A@         TEU@  A U  DT @                         P               @                                        @ @               P                                                   @   @   @@@P            P   T  @U  @U  PU  @U  PU @TT PTU TUT UU@ UU @T@PE@T@TU@UU@UU@UU@UU@UU UU UU UU UU UU UU UUUQU UET UEU UU UU UU UU UU UU UE UE UA UU UU UU UQ  UU UE UU UET UQT Q UT T U EU TU EU UU QP UU UUUUQ UU TU TU                 T                     UUE UU  A UUA UT               PU                             P DPPUUUUAPUUUUU QQ@UAQ     P  @     A   A   A   Q  Q U PU PQU UAUUDQTEU A  TQUU AP AA @      @@@@U@ @ PAU @@    Q   @                @  @A  A  A P A T ATU A ADAD @AD @A @ @        @   @  @  @ @  @  @ @  @  @  @   A            @    @  @@  @@  @@  @@  @@  @@  @@  @@  @@  @@  A@  T@  @@  P@  A@  @  @                                         @PTDPTPPPUPUEPPUDPUPUPUPUPUTPUPEUPEUPUUPEUPUUPUU TUE TUETPUTQ@UUUUTUUTUDUUU@T @  @   P   U                         TUU TUP TU UT PT  P     UQ U                         PEU TUU TTE@UUU DUU TU PUU @UU PUU UU TTUDAUUUUUUUUUUUUUUUUUU  U  U  UQ UU UE UQ U UU  UU UQEUUUEQUUQUEQUUU   @      P  @     T  P  E   E @A QU AE E E TE                       TTPTETQTEQTUAUUU@@U@@UUUUUUUUUTUUUUUUUQUUUEUUUUUUUUUUUUUUUUUUUUQUUUUUUUUUUQUUQiiiifyyyyffqqqqf�����f�������f����fff�����f���f��f�ff�f�f�f��f������fffffff h���'!� :1�'Z!� )2�2>3�2'#�23 �('># �('4 �(- �F'A* �F 'P+ �F'n5 �F'6 �F'n/7 ��'7 �'77 �'P7 �'i7 �'<+
 �<&n, �<-
 �P	7d �x� � � � f� � � � f!!!!f�!!!!!f!!!!ff�!!C!K!S!C!C![!c!f�!f�!k!k!k!k!fC!C!s!s!s!s!f�!f�!K!C!�!!C!f�!f� f!� �!ff� �!fff�!ff�!!�!C!ff!!!!fk!k!k!k!f{!�!�!fffffff�!h'*�!:9�!'Z+�!):�2 'Z+ �2
% % % % #% '% �<';�2 'F# �d-3 �d '-#�dF3�d2 �'((�'7 �<'77 �<'Z7 �<'> �<'i< �<&n, �< ':= �<	 d �2   �    \   W      �  ��  ��  ��   ��  ��������������� ���? ��  �?     �   |   W   �?   �?   �:   �: � �: ��: ���� ���� ���� ���: ���  �                 �� �� �����'�'���'���� ��> �� ��  ��           ��         �� �����'�'�������� '�> �� ��  ��   ��<�? �����:�����:�����[9��zU�[9[�zU�[9[����[9[����[9[�zw�:[�����?�����  �?     �?��<  �����  ������?[�����:[�zU�:[�zU�[9[����[9[����[9��zw�[9�����[9 �����:     �?�?�:�:[9[9[9[9[9�:�?�?    ��    ۪   ۪�? lk>��l���:��������� ۪��  l��� ���� �[��  ���  �oU   ��            �? �? �� ��?�� ��۪����l��k:����:�֫��: o���� �V���  �VU�   ���                         ��              ���  ���?�?\UU�Wկ�
��k��*� ��X%� ����� ��ڧ�  �j��  ���?  �         ��   0 0    � < 0 �0 ��?�5_U� 7��� �UUU �
�� �*�� �*�� 쪮� �}� ����  ���  < �  � �� �? �� � <� 3<� 3<� �<� <� � �� �� ��?  �         ��� ����< ?3< <3< <�< << ?�?������             ����           �WUU�          _UUU��         �UUUUU�        pUu}UU�        \Uu�UU�?        WUu�UUY�        �UuuUUV�      �UUu]UUU�      �Uu�U�U�      p��UUU?W�      p�WU�?\�      p�\U�?p�      \�\U�?pU?      \�\U�?p�?      \�\U�?pe?      ��\U�?pU?      \�\U�?pU?      \�\U�?pU?      \�\U�?pU?      \�WU�?\U?      \���WU?WU?      \U\U�UU?      \UUpUUUU?      \UU�UUUU?      \UU�WUuu?      ��U \Uuw?      �]W �Uuw?      �]W  �}?      ��W�  �_U?      \UUU  ��?      \UU�?  ��>      \UU�� ��:      \UUU? ��:      \UU��?��:      _U����׫�:      _U�5 W_��>     �^U}5 \}��?     �^U_5 \�U�?     �z�W5 \�W�     �z�U� \U_�     �zUUU�_UU�     ��UUUUUUU�     �UUU�UUU�     �UUU�UUU�     0W�UWU�V�     � _iU�UUZ�     0 pUU�UU��?    0 pUU�UU��    �� �UU�UU �    �  WUUU�  ��  0  UUU�  ��  0 ��_UU� <�   0 ����0��  �     �3��     �     0��          ��           ��>      0��    ��      ���   ��        ��   �        ��             ��            ���             ��:             ��             ��             ��              �?                 ����           �WUU�          _UUU��         �UUUUU�        pUu}UU�        \Uu�UU�?        WUu�UUY�        �UuuUUV�      �UUu]UUU�      �Uu�U�U�      p��UUU?W�      p�WU�?\U?      p�\U�?pU? �   \�\U�?pU? 0   \�\U�?p�? 0   \�\U�?pe? 0   ��\U�?pU? 0   \�\U�?pU? 0   \�\U�?pU?    \�\U�?pU?    \�WU�?\U?    \��UUU?WU?    \UUUU�UU?�    \UUUUUUUU?�    \UU��UUUU?�    \UU��WUUU?0    ��U� WU]]?0    �]W� WU�]?    �]W� WU�]?�    ��W��WU}_?�    \UU��UUUU� 0    \UU��WUUU�0    \UU�U_UUի    \UU��UU��    _UU���UU��:   �^U�WU�WU���    �^U�UUU_U��:    �^U}UUU}���   ��^U_UUU�U��    0�z�WUUU�WU?    �z�UUUUU_�   � �~UUUUUUU�   ��UUUUUUU�    0�UUU�UUU�     WUU�UUU�   �  W�UWU�V�    <  \iU�UUZ�    �  pUU�UU�?        pUU�U��        �UU�U�         WUU��          |UU� 0          �_U� 0          ���0          0  �          0  �         �            �
  0��       ���  ���?     ����  ����     ����   ����     ����   ����     ����   ����     ����   ����                                                                                               �    ��     05     L     S    ��     <�    ��:    ��;�� ��|� ����0�뿯� �Ϭ��> ྪ� ��Ϊ�  ���� ����� ����� �����  � �?              �    ��     05     L     S   ��  �  <�  0��:  ���;���|�������
뿯� �����> ̿���  �Ϫ�    ��� ��� 󪪪 �����  ����?  ��?    �?         �        p       p       �       g      ��      We   �?�UU   ��s��    ��=�    ����    ��U�>    �W�� �  �W��� ������� �������0��?𪪫?<��?�����?���������å�����p�����  \j�:��?  ן�: �  ?��     ��     p��     ���       p>       �         <    �  �   �? �<  �� �;;  �� ��;  �� �>  ��; �>  ��= ��>  �z� ��  ��� ��  ��Yê�   Weê�  �UU�����p�Ԭ�� ��=ԫ�: ������ ���U��� ���W��? ?���W������������� ������� ���?   ����?   ����   �� �   �   ��   3   �?   0        @ � �
@ ��(  :�   0�  ��  p�  ��  ��6  �{?  �� ���9 p��: ��� ���   ��  ��=  ��  ���  ��<  �          �       �k=       ��;       ���       ���       ���       �k    ��� ��?   \�� �v�   ׭; ��k  W�; ���  �� ���                                           ��������? \m۶m۶m� ׭뺮뺮kW�뺮뺮����������                                        �  o� ��������i���6���:�jj髩�ټ��>��� \5  \5  \5  \5  W�  \5  �     �?  p�  ��  �� �� �� �� W� �� �Z �i �� kj �� p�  p�  p�  p�  \U p�  �?                    �? ��?�i�篖�\j�欕�6� ��               �  �6@ �9  k:  �9 ��6 �e: �f: �f pi �i k� �> _� �?       �?     � 00     ���3     �:W�2     ��U�2     �zU��     �zU�p     _U\     \UUW     W���     ����:     � �?    ����
�    �����    ������   �U��:4   �zUժ�   ����@�  p�*T� 3 �^�JU: � ���V� � �����,��ϭ�_U,�7�U�5���_�Uuu5�0p]�_U��5����UuWU7�?�_�U�]7�
<���U�5�
���w]w7��5���WUU5��Ww�5�U���WUU5�� ���u������_UU]�?��_UW]U�>�UUUu�]��UU]UU� �~UUUUWu5 �_UU�_UU�  WU�3pUW� \�03pUU� ��03pUU� 0�3p�U� 0�pUU� 0�pUU� � pUժ    pUժ     \Uժ     \Uժ    WU��   WU��  �UU��  3sUU��  3�_UU��   ��WUժ:   �UUU��   WUUի�  �UUU���   �UUի�    WU���     W���     ���      ��                                        �?     � 00     ���3     �:W�2     ��U�2     �zU��     �zU�p  T  _U\  @  \UUW  E W���  U ����:   � �?   ����
�  D�����  T������  �U��:4 @�zUժ�   ����@� p��*T� 3�^��JU: ����V� � � ����,C�����_U,�7p�U�5���_�Uuu5�0p]�_U��5����UuWU7�?�_�U�]7�
<���U�5�
���w]w7��5���WUU5��Ww�5�U���WUU5�� ���u������_UU]�?��_UW]U�>�UUUu�]��UU]UU� �~UUUUWu5 �_UU�_UU�  WU�3pUת \�03pUժ ��03pU�� 0�3\խ� 0�0�WU�� �03_Uժ� 03�UUժ�  0�UU���  �_UUU��>  pUUUի�  pUUU���   \UUի�   \UU���    pU���    pկ�?     ����      ���                                              ��???���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �@�@�@�@�@�@�@�@ AA A0A@D@APA`ApA�A�A�A�A�A�A�A�A BB B@D0B@BPB`BpB�B�B�B�B�B�B�B�B CC@D C0C@CPC`CpC�C�C�C�C�C�C�C�C D@DD D0D  � �����     � � � � � �     � ��� < �    ��� ���     � � � �� �     �  � ���     �  � ���     �� � < < <     ��� ���     � �����     ���� � 0     � �3���     � Www_W�    ? ? �? ?     � ���      �<<<<�    ������    � �� �    ����    ������    �< � �    �0 �<<�    ���� � �     �<�<<�    �<<� �    <�����     ����<��   �\��|\�  0 � � � � 0    0  0     ��<�<�<�<�     �        �0< < ��?    �?0<  ?0<�     �0�?      �� � <0<�     � ��<�<�    �?  ���    �?�<��<�<�    ��<�<�? <�    �<�?�?��     ��?03�?�<�   �p5p7p7�5p5�  � ��0<���   0 � < <�0      ?�������� ?     < ? < < < <     ?�� � < ��     ��� < ��� ?     < ?�<�� < <    �?��? ��� ?     < �?���� ?    �� < <       ���� ?���� ?     ?���� � � ?    ������ ? ?      ?�������� ?    ?���������� ?   ������   �  3 � � 3�                   lF�F�F,GlG�G�G,HlH�H�H,IlI�I�I,JlJ�J�J,KlK�K�K,LlL�L�L,MlM�M�M,NlN�N�N,O,VlV�V�V,WlW�WlFlO�O�O,PlP�P�P,QlQ�Q�Q,RlR�R�R,SlS�S�S,TlT�T�T,UlU�U�U,VlV�V�V,WlW�W             $%  )*  $%   &'(                      !   " #  	
               !"                         	
              !"                                       !"                         	
                                                                    @         @  @ @                      P UUQUUTQTUUUTUU  PU @                   P        PUTQPUUUUUUUDUU TU  TA        @    @@    D        UUQTPQTTAQUEQUQUUUQPE QP  P@                      PUUPUUPTUTUU TUU TUU TUU UU    U  T @   A @UA @               UP  U@ U    @       D DD  U         @@  A               @           A@U UUUU  P           QT  U PU @TU  TU UU UU  TU    @  @@  @@P          UUUUUUUUUTUUUEUUUUUTTUUUUUUUU   A @ ADA  D      P TT @UT@UUPQQPUUPUUTTUUQTU UUU @UUPUPT@ @     U UUT UQU UU EU UU UUU UQ UUU UUU UU UUU UUU U     U      U@U@UQP@EUQ@UE@UQE@UU@UE U UUPUUUQ@QU @ TUU UUU@UUUEQQQE@UE  QPUTUUPUUUUQUQUUQUAEQAPQDPTUQQAUQ ET EPUTUUEUUUUAUUUTUUUUUUUUUUUUUUUUUUUUUUUUUUU PUQUQEUAEUDDU   U  U T U Q U@QT@UU@E@UUPUUTUAE@U TD@UUPQEPUPUEUEQUU UQQ QUU PU  TU PU T  UEPTUPUPUUPUUPUUPEPUUPUUPQUPUUPUUPUUPUUPUUPUUUPPUUTPETQPUUE@UUQUUU@UUU UUUUUUUUUUUE UUU UU UU UU U   PPAPUDPUPUPUPUPQU P  ATU                     @UU  PU  P  P  P  P  P  P    T  T @T TT U PUAQ  QQ                         P   T @ T@UUUUU@UUTUTQAUUUUUEEP @T P  PU  T  TPTUTUT  PT  TTTU@TTTTTATTTTET@UUUU U   U   U  U  U  U  U@U A AUP U UAU EDA UU UU U             UU TU        P AUQ@ U@QEU@EPU@TPU@EU@U                       @     UU     P UQPUUEUEUUUUUTA               @   T   T   P   @  @ TUP TUPT  TUPU @  P  P  T  T TU TUUUUUQPUUA TU@UU@AUUTAUPUAUUQUU PP           D  D  P  Q UPUP@EUAUPEEUEUUUEU@EUEPT UUU UUU PUU  P UQ PPP P@P P UTUPEPUTPQUP    @  D   T     PE @DPEPU TPUEUPUUUPTU QUUPUUPU@ P@  @  @  @  @  UU UUU UUU @  E  E P P@PUPUUP                                   P   P  P  P  P P TU TUU                 U   U   U   U  U U U@U U@ UP U UUUUUUUUU                                              @U  @U  @U  P  P                             @  P  P  P  P  P  P  P UUU                                               U  @Q  U @ED TU                                            E   U  T  U  Q                P   T   D  T  EDUQUUAPUU TUUUDUUQUTUUU EUPADTUUDTUPUPEPTQUUUDEUQETUUU UUTUUU       UUUUQUUU UUU UUUPUUQUUUUQUUAUUUUUUUUUUUUUUUUUUUUU       PUUU@U T            U  U  UUUUUQUUUUTUUUUUUUUUUU       TUQU@UTUUU                       UU UUUUU@  U  @UPUUUTAUTEUQUUUUUUUU                   U  @E  UT PUUU@UUT UUUUUUTTUUUUUTUUUUUUU            U  QTUUUUUTUUUUUUUUU   @UUUU UUUUUAUQUUUUUUUUUUU                       U   UUU   @UUUUQ@UUUUUUPUUUUUUUUUUUUUU                                UUUUUUUUTUUUUUUUUAUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUQUTUPQUPUEU PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUUUUUUUUUU   QQPEE@Q UU PUUU UUUUUUUUUU UDTU@@ EU UQUAEQUDTTUUU@EUUUUUUUUU   PUUUUPAUUU E@UUUTUTUPUUUAUUQPUUUAUUUTUUTUU@QUPU  T PUUUUUUPEUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUEUPUUQU   U  UUUU@UUUUUUTUUUUUUUUUUPU@UD@T TTAPUTEEUU QTQ UUU PUUU  UUUUUU@UTUUUUUUUUU UUUUUUUPUUU@UUUUTUQ UUUUUUUUUUU   @UUUUUUQEUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUUU UUTUU TUUUUUUUUUUUUUUDUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU@UPUUU UUUUTEUUUUUUUUUUUUUUUUUUUUUUUUUUEUUE@UU UU T TQUU UUEPU@UU   UUUUU@EPUUUUUUUUUUUUUUU@UUUTUUUTUUEPUU  UUTU@U T  UU@UUUUUQUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUPUTA QAEE TUUU @EUUUUUUUUUUUUUUUUUUUUUUUUUUTUUP@UUQUT TUE@ UU@UUT  PUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUEUUUUU @UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUEUUUUUUUUUUUUUUUUUUUUUUUUUTUUUUUUUUUUUUUUUUUUUUU                                               U @UD TQUTUUU TUU                                        UU  DU UUUUUUUUU                             P @UU PEU UUUUUUPTUE   U                             T TQ UUEUUUEEUTTTUUUUUUUUUUUUU @U                            U   E TEUUEUUUUUUUUUEEUA                                                            TP UEUUPETT PU                                                      UUUU  ���  ��������� ��� ��� ��������������� � � � � � � � � � � � � � � � � � � � ������ � ��������������������������������������������� � � � � � � � � � � � � � � � � � � � wYgYoY�Y�YgYoYwY�Y�YgYoYwYgYoYYYYwYgY�Y�Y�Y�Y�Y�Y�YwYgYoY�Y�Y�Y�YoYwY=ZZZZZZZZZZZZZZZZZ=Z%Z%Z%Z%Z-Z-Z-Z5Z5Z5Z5Z�Y=Z=Z=Z�Y�Y�Y�Y=Z=Z�Y�Y�Y�Y=Z=Z�Y=Z=Z=Z=Z?ZMZfY�'� 'd#�( '7#�(' �2 'd �2'2 �2 '< �2'##�( 'K#�($
 ��<&<&"&Z&�<'7"
 �'  �<'F  �<'d  ��'' '7' 'd' ��'
!�<'(!�<'F!�<'
!�<'<! �<'! �<'_! �<��&" 'K �('
 'k 	% d �([[[[=Z'['['['[=Z/[/[/[/[=ZW[[g[o[w[G[_[7[O[=Z�[�[?[�[�[�[=Z�[�[�[=Z�[�[�[�[=Z�[�[�[�[�[�[=Z�[�[�[�[�[=Z�[?[G[o[�[w[=Z'[/[[=Z�[=Z=Z�[�[�[�[�[=Z�[=Z=Z=Z�[=Z=Z=Z�[=Z=Z=Z�[=Z=Z=Z=Z=Z=Z�[fY'(�':(�'Z(� ')#�2 '>#�2 'U#�2') �('>) �('b) �('
. �F'-. �F'P. �F'd. �F't/2 ��'/2 ��'' '7' 'n' ��'* �<'<* �<'d* �<'+
 �<'<+
 �<&n, �<-
 �P	 d �d  ��    ��   ��   ���  ���  ����  �Ϗ�  ������ �����?   ����   ����   �      <                  ���  ��� ���?  ���� �Ϗ�?  ������  ����? ����� � ����   �      <   � � �� �� �� 0� 0 � �  �  3 �8 � 0 < � � � � � � 0 / # + � � �2  3  �  �  , 0 � �< �2 �� �� �� �     �?  W� ���p��p��������������� �� � ��  ��          �� p� \�: ��� ��� ��� ��� ��� ��� ��? ��  �:  �:  �:  �:  �:  �  �   �* �������*�*�������� ����
  ���  +�� ���
  ���  ���?  <��   �?                                      �    ��*   �>  <��
  ���*  �*�*  �*��  �
��
 �
��*   ���       �  �  "  �$ ��	�`"	(b&�`&�X�	P	V ThU� ��
     �       � � � ��$��$ �$	H�	Hb@	H@	ET�U�  �
 ��???���  ��3   ���:   ���;   ���   ����   ���?   ���� ����? ������ ����  �?��    ��     <                  ����  ����:   ����  ����?   ����? ������ �����  ������?�� ?  ��     <      �?       0��     � �   ����  |U�  < WUU � �_U5 �0  �U� 3   WU 3�  \U��0�  WUU�3�  _UU]?� ����_�� pUUUUU� \��_UU� WuUUUU��U��UU�_��U��U5W���0 _5kU� ����V�  ����� �UU��� � ������� ��W���?8 ��_���> 33s���� 0����;   �� ��:  0�����:  �|����: �0s����� �3_����� �<�_���� ���W����|�UU����_UU����_�_���W�W��ժ�����W���꯯�_�������~������������ ���ת� ���� �  ���_� �  ���^; �   ��^ �   ��_ 0   ��� 0    ��     ���    �UU:   �U��   |U���   �W��    p��      \�      \	   ?   \�? �:   pU���   �����     ���        ��       � �      ? 0 ��  ��� |U�    � WUU   ��_U5   � �U�  3  WU �0  \U��  WUU���  _UU]?� ����_�� pUUUUU� \��_UU� WuUUUU��U?�UU�_��U��U5W���0 _5kU� ���V�  ���� UU��� � ������� ��Wտ�?8 ��_U��> <3sU��� ���U��; ���� ��: ��W����: �U����: WU������ WU�_կ�� ���UU��� �zUUUU�����UUUU������U��{�����������W� �����_� ��ꫪ~� �����{�  ����z0  ����z0  �ꯪz   ����z   ����z    ���~�   ���_p  ���� p     � �     7 �5    �5  �    p  \   \  p   �   p�  �5   �U��_    _UUU    �UU�      ��                                            ��        �     �  �    �       ����?      �\U�   
�ʫ���  �
0����=     �����  ��?𿫫=  <   ����      ��?    �� ���       ��        <                      �        0<        0�      �� �    �        ����      �sUU      ���5      ���       ��z      ���  ��? <0�    ����       ��        �        �       ��        �?       ��       <    �;    �    �   ��   �? ���� �����,�������������������������������  �?  ��    �    �    �;     <     <    �;    �    �   ��  ��? ���� �����+��������������������������������� ��?  ��    �    �    �;     <           � ��� ������������:���:���:��?���������3��03  3   3   0      � �� ������������������������������������3��3�� 0�� 0�� 0��   �  ���    ���   ���:   3��   ���� � �_   ��W6  �W�W5 �WU�g6 p���\ \?��� �̼:  ��3�  w���  W���   �      ���    ���   ���:�� 3��pU���_U� �W�5  �WU6 ��W�5 �U�WU6  ��_�533��\f�̿:pU����� ���   ���                        ��    of?  ��� � g> ���� ��gf�����9gffff朙ٟ����?��?             �   ��   lff  ���9  ���  3;�  37g ; � ���f ���� lfff ���� �gf�   ��        0 �   0� �   �� ���� ����; ��0��: �?�� �>�� ����   ���:  𬮮� 0��3 0�?�0 0   �        ? ��?���:�>���8�;�?0��:�?3��>�3����3�  <���  �|f��0��0�0   0                       �?  �� ���������;���?<��?/��;���?�����  � ��� ������ �� ��          �� ��? ��������������?�� �� /� ��  ��  ��  ��  ��  �� �� �� ��?  �>  �?  �               �     ?  ��      �     � �      0    <PU0     CU1    \�C��    �P��  � p���    �� �  �U= ��    0� �   ��p1    05 �  �   ?0p    05 �  �  �@�p���?  � � �U�p����L ��� 0T�������L ��L��ż�VU�:L �\Sp1�jUUU�L �p�� p̪UPU�O \<�5 \�ZUTU�N pA W �Z@U��N �W � ǬVP���z  �     ǬU T����         �UU���         �UUU�W�: ��      ׫UU��W�: <      ܯZU��_�: S     ܯ����z����     0���������     0�����0�     <������pp     �:���Lp     ��:���� _     ��� ���^����      ��� ���5p=      ��������Up      ������? �p      ���� �   p     ������:    ��    ����?�     W    ��
?��      �    �����             0���              ���               ��                                                    �                00                L�                S���            �\����           �4𪪪�          �4��UU� �        0ͪZUU�:�       �3�jUTU�U      L�VU UU�SU1     �TL�VP���W1     �Tq�U T�����1     0Uqk U���>��     0��jUAU�� �     L��jUUU�� �     L��jUU��U� �     S��V���W� �     � ������^� �     � ̬���z� �    �4 �����z�  �    �4 �������  �    �4 <�����1 ��    �4 �����1 p5    �4 ��: ���1     �4 ��: ���1�\=    �4 �����*�10]� �  �4 �������1L__�� 05 ���*�p�\sU= 30= ��*�p�4��� �O ���� p�5�    P �¯�? �UW�?  \�  +���  �U\ 0  �?  ��    � pU5      �      ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               PAUSE$PRESSaSTART$STAGE$ONE$TWO$THREE$FOUR$GAMEaOVER$HIaSCOREb$YOURaSCOREb$CONTINUE$END$ITaISaNEWaRECORD$eBONaTREASURE$CLEAR$DRAWINGaBYaBANYONG$MUSICaBYaXIAOLIWAI$PROGRAMMINGaBY$XIECHENGWEN$ ����� �&�+�5�?�K�T�X�i�w�}�������6�F�V�f�v���������Ɓց�����&�6�F�V�f�v���������Ƃւ�����&�6�F�V�f���v�������  ��  �������  �<<<< �� �?  �<< <� <<<�   �?�<<<<<�? <  �< < � < <�  �<<< �<<<<�  �?<< < <     �<<<<�<<<<�  �<<<<�? �� ��00�?<?��<<<<�<<<<<<��3<<0  0<<��<<<<<<<<<<��?<0<�<< <0�?�?<0<�<< < � �3<<0 ?0<<���<0<0�?<0<0<0�����������?    ���<0<<�<<<��� < < < < < <0�?�<<?�?�<�<<?��<0�0�3�??<?0�<<<<<<��<<<<<<�< < � �<<<�<����<<<<<�<<�<�3<0��<<��������������<0<0<0<0<0�<���<0<0�����?�<�<�<�<�?<?<??0� � 0??��<0�������?<�� <00�?    �    �                              ��    0 � ���� 0 ��33030�3�                    �  �� � ���� ��                         �            �  �?00�?���?00�?  �            �              �   �   � � ��� � ���� ���      �   �   �                         �  �< ���� �0��   �                         �  ��  _��WW�UW�UW=��W=�U]=�Uu�W _� ��  �                      �  � �:���TUj5����: �  �                         �
� �*������������� ���  �*  �
  �  �                            � ( W��f pU=�rf: pe:��j( �  �                      �  �  ��  � �  �  ��  �� � �� ��  �  �                       ���?� � � � ���?                  ��� � �d���<�P������ �������\�x�L���^���cdNd7d=d(d)d*d+d,d-�2�.d/d0d1d2d3d@dXdYdZd[dpd{dsdtd�dld�d�d>dvdu`���F�d:d<� ����wi ���� ����'�'�� E�`���F�d:d<� �����wi �橴�'�'�� E�`� � � ����� �����d<�Q�R�� �� E��P�S����O�T����d:���2�� ����d��	 ��Q :�P :�O :�}���� ��R :�S :�T :�dQdPdO���'�'��`�O�T�P�S�Q�R�<����	 ����Q :�P :�O :��:���'�P���� �� b� b� b�'�� E�` E�K����
 ��_���� �� �q�
��K��d�; ��  ��m������3�� v� b�
��a�; ��q���
��K�dq�ũ�q�
��_��� v� b�
��a�; ��q���
��_���q��dq�
��K�L!� v�`d{d�� ��i
�H��i�I���J�8�<�K�9 j�d&d: C���&�H�i��I�� ��Ii;�� ����r�I��Ii;��H�� ��Hi��dr ��d: 3���8��9� �
��g���g���ՊeH��ۊeI� C�����d� s��H��I���8�<�9d��d: C� ��`d1��: ��  ��!ɿ�� b� v�d:d1 �d1����怀�d��� b� b� v� 3����� �dm�D����m�:����m�0����m�&����i���	�Pi�P��	���m�� Q�`�1�-�
�1 3����
��g���g���ՊeH��ۊeI� C��`�w
��{���{���z:
���ȱ�`� �����������`ƃ�F���Ƅ�F���ƅ�����������������ÊɊ��������ϊ 	   	   	    	**H�Z���& E� ���8��9� �������� �� Ջ��r�������������� ���9 ����������9�� ����D� ՋL� Ջ Ջ����9��� � ǋ�i�� ������ ǋ�8��� ����� ՋLe����� Y�d�'�'��z�h`�
���������d: C�`H� �& �����&h`H��'�'��h`�Ԍ ������?��?�� ���������?�� ���������?�� ? �����  ?� ? �����  ?� ? �����  ?� ���������� ����������� �����������  �����?�  ?�  ���� �  ?�  ���� �  ?� ������ ��??� ������ ��??� ����� ��??�               ?������� ?  ?��������?�?  ?����������?  ?��� ����?  ?��� ����?  ?��� ����??  ?���������??  ?����������?  ?���������?  ?�� ������?  ?�� ������?����� ������?��������������?�����������?��?���?������� ?��                              d��� �������(�8�\�9 ��d:d<������ ��  ��� E�`�����������������������������������������UUjUUUUUUUUUUUUUUU�U�UUUUUUUUUUUUUUUUUUUU)UUUUUUUUUUUU�_UUV VUUUUUUUUUUUUUUUU)VUUVUUUUUUU�U�WUVUVUUUUUUUUUUUUUUUUU�VU�UUUUUUU�U�_]UYU�ZUUUUUUUUUUUUUUUT�Z�ZUUUUUU�WUU�uUeU��UUUUUUUUUUUUUUUTUU�VeVUUUUUU}UU�WwU�VU VUUUUUUUUUUUUUUTTE%U�UUUUUU�WUUU}wUUiUUXUUUUUUUUUUUUUUQQUQ�fUUU�UUuUUUUuwUU��UXUUUUUUUUUUUUUUAUU�VUUUW_U_UUUUU]UUUUY`UUUUUUUUUUUUUUUUUU�UUUUW]�UUUU��WUUUUY��UUUUUUUUUUUUUEUU�bUUUUW�]WUU� �_UUUYU �jUUUUUUUUUUEUUQ�YUUUUWU�UU� ��UUU�UU�UUUUUUUUUUUUUUiUZUUUW�uUU�<�WUU�UU `VUUUUUUUUUUUEU���UUU]u]W���S�\UUU�jT`VUUUUUUUUUUTE�j%"VUU�]�U51�0�EQsUUUUeU`VUUUUUUUUUUU���*XUUU�u]]�W3<E�UUUU�UaXUUUUUUUUUUUU�jU�`UU�u]WWsT�����UUUUUVeXUUUUUUUUUUUU�YU��UUu]���LTì �WUUUU�j�UUUUUUUUUU�YE��UU]�u��L�����WUUUUU�U�UUUUUUUUU�jVE��UU�u]�5G5�����WUUUUUUVU ���VUUUUUT��VE��VU�]W�:G�����WUUUUUUYU   hUUUUUU��VU��V�uUU�>G������UUUUUUU�ZUUUU�UUUUUe�EVU��h�]UU�?̰�_UU�UUUUUUUU�jUUUVUUUUi��UTU*�u]UU=�0��UU}UWUUUUUUUU�ViU�UUUUY�jUEU��uUUU��UU_WUUUUUUUUU��VU ��ZUZ*hUUU��]UU�
���WUU�p����UUUUUUUU�j   UV��UPA��]UU�*���UUU��   _UUUUUUUU���������UAE��WUU�� ��UUU7�5   pUUUUUUUUUUUUU����UEEU*WUU���_UU5�5   �UUUUUUUUUUUUUe�V�UUU�WUU����UU�s5 ���UUUUUUUUUUUUU��ZUUUU�UUU��
�U�U��s5 �p�WUUUUUUUUUUUUe����VUQ�UUU��
UUW�_5 �\WWUUUUUUUUUUUU���*hjUQ�UUUժ
_��WU5 ��U]UUUUUUUUUUUU��(R��VUuUWUժ
_?��WU��U�U]UUUUUUUUUUUUjU��ZQZUuuWUժ
_� _U�U5WU�U�_UUUUUUUUUUU�V���XUuuWUի
_� \�WWU�U}�UUUUUUUUUUU�Z��eTXUuwWUU�
_� \UWWU��WUWUUUUUUUUUU�jj�ZFTUuwWUU�
_5�W� WWUUwUU]UUUUUUUUUU�Zf��UT�ww�WU��_�U WWUU_Uu]UUUUUUUUUU�U��ZY�W}�UUU��WUU� �� WUUW��uUUUUUUUUUU�����ZuUu��UU��WUU5 �5 WU�UU�uUUUUUUUUUU�jU��V]U�]WU��?WUU5�s5�UU�U]WwUUUUUUUUUU�ZU��Z]U�u�U  |UU5_�UUuU]]wUUUUUUUUUU��ZU�V�U�_�  �UU���pUUu]u]wUUUUUUUUUU��VU�ZU�W_�?  �WU�_? pUUuuu]_UUUUUUUUUU��UUUUUU��?   W5�UU�  \UU�uu�WUUUUUUUUUUU�VUUEUU5    �U� ��  WUUUu}UUUUUUUUUUUUfjUUUUU�   ��UU�    �UUUUu�WUUUUUUUUUUUU���UTE�   p�UUW?   \UUUU�_UUUUUUUUUUUUUU��YUUU  \UUU]�   \UUUUUUUUUUUUUUUUUUUU�UUUUU= �_UUUuU  WUUUUUUUUUUUUUUUUUUUUUUUUUUU�pUUUUuU �UUUUUUUUUUUUUUUUUUUUUUUUUUUUU5\UUuU]U |UUUUUUUUUUUUUUUUUUUUUUUUUPUUU�_UUuUWW�WUUUUUUUUUUUUUUUUUUUUU�W�_UUUUuUUU���]�_UUUUUUUUUUUUUUUUUUUUUU�W�_UUUU]UUW��uuWUUUUUUUUUUUUUUUUUUUUUUU�W�_UUUU]UUWU�uuWUUUUUUUUUUUUUUUUUUUUUUU�W�_UUTU]�U]U��ըUUUUUUUUUUUUUUUUUUUUUUU�W�_UUTU]�U]U]W7 j��UU�ZUUUUUUUUUUUUUUUU�W�_UUUU}UWuU]]�
���VU)�UUUUU�UUUUUUUUUU�W��_�UUuUWuUu��� ��Z���VUUUU�VUUUUUUUUQ�W��_�UAuU]�U�_U*����*��VUUU��ZUUUUUUUUE�S��_�U�U]�UuUU�������ZUUU
aZUZUUUUUUU�G������UuUW}U���� ���hUU�@�j�hUUUUUUU�W�����WWuU�_UUQ�   ( ��ZU) �j
jUUUUUUU�W������WW��UUUDU�  ������@����UUUU�UU�W����U_U]uUUTUUU* ����j
PT���VUU�*UU�W����U_U�_UUUUEUU�  ��� Eef�jUU) UU�W����U_UUUUUUUUUUAU����Z% Pd�
��Z� UU�_��_�U_��_UUUUUUUUUUUUU�
 TU��* ��
��UU����_�U_��UUUUUUUUA T�*  U��*�
� (�UU����O�U_�W}�WUUUUQUUUU)  U�U��*���UU����_�U_�W�WUUUUUU��� @UQ����
* ���UUUUUUUUU_�W�WUUUUQAT�
   (  ���� ��UUUUUUUUU_�W�WUUUUUU]��
�   ���(  ���UUUUUUUUU_�W����_�U������ ��*�
���AUUUUUUUU_�W����_�U��?�U��ߪ���  ����EUUUUUUUUU�W��W�_����_��U��_U��( �����UUUTUUUUUU�W��W�_����_��A�WUUUU (
�TUPUUUUUU����W�_����_��U�SUPU� ��  ��UPUQUQUUUU����W��������E��UU�* (���UQUEUAUUUU��_���W��������U��U�* ��* ���UUUUUUUUUUU���W�_����_��U��U�   ������UTTTQUUUUU���W�_������Q�WU�  �������UUPUPUPUUUUUUUU�W�_����_��U�SUU�
  ����UUUUUUAUUUUUUUU�W�_�}U�_��U��WUT��* ����UUUUUUUUUUUUUUU���_�=U�������_UUUU������UUUUUUUUUUUUUUU���_�=T������UUUUU�����UUUUUUUUUUUUUUUUQUUUUUQUUUUUU   UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUQUTUUTU����������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ���ة��  ��� � �� � �� �ύ& � t ���d���� � �������� E�XL �H��'��'�(��(�)��)�*��*�+��+�,��,�-��-�.��.�/��/�0��0�1��1�2��2�3��3�4��4�5��5�6��6�7��7� �	��	����(�h@H�Z�' )������ �� r�׍# �$ �% (z�hX@                                                                                                                                                                                                                                                                                        ;�n�׍#  Z���& E� �dTdS��R��y E� � � ����� )� Ӎdw��d�idzdm��� ������ �� )� �©�y m�dxdOdPdQ��в�q�dwdz��dz E怼` �� q�dAd>��BdCd'dDdF�F�E�G 4� d�` � F� �� �¥p���Z�l�����y m�dx E��� )� � ��L�í  	������L�� �ĥ3�5���C #� d� �� �� �� �� �� �� _Ԁ� � �� �� �� �� _Ԁ� d� �� �� �� _�L�¥�� d� �� �� �� �� ��L��d. d� �â ��������� �� E� � � ����y m�dx ���w���wdzL��dwdzL��`� �d�	��  �� #� b� b� b��������� E�`�w�����y m穀�x���y m�@�x`� ����.�	���
���� � � E���� E�I� E�����`ڢ ������x������	 � E������`� ���� � E�����`���� �ˢ �d����	� �⊨ $ĩ��d����`�  	��L�� v� �  Z��)��& ��ydx ��i���Ae����:d<�  �� b� v�  	��� b� v� ������  �� ��`dd��8��9�w
�������������	� ��ȱex�� Z�
���ȱex�zd: C���`��>�>��	�i���d>d�i��ƥw���@`� ��/����� ���� ��`�A�i���eB�� ���� ��` Q� 5��8��9�A��B��w
�������������	�@
���ȱex��>�?� �?��
���ȱex�d: C�����?i�?�i��� 5� Q� ��`�'�]�
�'�����;� �C���C�AdC �ťA�,�i�A�dA�Bd>�w�%�@���@�d@��>�� � ����  �ƀ� ��`ک���� �d����x8�0�x��� ����8�0��(���եG�%�F�$8�0�F�G� �����8�0������{�	�|8�0�|�}�` ��i��V���ei�j�~�i���W�f�8��kd:�)�<�U� ,�Q :�P :�O :� @� g� ��`ڥe��f�d:�U�<� ,�d�� ,�ʀ�� ,��`ڥj��k�d:�U�<� ,�i��
 ,�ʀ�� ,��`�V��W�d:�U�<�Q :�P :�O :�`�Z�U�<d:�~���� ,� � ����#ə�����
����� ,�������֩ ,�z�`�d�*��&��6��(��$��*�	�0�����P�� ��&�P����� ����� ����� �����Oe�O�Pe�P�Qi �Q�`�(�x��( Q� �� �ե{� �ԥ���F�"�G�#�$�F�%�Gd� N˥"�F�#�G� N� �� �� �� ��eD�F�eE�G �� �� 4˩�: �� �� �� Q� ɥ{� �� y�`ڥF��G��)
���ʅ轂ʅ��8��9�.�J� ���`�Z�.�a�w
�������ȹ������ �d���:��:��:��F8�x0�#�I���G8��0���I��� �ɀ��кz�`�{���E�F8�|0�:�I��1�G8�}0��&�I������� Y� m� ���y m� �� �� g�`�F�.��� ����d���� ��`��i gǥi� �ɥd����l�`�d.���pdm �� N� �եGi�h�F�g ]��`�/�?��/ ]ʥhi�h8��� ]ʀ%��:�F��G� ��dp�d���i�d @� gǩF�.`��8��9�g��h����ʅ轂ʅ��: ��`a���]���Y���U�  	����	 � �L˭  	���� � )ˀZ�  	���� � )ˀI�  	���� � ˀ8�  	���� ˀ*�  	���� ˀ�  	���� ˀ�  	���� )ˀ `�D��D`�D��D`�E�0�E�E`�E�l��E�E`d���F�H�G�I��J��K j�`�F��G���8��9d��d: C�`H�Z�H��I�dd� �����2���%&�����(�d�i(��i ����J����d�H����Kкz�h`�)���) �� � Z�`� � ��� ������`�Fi�8�	�� � �������� ������`do� � ���L���<� � ��L������(8��(�s����(�(�d�� �̀[�� ̀b���<��L LπB���<��< gπ2���<��, +π"���<�� �π�	���	�
���  �̀��� �<�P����L� ;�` ��8�0�8��(�
�(8�0���� �<�P� ��` ��<���8��&�
� ��do����(���� �<�P���o`ڥo���L�͢ � �������L�ͩ� ���:�( �΢ � �������[�� ���:�( �΢ � �������7�� ����( �΢ � ��������� ����( ���`�<��J�J�P� $π=�� +π4�� =π+�� Lπ"�� ^π�� gπ�� yπ�� ��L�ν(JJ���ڢ ���d���=dM��JJ���8���8�eM�M�x��8���8�xeM�M�L��M�L����з��x�L��� $πS�x��40���(��
 �π: $π5 +π0���(��
 gπ! ^π Lπ���(�0 yπ =π ��`ڽ��(�� ����8��9��
��8��9� 
��0х�0х��: ���`��P`��(8��(��P`�(8��(��P`��(8��(��P`���P`��(i�(��P`�(i�(��P`��(i�(��P`�  	�������s�.�s���ds�2�\�2�2�$�  	�������t�G�t���A ��dt�:�*�6��*� #�m���������� ?Ѐ GЀ �Ѐ �Ѐ ��`�Fi��Gi�( ��`� � ���
��  Ѐ����`� � &�` ?Т � ����� �Fi��Gi�( �΀���ڀ(� � ����� �Fi��Gi�( �΀����`�� &�`�� &�`�	� &�`�
� &�` ?Т � ���� � �Fi��Gi�( �΀����`ڢ �ə�6���7���� �ǩ��� Y��� 4�������3��� �Ѐ
 �Ѐ��о�`����ڢ �d�	��w�������������� �`� � � ���t�d���h �ѥ[����]��� �	�$��8�
��0��
 #� 4����%�<���� Y�)������8���0�
�
 #� �Ҁ���� Y� �� �Ҁ��Ќ���� L^�`Zڥw
�������轲����Z�d��:��:�z�� �����������(� 2�z`�x������0���0�8�0�����0�	8��0���8�0�'�I�����	8����	�8������[�� �[`Zژ��d�	� �� �� fĀ* ��d�����7� ހ $� �� �ǩ��d�����z`� �Ω�� �<�P�`�+�Ly� �إw
��zӅ�zӅ�N
���ȱex�� �ə� �ӀX�N )Ԡ ����ȱ�+�D� �d���1��d ��ȱe�xȱe��ȱ��ȱ��ȱ�� �����ÀȀ�`��a�̞!������w� �Ӏ�� �Ӏ�� �Ӏ �`ڢ �d����	��d��������e�������`ڢ �d����	��g��������`ڢ �d����	��h��������`ڢ �d����	�
 ����d��i�������`�w
������z
������N�ȱ�} ��%e�|���{ ���z`�{���*�0�&��0 ���| ��|��� �Ԁd{�	�p��� y�`�|��}���8��9� �2��2���: C�`�,�3�	�, V�X���X�dX� �d������ %�����p� Z� �`�-�3��- o�Y���Y�dY� �d������ %�����p� Z� �`���D
���ȹ�ex���
��}x�xȱ}��� ��x8�0�(���0�� �� �Հߩ��d����`ڢ �d��� �եn��� �������`Z�w
�������ȹ������d������F8�x0�$�I���G8��0���I������n�dnz`���� �L���� �L���� �L���� #�L���� '�L���� 4�L���� >�L���� K�L���� U�L���� b�L���� l�L���� y�L�׽�� � ��L���!� ��L���"� ��L���#� (�L���$� S�L���%� ��L���&� *�L���'� ��L�׽��(� ��L���)� >�L���*� P�L���+� ��L���,� ��L���-� [�L���.� q�L�׽��/� ��L���0� ��L���1� �L���2� 5�L���3� �L�׽��4� ��L���5� ��L���6� ��L���7� �L���9� �ހd�:� �ހ[�;� �ހR�<� �ހI�=� �ހ@�>� �ހ7���d� �ހ+�e� �߀"�f� �߀�g� S���h� ��i� ��`ڢ �d���#� �d�!�x�"���#���$���%�� �������`ތތ`����`�x`�x`�x��8���`�xތތ`�x��8���`�xތތ`�x��i��`�x����`�x��i��`�x����`���< ހ'��)��G݌���������	ތތތ�x`�\I��\`��� ؀�A�G݌� ؀ ؀ #�` ����x���x��)���G݌�� ؀ ؽ�)��F�x�� #؀ �`���
� >؀�� ؀�� K؀�(� l؀ K�`������������d��� �d��8��� ؀ �� ��`���
�ތތ�������)��x`���
�����H���xi���i�ڢ �d���%��d��x����%���������
 �������`�]eFm�mz�])� � U؀�� b؀�� l؀ y�`����v�]eFm�mz�])� ؀a�� ؀X�� ؀O�� #؀F�� '؀=�� 4؀4�� >؀+�� K؀"�� U؀�	� b؀�
� l؀�� y�`���<� �؀ �� ��i$�x`��)��)�� �x�!���"��#��$�% �ש�# �ש�# ��`���� ؀=���� �������G�
��� '؀�� U؀�2� ؀�9� ؀ #�`��)�� K؀ y�`��� ؀)���� ؀ ؀������G���������`��ə�)�x8�F�� ؀*������G������	�����
� � ؀ � �`������\ �����9��G�x8���x�!�'�����
�������xe\�x�L �؀� �ތ���G�:��� ؽ��n�+�����\0�x8���������e�x��x`��������� �� ��`�������� �`����J�� �����������w������������i� �x�!���"�0�#��$��% ��`����!�G�:�G��G�� �ތ� �����x�F��������`���( #؀�<�G݌� ؀ ؀ �`���� #؀=�"��'� �������G�
��� >؀�� l؀�<� #؀�C� ؀ �` >��x�x` [ܽ�)��x�x`�6�2���6�� �xi�!���"��#��$��% �ש�# �ש�# ��`�5�2���5�� �xi�!���"��#��$��% �ש�# �ש�# ��`��)�� ؀ �`�d� �x�!��8��"��#��$��% �׽x�!��i�" ��` ���)� ؀ #ؽx8����"���)�� ؀��	�� #�` P۽���x�x` �۽���x�x` ��x8�� �` O� ��` O� ��` �ڽ��G���8����
�{i��`�u��v��dv��vڢ �d��7�������� �����x���x8��!��xe\�x�3�\I��\����4�%�F�4�� �x:�!��i�"��#��$��% �ץ5�/�
�5�������e�d��e���e^���	�^I��^��`�u�*�v�&�x�_���`�F�a�G�b�f������v���u� `�u���A�x�a�(��x��x���b�n�b�i�ތތ�_�����W���b��b�֩��u�E�x�_�(��x��x���`�-�`�(�ތތ���������`��`��du�e����`���P��4 �� ��x8����xL� ��i��x����x��xޠ�u���n�6�:�d�6�� �x�!��i
�"�*�#��$��% �ש� ��# �ש� ��# �ץ5�/�
�5������e�W��e^������^���^�鞠` O޽x8�����)�� إ5�Y�x�5 |�xi�!��i�"��#��$��% �׽��" |� �ש�# |� �ש�# |� �ש�# |� �ש�# |� ��`�_���_�d_�_i
� `�4�8�<�4�����������i� �x:�!��i�"��#��$��% �׽�����e�e��ec���	�cI��c�콌�G�
�G��G�� � �x:�!���"��#��$��% ��`ڢ �d��� �������`� �� �d����x8��"� �������`ڢ �d������ �������`ڢ �d������ �������`Z�x�����d�ڥw
�������轲������8��9��
�����X��Y�0Ș
�ڥw
����
�����
�ȱ
ex���: ��z`��&�N���[F\�\�\]a]�]�]Q^�^�^�^�^$_�^�^�^�^_�a�c�die�eef�fef�fgug�g9h�h�hQi�i�^�^�i�l�!"["�"�"7#�#�#�#�#S$�$%[%�8�8�8�8�%�)� � � � � � � �  7.�.k/p0�1W2l1l1�2#3w3�3�8�8�8�8�8�8�3o6��������	
	

������?)
E@����ڢ �������8��9��: ��`Z�
����ȹ��� �}�ȱ}� s�����z`�0(��d��0��8��9ڢ�������: ��`������ ���JJ�`H�Z����dd� �i���j�����2��:�������%&��������
���Q����(��i(��i �d���8����d�����9Ѝ��z�h`H�Z����dd� �����2��:�������%&��������
���Q����(��i(��i �d���8����d�����9Ж��z�h`H�Z�������L�����������LA�����2������L����r�����L������LA�����2������L�z�h`H�Zd�@�� � � ��������z�h`�Z�P� �� ���� ��z�`H�  ����h`H�Z
�����轾��� ��$��a��b��c��d��e�8�7�; ��Ȁ�z�h`H�Z�7���=�7�y8�
��U��U��<
���ȱ���8��9�;�a��$��b��%��c��&��d��'�e��(
���ȱex� C���z�h`H�Z)�; ��z�h`H�Z�)�JJJJ�; ��)�; ��z�h`e�]�[�� � �@�`� � �@�`�H




���)�& h` 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P���@p�� 0`��� P����������@@@@@@AAAAABBBBBCCCCCCDDDDDEEEEEFFFFFFGGGGGHHHHHIIIIIIJJJJJKKKKKLLLLLLMMMMMNNNNNOOOOOOPPPPPQQQQQRRRRRRSSSSSTTTTTUUUUUUVVVVVWWWWWXXXXXXYYYYYZZZZZ[[[[[[\\\\\]]]]]^^^^^^____________P���P�����������DLE�EFl�,���WPX4�U���&�+�F((AZ�d7K<�<<�(7_P���   3  3 ��? 0 0 0 ��< 0 0 �� �  �      ��     � �   � W0   ��U�   ����   ����   �W�   �=?0   |�0 ���_ \}]�5  �WW��? w�U�3 \UU? �W� � <�                   �      �?    \�    WU  �W�  �?W�  ��_�  |��� ���� p=��0 \�WUW �[UU_�<|U�^1 ������z�% ? ��W
     �             �     ��    p   \U   ?\�  ��\�  �w�  ��� �w? ��p���pU_U]�poUU}���U��� ���
   릖    ?_)     �      0     �?      0 �   0�   0pU5   �p�?   �s�?  ����?  �w� < ��  ���W�?�UUUuU3��UU�U3������ \U�
   ��?    �              �      �      �      � �   � W0   ��U�   ����   ��� � ��W� \�]�?0 W�]U0 WU�_= �UU� _���  ף�   ?                             ��        �?    �    WU�   �W�?   �W��   ����  �Wu�5 �UuW� 0|��U� ��UU��  ���o�   ����      �                        0   �  �   W 0  W�  |�   pͿ��  p}��U �UU{U� �UU}}�  �W���  p]7��  p}7�3  _���   � �    � \   \p   ��  � ���� ��?���������?��?�� ���� ���� ���� ���� �����Wu�5�Uuw�0|��u���UW�� ���o�  ����     �� ������ � � � � � � � � � �* d�dҜ ����d�`�������� 񥧍 ���  u�殥�ũ� ������ 񥴍 ���  ��滥�Ŷ� ����J�������� 񥋍 ���  �磊������ 񥙍 ���  "�撥�ō� �栥�ś� :����� -� ��`������ȱ���ȱ���ȱ���ȱ���)
�������������)0��ȥ���������Ȅ�d�d���� �L� ��� �
��� �d���Ȅ�d���������ȱ���ȱ���ȱ���ȱ���)
�������������)0��ȱ������Ȅ�d�d���� �� ��� ��)��	����d� ��`������ȱ���ȱ���ȱ���ȱ���)
�������������)0��ȱ������Ȅ�d�d���� к� ��� ��)��@Ы����d� ������ȱ���ȱ���ȱ���ȱ���)
�������������)0��ȥ���������Ȅ�d�d���� е�� ��� �
��� �d���Ȅ�d�����
����������ϱ΅�ȱ΅�`��
����������ϱ΅�ȱ΅�`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ɠ��d���� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������ơ��d���� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ư��d���� z�h`H�Z��)?	@����;��%����������)@��J��������8������)0��Ȅ������Ƽ��d���� z�h`� `� `�˩��� -�`H�Z������̩��˅ҥ�)?
���������d� b�(z�h`dҜ* d�`�ӱԅ�ȱԅ�ȱԅ�ȱԅ�)
����������ĥ�)0��Ȅ�d�dť�� Z�d�`H�Z�����L%���ɥ�;��)��ɤűê��)@��J��Ʌɥ��8��Ȁ��)0��Ȅű�����ť�dť�)����)����
�@��������ɍ( ������* ���¥���� b�z�h`H�Z�  ��  ��d�d������ � :� �� "� -����(z�h`H�Z��� ���� �dѥ�)?�ѐD�� �>��
�����������������d�d�� ������)������ ������� � -�(z�h` �� � �� � �� � �� � �<� � �� � �� � �� � �� � �<� � �� � �� � �� � �� � �<� � �� � �� � �� � �� � �<� �     � �� @ �� @ �� @ �� @ �� � �� � �<� � 
� �
~� 
}� �
|� 
{� �
z� 
y� �
x� 
w� �
v� 
u� �
t� 
s� �
r� 
q�     � ��@ ��@ 
� �
~� 
}� �
|� 
{� �
z� 
y� �
x� 
w� �
v� 
u� �
t� 
s� �
r� 
q� ��@ ��@     � �x�� �<�� �x�� �<��(<��<��(<��(<��<�� �<��<����(�� �<�� ������(�� ������(��     � � � q� � d� � � � qp� � � � q� � d� � � � �p� � �� � _� � �� � �� � �p� � �8� � �8� � �p� �     � 8�� �8�� �8�� �8�� 8�� �8�� �8�� �8�� �8�� ��� ��� �p�� �8��8��(p��     �(�� ��� ���(�� ��� ��� ��� �8�� ��� ���(�� ��� ���(�� ��� ��� ��� �8�� ��� ���     � ��� ��� ��� ��� ��� ��� ��� �� ��� ���  8�� ��� ��� ��� ���  8�� ��� ��� ��� ���  8��     �  8�!�  8�!�  p�!�  8�!�  8�!�  p�!�  8�!�  8�!�  p�!�  8�!�  8�!�  p�!�     � �
�� /d��     � G#�� K#��     � �#�� �#��     � q�� �� ��� ��� T�� �!� ��!� ��!� ��!� K�!� T�!� _�!� d�!�     � ��� ��� ��� ��� d�!� ��!� ��!� ��!� ��!� d�!� q�!� �!� ��!�     � ��! ��! ��! ��! ��! ��!     � w�# w�# w�# w�# w�# w�#     �(�3�F�a������������2�9�@��5A �   �G� �5� �   �5A �5A �5A �   �U� �F� �F� �U� �F� �F� � �   �h� 4�E� 4�V� �   oA �   :A �   �� �X� �   �� �J� 	�J� 	��� �Z� �   �A �HA 	�HA 	��A �UA �   
   i   �( �  �  	
	�
	�


				�				


�

		�
	�				


				


�


	
	
	
			 ���������������  ��  ��
�  ��  ��:���  <�  M�_�n�������|���������� �f���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   E� ���